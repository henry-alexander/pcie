// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZWdf4m9/UA+PizLAc/79TxmaHKuh87Teq+fKUrx66N/01BuZnPbmE3A/Ooa/
dckgRdxLdEqbUCSTWRDRzcezCIA2RIB1kSpFLLtwUolarI54f8Qyqiv2lB2i
9/xZaYXekenpeQnz3s6y3ZHnVRdOZdhPOyOY2T7B0JVs8NNjqbbGX+HO9ClL
EzLI7qvIBSawMS57yomAJSk0yYMSXheM2eiEXgQEvOSVgxXdueX9ANrHgzbU
8K9E0WIXYMXMJRqyYO9RSms6/9W2n2aeFyXyiCEjfNYuuGW4soQKBHoxIw2h
bGiFMUfVLhZ0J35IikfkGTYTd65DaiJ+zqwQR6AiLw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IEowuadQY54KnXBfpfw+GmhoppTN6qWD6x/GivZ4iO8jOcC2nen0sCHEou3s
mQl26WwB2Lzjd1ev9vjNmUnwqoFXVnskh+xtCS6xHagB0Md0PlcpHgG1z3r1
FHmOB0n3lQSYsOhdD0Ub9s39XA/KkP0ZCk3KCVcKLuGyi3Df7CAsb2QBjOs4
ZfKHN7j6qup1gexgMJF7WCTjDGuTJKbwRgFwoyZTJWYib3/qvvwttSHXwh1+
P1LMbAIk+c2RMTpalTCTFwXu1LHiJdPnakX9T1DOBHxbjBK+iy7WIC94Ujjk
nYSZvkRGth7FFQPaOz6J3vk/ir/H8VvCzxVwLX1RyQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nSz5xsNSybZN7WvYWTTOZfZ/x053/+cXEsUQNS8jhjDd7bJfTINlSmrT3Png
LwsdJALRJj8rdk/jpsmGCffO1mQEQKBIiyA8c+PJJnJpHcd7J860XfhtCunQ
A/RbK1tcAIcUl9Je0o4Hj/8MVChz0jaUVDtZV3W8up0UQE0OElHfU86wyP4Q
9U046W20vb6U6HT9kFIT1ruIVy+E9aLTPRHS2+jBRZPD3T9d416OlGR3Mpw/
MdZuNJR2u0Qd8VRe7Jc8tJRG1OFToWzP8j/RsCpLThz/OPZk0svWpdH/j67j
UcovhuE37ehDdhFQulvVLDwpD33qwagmAPdDLGJAlQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bH55Q1y3Yb93/PFLIV+qkId0bLRlQVe4e62LidBmxlYwiIPVr6HSzIZjwZwf
n8tQKpiV0jXV2J0RsPxi2DoRzsRumZdDXQxIBLfO52xRT5TAe07AzveiICue
m74WSDGyDFWnXzjBByUIgBs/Txt3ikwVQvLNDgrMRfIRroYAGc0=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
R4GfXeNXymQiwws7bq9GzCULV6kjnTagrs8Hv75P0yuJ0u6tWYdpuNgULXgl
aCqnyEmaCnBGdsa8ij1tXKmKkf54DwCfsu9CiLbI6EiFHeOJhBf7HAk1HULr
ghzLX+bRZN96W2qsmLPaZI2aKyP820rSioHTpapDPruI9UGKjbnGPSNIngsQ
NZK5v/ulateqnEOfn9VhGuDS5ueIlIMjDuyRRnt/CTGKzt7I/eGUa2Fh2del
wr9FLSgf9wKVeAzCxOWigh41UccCi0NvtGApafBIegBmYv+ddw/cNiizX1yn
Eo7LPMWPtYkz+PQY2+JnCNjLdVqzIynQtSzNhLWWxMeinUSiBDpYJ6IYaFXz
njNzspBlp2Hb1ZFZVqTgaeAGWj8DCCRfOzUJxUZMcrVz0BdHDicnjR9/WBQm
HSsfoWaI09x5AGQP6mj+U4ilYMFVLX+pvh7rGp8wmvv0k0Auo9MGFMoobm/A
Tg6cVKPvF7d0TiRG6QDkftPfqehMUtgt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r7KP18HrHBxnbPDMOlUKosYJpXF8boenGHM/dlrfPzPAtzGoWBqHtiMvTGqq
5WH8BfxdWqX+4DwXpZm4HVhqb/uI3J0K+2kvHc6J2eXJ4y4suZFqz+WFG0o4
wqNxDpdGb6tB+uND5+PkywTtT8/FMMcPsHqVjXXP6DDGyda8Wq0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dr3hoAS8EhrnxEnSCqO2HlzcNdUNNSA9540iukBVmWXzrZgPdDa0wr5Jhjb8
sIzMCOdk1k/WyqP7HtZAo1rxbyIbuAxiqWpiSnneRXcB89CL3j+UMfgGwljr
Ljc0tRSmcOC9st6ik4l3/2YMw/210mzz8sLKrs5Ix1zRGpuU1Yw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11216)
`pragma protect data_block
aZ5V4BzJ4s/woifv9NE1TXFOFUaSQQ/WHHE+OzNAaqNGlL4RSmw9HdTv1YTO
v4/vT2E1+wM2Vm85FWVcJPrm9zefxBANey/ZL5eUxRoWadtnpR4KvJnwHTU7
5F5EBPHEcIni+wkP6/7Ywa4wXJ/ZfM+NCiYoN6wVoq/6pappzUJO0kjvAbuL
hSXBs6BpebsFTIRVvfJugMhaK4NresV8Al2K64I4AJ5AOvTxr7tvu0dVX3np
OxTy5JLN3riVCSSUVMm7oO9vmg39EVo737N9IS2xz50aKTwCyY1W8oMvGqdY
uPcQqsmP31dXsT4+TpsTipDlGnQpdk6fxA7C+6NFCCEmjikiOp2SleuYFODO
a/5qr89FT+Zc5lUCmz+DcbZNaAvvjFbBoi3GCGDypoDg4Q8REq1TS/MCEXge
q/p6TlbqRQIMr/DHBdBPh1sDrnBDxfywOnQsNaQgisDNbr8WMpLzU9zf4sqS
QMdS7WM5ZFpJHuL3v1QmDGdNSMfLzV8RLntV/4+B/y6lepx/33byb87OhpDa
4jLKQ+R5LSiT47qf2ua/kHDm8Bg3JxHQOCIBg0WtTulLWEkm8y/U1wnGVaog
lvDnvL/3mhr98eMkD7WGmMJymgEge0KOoc+xFvtOONVD8bKshfWhfqyvYU/i
ujS8wVeqQ5rFliyt6H4XZAaVV5k9v4ow/E+UcdCap9c4eSqMhr1MJNThy4Bg
HanhEPvKVyBs7CbGL4rznBA/JGArYclj395AcYK+Y6z2b5H5UH3GRZkxwihd
9Y9jVDMZ7visFYwnDHRsV75V/DLjkoChX2Oekj5IVlCrML36F3/eKj7AMlz6
vu4ZZioNZG6m0VnYj4uNGvrrY9Q1DsU3j0Ckbnl7XEijIODumZQh/KfJWL0w
kHxw7g6g6dQDPYJKu0DNXtOgamJZjbveSCvh11tpLfrUxgkQjyZT2bvcumTi
SFtLIjxUdC7xHNXsgLf/6d8zD8TdMEvDXIFs28lDnMgs5dW40r02pzfCRvvt
VVoLaWAU6d/b0aGtsptOSF0fE9pXJUZqF8qgqy7MbcoeCESFPqmweKSFUvGp
luodRdufHm8vEuLcSt6AzbbViLSl0qHc5eLEdPjFzCNiw9g8DaivZD+bdY7b
AXutIPufFGw4LvvB5aSIrZ8Cb19tRZEpiDpG+uBiK/v9COsK//kb09KbknUt
vcva5IVaAtlwKgKOUfHWYhmxTAIxscMr0J0fjsfjDOn1eMtRaAaAeW9WcRGO
4eBdYAWG64dbLRQvgG4GhvDS29jBrZfXUbZiUmqJCdRdU/KwhzOPh1WMEumu
Kzc5zWcTdIZHBJ4Y98apEyIWkW9RFBFrgEVn/AgB0EHBt7oWAFuy1Q4Ulq05
4lXck0h3/rE2G+Kaaxe4iSMmi2mKBhjp8jQ+G6eNncsh9yPs1qWBUmx4a9Qw
h7ofmoyMmIYrjXQdlhj7tJTFOA3qm+mgiGkuIvMLCyJ4gFTamLYfja7VMRSv
3ri77s+1YQzLZkwN4Q5j/MsbCdnE3fwvZPa9O8KdPLpIO02TEoFgG2r9bGTT
1ecAGbZYNmEvhsC1Ng3/XML+1iNXvQ+ZL5KDz/vRqUNRWFx+5qR/w6+4RqW6
NX23c3MyaMiJNOYUG6FTnTBmt99jPkMOLjRWeSbOCr78VyzCLimZ0xZ8++wO
BfUMkbjSU0Wy8Xwz4Cz5+VUg4YishGJLHWjbmPLNUxW/QzTmHnhrajSsrj6W
fBFICjwVcixatO3NAa74KDhaUZx2pZMK5FsPn+usZj0Gl+6W7xGFei4b8E9w
udftZhvcaQgyiDBhEz2TCFCN5+bueE57qsnpIi77fmmYYwp88dS2Fws0h+ru
dmFUlwgs1WJfrV3L7B8J6HImmKNroPDBN3Jd8UwOqHczcfnp+bTdqEtCSKS8
CPbaJ9iYWjLPMeBWtTFFCO8qA0yrWQmUpWt0xXuWCxkzSdXZcdxd2E0W4EuP
xuXM0QadbiJSJRWH0jvPYsyxCA6hZU6Lh81/HhAPxrsdzjibH0vCXEo7rqHk
mCVerJSorA1q1bGo59P7wN+BAPTQrIeSqjpcmhEGxz93JdVWTbDA0ABlNtzg
xe7G4vqYJ/3LFkVC71pWLeROYjgG+A267PMzAhbCa1aYRiAl5oJ9q6HkgXYs
6VeNnECHcCQSkiV58+l0hen+dEiKVJ92AyAgi9oHBm/d53TopTVB/KnmMm5S
+n6ezYizRjfRAIzUTChIIcgXTcxstd3h/FvZD/+3weuqw9sgSqVwIvdtV+e4
R6IH6ga/gpznEUny/kIw49Owbm19Hz3Izj2o18mUg6HftYA9woED06mLltDV
gcKYUDVlKtdqV6BDyJS1bzHpA9sBE4ICvCrYhm2/GB+KLK/Yu69et3CQ3Z63
YKXLXN/p2xcXlc2/PwUIkfVsNSlUrqd407glRl/EYSNoKWlRPZ/g1zn0SpsS
0eVWIp2BbMzHvpZ+9DNi4nXj666W2KmpR2h47uEsLR4dfa1pbNz5hgryo0jU
s9Egdxyb6os4pV6YKNlUTlKmjPsmkxxErFLLia5JbbzMmUcfdEDcrLhu0o0L
/NDda00Gcj9TBA9E+04EKUmMqhvxDsGiwHLeBKkOvdDDmFLqc115o/1IhUYk
cGW6Kv0JtgEhYLLWcXbVE6KWKZ59tBnI0YTeViChswz/qPhOeLhjy/G3hfRU
uPwkJfXMmT8nWV1OH7ZT0FUgFSnpFmffB5Ci4jXvlNVeF58uP/eLV7hX9JdS
mekKTVDjv7FzKZSf04BnaOzTTr6qKgAeNOTpkUC4RXI2txpYXVY+lRiAss60
CJxI9SfNLCSM24axhAu/F+729pNbHJoF1PuJjETaARpaJ8Kk83efHbKZxqGZ
5M9PYAfNlrdlkO+SVs9VI7s4JIxa6sqYGfD5TaHur0Kx45DkLKK3LZgrt6Qz
xFT5lPKHRExA9eaeMU9s87VLZ1Hls+7CJsH3e4/9OkudEv3tQZW4GQwM/zUg
jqTmn8NLbHkvkH81O+B5ujPfHJeTeNZwV58Tm5CGBhdgXRMpFy0lvkcH4FiC
2fA5K4QhCZhXVHJdO1Im7wddJ6w614olsDDAfY22tqjNOl9z8gjYB8QlOEwV
P9485E9YcEqkBMKLKwxDw98KZXfuW0TpW7iXolVWm7enNQdwKwekBYO9b6YA
yewJnoNmK7JNknXGcFXZkpROvfyBoMk2cPfYyoQT3gWrCFtMsWAyujv6XVSb
L7Uqtq+LnE8rYJ3Y0AdYIF/F1Oo0CyGjxO7I7m7i54XndjoepbfATQnT+pwx
nm7uzgm4THrDWnQrt0WvhhTTZP/h61kxs0kB1H914mtak1Ouu5xgB0+NdiNh
hU1py9ZDSayazKz2GOWnQ/XfBW8xhR2eYjygZeBcgd0BnJfs4dsadCPsRsl2
JwftB3MepxE7Xc9UGbPDaD22hPMEoLco316fDHw5Y/RbLvU38A4hqYCTZyZH
9CuAws6hUsATNzEPTO6fw7gKpyaI7pDomYw9UMwR+uHJQB6uRNeDsydQaGi1
qyVQWLjeYq6OUCUhCtiKFjiO7QhFe8g3BVCqpRRNLMNItqO/LLwHbf8YX7/o
Wp1tnl4ta/XiPf0m1t3X4NZCHfsodSvmuk955fa8st7T/nCZhlUEqqwnvvAs
SndaToydjitZtTx3/Om8ZM62stctUOPgKVjxnArs/w5nYlJCPPX8sFLA/Tmf
6HirABBJsDiHO2NYoxQPuEp1APmaYqvtlRnOBIhYIlHVg/LPM1hau4c8/yAt
sg5g2LwHDTYVKEhfelSteUs5Wa7KWC/nvxUyUHQAj/oBetsY6CW7uM9vcS4A
CEGGSV94YkOOpB4CFm+2a13EWWlJaBcvYOOdETQBpPGleYdWwL/WgrMhFuhq
i6ca2VAADhGpCbdngru+sLqGg7bJ/DQ5ziANJPwb+PK7dn37cbUvoWLYNJoR
8wHeBqq5TPueqY/CL1la84BFr7AoLum5RJ7Al+BHeMAiAbH1SPL6eAsav7IH
YdNs9b9ktow2giCLMQwDjwyt/Af+Kjz6TpQRUKy+M/3bcygZ8XTrCL2GW717
wJRV2RWaRJtULz1w4BgTrbY92UewBTvslgczs6UdozdqFdjl6EPyKohAtuE4
rhM6HgjPfHpNcmWOvam0a+eZvLnRYvgaZtJNAs36HTZbL7kl/sLbI13gsv7P
voD+oyNxpJncO0boNfY6QlFM44QTSldrCuPaRbXcmwWYdK+NBnwOK4lYFNRL
HoFRNLKqRurkdP6UpL4pYqrKVIQwk01TyLMvUrZTRc4AY4gqhqliCZvPw+9Z
MaNouSzsIORzPSsVO5LythSlDGCtSKVCtgpsrg31WUFOGgcQfiUYpVLrSxG2
HXUhu3iNPCLLUjp/LzjkZ7HacdMm2KSRXavUAMolUh78OjLbyQO4h/sEWFjK
pHFxrPjUHmylEdtt+Wag8lBFR1G8mvxFLri6gxH5/JEyZPj1kGIk4GTt+TqH
yoJVSSoUz5g5V+mxWLcwGXxiFMH50U4yNt72koovPnuutL+kAibhUaDbyE9E
kr4yL4PW+3lpKTBmMs+ArSu5RWiY9Y22WlS2diSEKaUwE5KY2YwRDP96dXki
glySXJ0bpfFLEhXyyXVbNG9TqALv1UECA5rWsraKUNrjZdnSZnBwP0XGRF4G
yg4d9sJ+hzbjHK7bvNkCJt1sglJSBeONS8vwryZpDRvxvQQcj8FGNhS2tdkG
+hd2VY44etZtCrTQOEyhJykLixABAu61E3Cv4yJn4CpSzh8o9tX5vEPYfpzg
k2zMAoPFrSm6smrWvux3L7qUQiORayfloIacOTcaDugA4UX3JWSwd05uCdLC
DmG4GyNP3LecdzWIxx2Zpg29IjrKy3WQ1s1xsRMf0p3/6/2C7MGzlql8X9xu
H1Ct8MQBKFazJtYy6rTtl+lzlWKlGC05hW9lhZn4NQ+o5cWBipIPkvRExqP/
KVE6bh67nUW71CMZClYwpAFOshInNu6MYElziEYlrIdTn1vGGAnmeiQiJ2Ba
ktIG1MQQp8YDqoiuRMZbmfekYJyc4rMtWF1ejZ4sQfd/PULXB+RRiA0MTEuZ
RP+jL4gq6eWVG1fj+RvRl+c+zQ2yAdE0LPu9WBAXVRZeNcCiTH+ivy6Y9m06
3AQ1i2Aq4iMiPR6KMhIEgW/rtSSCz9xEEPins1zjVImBufX8CcZhnS6ROhGN
6dZmii2PecZd732FeadtGtPG6Tt+p1iY1mvu8dFn85MHwyIg6NQKGNIkB9pi
BtIGE2wNGE/bBS1icGP27LIBAiZCunai9kFPuuwHfwFbPqjbYLH3phdsSNe6
syhhXVAhaFgiWQSw4Geau0T+MVLbCPMlYr9jUXIOhnORnTRZR/YJRvjzPyOT
0Gyn9wF3/4/+So73QW2ltmUxqlrJJNnpqZvEumHzqg7zx58eL00GwiAEHQ4n
3yehKvfnEhTuVja+hPLwR52g40+HZwcVlf7hiQv+y9dTWUXOo4vTZ+RSNM0e
UcNdpQ896UUcv1BUk/6FFMG/I37SYGMLcA3cWY50V30QFOA0xZbpNIA+ODTk
X5aLGqU6xPebbej856vMK2Ax06SRyNimmRBSfK+5agSvIb3TmmcOEA14b9qk
aE1fdsXQS3mO/UaRVeKK/FPmxHC7ujXAoiIgjRUBDucRS85DIMeOGTi1qLID
dpVpna9goIswGWMaVBpHCyza0QawXuq4h4f1FHFXyCo0IIi4Ix2gVSkfHzkG
rQS96UJ29pnn6aQ5NoeW4eEvsZXnz8wJ8lWCqp9eyP/yzpazW/sOR0/zEAIA
9JbLCRqacDqP5NlZ85XYjMQwthUKJ80PvR6txIgBn4RoApvTamHs1+egRalq
JuuIMIBPjExCALnS3IrqTfQzylk44a5vwHYxXtd0wKXR9ojCKiwDKFPViA9P
UDS6n1vjuu1Se8QDAsD3TO8Wj45L6nr/4UlDVm83glaix2ZnuSz1wrc6/hbd
u7EqZTlNY4/5o2BbI1Hv0VS0Koi/cTrn5xFQY9Gxxe5q7B8m0x/hyLW/NLTp
nkzR+T6vQPsMKFNwyNFDHBzZjjsRBnaBkclGlw/19NFgNpMliZkxtULhWGQS
B3tkcDSBwNAVSs++Yv1msrJTNOTUiH0NQQ/vIrQ1tr1mve/n8YmC7n9d6DyO
qsA9ynn/HrufuA7pdOeXwuhDmUbEg+ir02bNywaZDDz0gDWRqt2BP5RdJUoe
7cAXJBHoU/+FHtOrbngZLkSf/fdGMXpKIg1DMVzaGqIKZHHhyPqbgUnnByIr
myudUuuPFHTufdIxO2OhnDzQCTMESS219qDvF2naNWxAovjwyrO7tXTY+rZV
79f6t2CETYOYb/CfJxLUwOD6ZI8evQ/WZ005vMc5rwMIZUvxqnVCIa8r3TqG
rAg9e+sko7tVNgplZ2Z9zaUp7hn+rxFnDAjlo3NG9Er+1jJ09AllNxegi6jc
hMu99Z01kYmZJAGvRIuHB9iEXkngxCIeS8nXdlDMtYrdrg3HHTw7tzndRbU8
YpnNPE4WOaxiW474BKHzU5a4Q16+3M6FKnwCLf40689cANhyelpB5cuWc9Gs
npd6n18jOMjn/laLorPRDMTTUgiLNfmTj/e6oLe5fK23zp/FTEEEa3X6QkUm
Fsqv9Kisa3sMQUOEyK7ad6XCN+nMwiiFiMCME1Ukpseyp8u4GpRUSOZiqolr
10x7cwlJJUif3+A39LsClmuenCO3m6x9HAKdk8CRbTdw0EZ4QcjT/81p6B76
H30H7SOJc8Him4VIfEUZ3RvpZhJ0VyQSgC9zAadYKYe7VpJxQVpLJ4pDwLW0
vMyiBbLHMaBw27UW2E0N8zkkEZptlXCp6ip+3TLoAY0XaUIDkPno9khM82Ir
ZO1t7fWnL+2+tErXLvlSg3UVaqo5xbPKL3sudN8COlFN13iSHy2ttfvINvNt
j48ImTP22SoCgdWLRnDT46IN5LV1BGiY/NqejiKImZ4fsDrCbRqaJyc1qTnp
kFafgVEzJThEIrt7i5SGNLWrHlDjRGaIv6CxpNwqcGBf5mtemxdUD+hqkzee
iLRRe4OIO/ZFALIU4KVlZhIwFULxyIWYmkyMMyzd8t40Ovtxy/mQKieiW0rU
4utwlEfV6kx4frUNc8aQ/xLqqZTRsg0C07E0wxfsG+igpld/LDRjvZT0JhLz
NJQv1BtqUW/EUyRICNZH2Izw6zrXJLNGk2Qv6B/PUaCtJk6Ij/e+NbCUBa4w
doWjm7RUN70oUwFFObXw21fdIMAhXDVnwcBEnffj0B9jtQvGphx6Tbcbuoi8
C5HVPEB3k41wCbhoF/pCV18VLdqMR9to/6BFtD6bZgTiup2OmZMvtOMrkKVU
X8C8UxbPj+5oWpeoaxKSyJnmyWRZEpIqqvIrqRWXHgl1YCDadAjod6QkrMfR
9GltSjHnCTKju/vPEQ3yvWvCCJ1JFL9jze1ExNHRuZjayfrBG9a5Exv8RgDc
jYFLGO36z1m3O7TEHyCeBUurLEYZ9d/1cRoAtlGn1ZFaxhARV5gvorClAqAp
kdn8bv/ClSctQw9v7hz9CVswBVDxPjeB0bwNGVKJYSg+rHjicnQnJ4HumJSi
RS6tw4wFQx6YrbBdIzNuiwW98SPMXftcxFANCYDrD0S1Ld8q4t6xJ0Y2fjqd
1WKq/yQebO927o/hAVQ9lINTTgdb3BQRATs35Vhc1ZRVxznJRE2kog2hm94G
lNDQZqYRiujRA1+SUnBKlCP9mHXgmPYpIW1Uh4oe7XJQFb+iyjGo1jn/UXAU
diY4LFadoUApzK88TtMK2yXt+DdKadPR/nN8TD4rA//JPhjXx6qfC9dMf041
4EjOr0sUAwmgUOKy8RbUpm6pKnj8m1tG77W37+3MpJaxLPybtEgE6sgBjbhC
lQV8RkEAvtaSWH5msWc8eKgrc2RPQ8XwbDJ6I1q7OND9b9bkajX3vs82R18n
FQdL4lfukKQXjP7d+Cn/XOdjsUzzKh/nUeRNaSV9q88pCJlKCJtqnt08Wdo3
hKcZQtKSp8er2Eoe/91UdqkmtqZlIt+1ocec0tYgbrt9h1VxijX6/AmkeiCO
oZ7se0PxGSiHLyWtmfY9KMtvvlchSW3GPfyj/02/ZLHPuNKQRM8deXa+/1Bg
+lQYfPwgYGNR9UkraGcNVst5t8JmUIAexK6+DhfPxu4zFjt0YvnMqJcTwjbb
paw6uAS8Ys5Jw6cnLWpDRUfSGXVYcjFE3m85iiaZuqXlD2Ui0ilsXgTslNmg
/bVpmsY5B1FPB5vCIwL9tNNtNH9cGyp58N3K/Ab96IDkd9TKL86COiFhn+Uf
X4Ez/TGBo9Jamt8L8D+OGW9wRytsOo1uo6CvLevzSQ/XYTFwhRT8B/jwgHBe
Vjz7Zm8tutTwB2Po0uMvemNCYXRPjc78CTMNlmi3YWoHNHMDY4QDnmKBFTyF
kp0EqxHOyMBGKVp2zZWxQwAp7ngarFHverk+L/3FIiXNvvLNFPK6WwITavXR
PMyYrEd2Q5pXldUZzpKLGzWeQKt//DIAgu4NXlR0/28h/ctekFQ2Nz0AydJb
sF+DM0a5AR0VBOYg7m2kHWIqTjlDtOR0eDhg9udDbrBfhIj0XdcNqQ/wGBr5
FSsxb6O7KxfNNWMo6A3ZwkeoatXtNe6SSVYg5Q6odc23b0rcmivHz3WUPFKT
JTEOYfNZIjvphx1f1oyXNr7/VDbyRvo6oL+cD7SD+lqbjLhGSnNTmNQ3GoYK
wQo0h/PhrGsULIOWn5Pn9vWiU3Aa8GXOWJmle2tffc/FHiooTn3yxqGM4j2j
F7O6Pm+imiJiP+t+QpvbLdUCf8FX2iIrfMa2+PSYPVO0Vvdpfu+WRk2/7Zc+
kHhbItkVMEhb1doq50jL2a72PTmn5K5VG3LjjkRkok8p9S2/stOhNsqqXtVp
MrAz+1H2DdKXE67zzcE+oaWNEFfUWfi80hZPyq6ltwiABhbcmD5eNZe6nbDi
j9Tfe/YPcjjBHw/yTA3wWOn77+i3YjdL1Ys2jajFnhFvtzATBX5KTnsqOZId
Dmr1Z61+BzONzt5ucops3KuqXWKaaINuUUL0qOS8anEEET+hm3/QnI/TmbQg
cBN3hWarc7hhXBzDv2H/Ehay3unclDicK1zPot2yD2F3Roc2P2ybcDO4UtZQ
2o+BArNdOPrI7wxhWf9Xv/3bdeTJkI8f5ZUmkem9qQ5Whpw2VAuCFicpIi5s
78JiVc97WLg8wFPHvpBlpYixvvyHZ8h0ZbnqOFyFWQA5lgkwrIygSpMdogz9
0LOWY02innUlEpeV37N+kH6fKxdZK5dID4aWfH3+F98WpyEJSc4pu0cREK1t
WW+u9wg7GcJbHwMDaDMJiD++Eru0JisSL/iQLRW/RqHTnHYgxSO3atKVlNXv
IwssbVU4io4+AL3jLfzNqn93hattYhFOvYQ1PAgPN9q0iWBDpD6IEhchkqzQ
rUuo3eYZ6RDA6lo4lDXOqP/9ykRC9O3HDv0RoVDdeKdz/4nnaxE2MmE72grx
cdC294I/HzNrvmA7qN875K9LPSQRjmHHcT5tppDt0ud+1M5iqnu5eMyexDy1
eIfR+ZqTALlzIMUCv1NjCRHkF+BKfNop4SJBl36DS+0rUXar5QCFu+bM4Hu2
t8MiUiffQVPKdHD3S66Tm3bg1SGJNJRhSi74ZW8J1ozKgyakMWU4P2IbyWsy
t+De145jABxpXYUi4dJ+Cr0vp9EmVBru1uFh8yFLapCnv+LAJKGY3DgVUGMU
j38papoGPip8wPNRZS+w+PHm9SSG1UXZbCDj2yKIdcp6Z3YI3JCUDjgr6+q3
EuXNnEQPZ2lc3lwOK9fxUhlxN+t2W03hEp9EabWhiVaS+7onSwoLCSxqXcBq
WMbuaxDeGO2uJFe32/h652hzDhwLM1GomCH+S49zBiwxsOyYrKKrYWSz6G8n
MThjQEV4Jc7POdjZYF0MxWhDnQCK4NaAzhfz+MQiaTpo4gavCFt0mOghO0/n
cTKBWzpHAAfvTNSjbFWCunlJ7Y4pblFNCqkuU8Y499jP3zqzyo8gxZEzhzve
/FehFO08b5huacvkN0yg+pojSniIxH0XNc13LP3v+uTau46GrqAyUqPRfGsZ
u4vJnFRW1hwpOts3ExdI8KqB2WhDXoX2Au/kIWLgDu/3Gn8TEtGYmQr/b4iK
/8SBLyZq2Huv/kvif68PR88FoyKEqDWBfboEn/B19q7oUyq2gwY+jXzP6eHd
DW1MnQIRVXox+ygARS+pE7sMweahpVvJlmODDI4g+FDUmbnXgo8ksf5QEdYE
8+Vm+Vh+v5yzKqca6ln9DiFjF0pi2+Y1zelfpAukD22wAIjIXoSvxyUAmalr
zQMg/57+C/7NRzWG1Z/xIXZpxW8pzwKFUu3y1jD8HiJgfAU/i9AxhmCPz8Tv
oHrBMqEoLYctagx2Dxh/SaTrHoIDQhLvp+dv4qK1fvaf1pHt9jX273uIFx3P
b+UsgpJ6HcoI8b+uSpg8piNAVXuh1mf3ZE3unoEpX+JdjhpLve5T/SFNRsUt
4TNi5vnq0WAZCd56J5EaKVfFYoA+lV6ilrA7tKq67Se3WDAtrz2k029Zuxyt
P34F5F4YVaZW/rcnPH5sogWEdC6lRBHqH3cd7WdXGYOOtIJ+KhdCodf3fsWB
cbVABoux4sPYidyxQGxsHFIz3dqO38B2pSilwBb4foG6cn0HY3AEDDecp9FF
193d08s3oRzHQXFQK1VlmIadNiV0aT2W1LrGe5v6VQk9Z1Tj8wfdmjAeg/P5
iOTuJJ+XI48sFLeZ650jzhAXCcXLdNbc34qJQ1Bxasp86Y3qT3xZnZu/ajWs
4SbXJwqa/JtDXOS+pYQySbuzWh1RktA69UUWCobS8T7syK4e0areKshgYJ57
pEiUCmwPLyG7vbbywresRBXOVO6DlyNHiCvjpM9LO58pLt2gxl9HqA12pY/4
Q0h6/pj53yvVp3JmbI07zWGuhxdLKVdWbyVHZjxCoA2I0WY92xwz1a5nAGYD
j2DOPDO0ovGdVfIJ2r9O5e6GECDavF6iYOLS98xXIX2DSU2a2tP1/oGO18E4
jmfhh5wQGe9ieEaTWMFmO1rs4pmm0TQuHuSPXoYxX44Uk9U7Ut17NqUwkL1k
qUGfMc4KxE0AVpjEUYVl4j407uDas2tAdBqe32Dt1mZQsoHwLAbVla8pK0LY
+rqXPiT1hL4gjE8aLKRZuzCuCu7HfZqfZSBIK/ro+qEWd1BakhANu9srLcSC
v7+Hucvy+cXQmeBT+DGEkbruizBN3wsPD45OlFUYoz8bLF2RxCPr6iEHoV8z
qHXwCWgPoC10wq+8p3P04zXvooRj2U8dHCABG2yBhXagF/PAt6qIxkaK4bSV
y/hMyLDbhc5v70v6uMlJA+cU5wujKa9xszbKNq4dUmkim1puko0OILlA7wb0
4YNrAn0wxgfvjW1Q2Y2hvGB/FhWSsLGaf2xJhZO9SJKUO8XIoc0sew7cKmPr
l2bjrVFY8n7yFqQTDwFa5kpBy893ELzVNfFy6seHxyV/0sDcoVawrHo6uTbD
e0NPTkVsDM3++lLVrdJBzopPYGFTCJsE0WRGFgMwNSogLkfcb3jhNyEuiDef
aIXNMdalyFUA1xj2kbYHxOc78BTeP0/KeaFHU+Hx5bvoQlHXqN/S0tWvC6Mj
YiAssGgbH3UlF24YC7G+ccWU7LdHMGDXGrQF/j86M3eGK6BJx4AMObBMiaiE
a9GEJhDUk7njUbh9zmoXkKxq2i+vDiKpSQejb5yT3EcM9GF5PiexfF/IvPt6
fP7bDl4hKoZuc8oc2KV9xuyxZOq1NYWW0menmTEew6fRDLtuGFaWA4mBB+LL
mUUWTlcKoAWXmILGpAn2DeIGlO1wdkCcK/If2je0cIxvN2xabTMsFr710HWp
ZkEqXUuutYtNDQxiq0dBg/jZh/G+c2s0yIrhKlf9PlrHilfPFTihyvdi1bQq
NM5RwZ9o7CuACPF0wX1HYyYMgyRR26wAy0FJoMYKUmpqWf8izFYBcIakkSIB
KiEaAe/wvFN3k3A/HSs+cygChwzMH4P5IHHQZ0Kh2O8D46Y+C3XfMSNvgiRX
9+tgLz4xn4jviiOMSPhz/Vc3FUmlWFvR0y7lkONIi+Vt8jvszOkHpqxHQDCw
G+vGN9NGbM7ZYZLonA55q01p59V3ljTcVwk7vWol1zWqB0CFS7269DHLP3fT
496qqlbkAjLrbtahTX15Hz4mKwupWtDL8Ag8icZJSAiyfpSIU0tKH6WKjMdk
7Ja5I26fDtASln3++jOp+nX/ckzlD9JCCjNrgNqX+qnS8eOEiJ5xvy3gYQkh
Sve5c3n/tBz8w2UfPuF50/yssqq9J1Nrwr1nvjQChKowDzQbUVV6gssPBi4Z
8lp9axWr924FOHYIY3Vfu5GGZnpi9V23R5uaR5UBYrkhj8Rl4MYe4/LU1f22
eA4PfCdVniBpo/kRv8BP4LKXVB5kbTbV47W+VdIVtjBrHW624T/DBHT5M++8
AKNJE5SyH4UhfKeVrt/CFqStevettawXndDNwrjXJDkwD4D51z2LiQsgQfQJ
hTmCUf1G2eY21yOnvtBaNv9vCMnqY2u6UFgw+YJFFQW2zN85I61Ursd6gqUl
z7CKcqmIwjAjs6kkNQZbujtca13AdcSZzBx2EuggZFkfBVGrFOlLOXR4ErjN
TiO3vP0KaWr6emxLfn2NKh/BVAqups7VGto519uRAAbntyUQSoVCVN9e+Wlf
PM0x4rw3+BVLmp0ENiular5XzKeFVmwAPwqtysn0iGvGxFzgpYr0aT6bQsyx
0EZ1Iik6R1/PZ81tbajGH+IXSMxPxAQ5wbiyLYtjzDYnEVq/eQ4jHpUTubm9
YMmj4oEYUFqyfPa1sxWZsVTW1xl9jgqfZR8YekNOvkpIWw8mFodqWpyTAb1V
YndU7aBSjZVwsJtmzOQhH8GuyNkqKT3hrkaAZbGFRfq91f2QHXyw3ADVXBXJ
rrmw+04P2wR3paNsSjOjhulXsxh9D6vsMxP9kn2ftbmECZurn8rEkbnycMPQ
BWshq6p01UJW3jM6NXgzDefovAz9bmOnl4XcCI7tHW3AFIVk6lNlQyi5v/IT
/m8CD24tYY673AY9qre1qhAstKOvVvzFslFN8DuNZZGY52PidRQmH+1zeKhc
vo3Vn1E6DzJ8f9/EuZFCTaLjSN13jFY66pqsT2KfLZrZD/LazuOuBAXRERz8
rHBGw44cW6+hyF93hBOCNpiypwbQvcm/SQpBk5/IlE+BSV+FmBxjFti2kcVG
ZhqbmhKZYgBIDodGeBAdrx1ReBq0cWDIAHcg/fuMNyZfFCKIWLjvr7tCJa1K
9OjyNTscThjoFcnsdhQ6bGUrumONNbnGanX6dQH+5V/txOptxuXINwnLhdrs
XVrL6lqn5GGBgsN9D8t4g3vAnJZ66mecNKYSTtVwRzL7YKnGMZdm1f1ThcfS
eQjCBCupwPco9ELRcvpf93VHPkJ/NU1mJP5sZe2nyP7i+uA+bVBMyBH3hw7q
f3bRVSlMQCQaK0QkbEkAPYKAkAjdX9dangvRzbwy5fqY1NoxFWgEznli4pYC
FLwP4HBxWXGUKqBdhDA7mtnkmplaNJukDfTnG5tOU+yxnAJrCwtXVXBC0hBw
VRl8lhvl7cFsJYT59JVWT4mz1tV3WHInz/uajG96XQB8RNlG3HIksd5bjT6M
GAVMkyDLGko7KCo/QeVjZEo0in4BzSfbPEJd3+d7agRxsd+SgG/mIRNIdep8
aMf6zZIW7Q6Set/PaS53jZzc2aGxH2hdL0cjGOCsuLPXXd7Dn581uYNkeNOu
+wuM2YHn+FUeFsBt2dVkGk+ycHjmxFcgmVWal9nis+EwyEhsj/iQ4j3B9HKG
LuyCYsrSzPYFVLjkscfNqbYWFr0ydNxr3B5GbvMRWPddy2EuHBqxwlAP7uTj
0CyheWa0K0Wgtpz6d/83OSJmJZMhG6NcQrpE0yjT1yWZliIG29JMZ1C9wTMV
qP9wI9PjwhryQNmBHADodTraB6agi4cLTP5T3y6rPWJhEsHH3Bl63xZdRQi6
chlbckCjHXvcenagz4oNeOey7FKa8VSL5iResVarpVYIkp+Jy9KrBTmrsvFn
ekKWVSHSVRKkrz+iVNW669E2g6DcyOVhCs6BwHB49vxl/8ahKhXIAtv32xHs
EnKRIYDpDM2xLXscdcjVzZSqtAupKTfXU5b3qtEJzgNIlIh6j3nnWiPJh3Iq
/k5usZJNJowkPYTP5OA0VGmCgPelCuPEATjVoLbtcuxqlzVP+JAdw5hg8gXX
JMIS05HTFPvjAceZ8/KJvKG5eyT2CBe4NYkuf/Q7/3QATq9v7uEjtAnMfk6g
VFqS66uWvxjDnhNry7OqRYRg7L3Pb7gFnnVWIgPJgybx2qaj7MGbJJ2uagol
jHAyUsF84xz68WddblbOZp8xNWwcm5rUvmUa9gV8nqiyPVk5evfVfBhhGOjn
lBWFxojIV1yipz7xyTKv4A9ct3iGMgCY15kCM3l9klZIGuCb6qUK0xJlXFh/
QQzzY+MHjA127qGZ8ixp+Cl23v+DYGETEuRYEqINI1MLJtHV/SOF6x/gndMG
MM34nfiSC8n1M6triZtxtH/AO1NJmPKdxkYeT+chGpEjYAWy53yXPMj6Nklt
C4hP70kyg5tQYRtsOQJ0TmGM+IgsSa41LrY1zv61uSnSSDdziQLSGk2PxxpZ
J+TmXfQ8UgKC8XevWT1uHMBEF6hKjvnj6P0mTthBe/mlrao86051nvVAH3es
7jeVaM6UM1LMunlf2Amv4EHXVPg/viQ4zGpgbJ6aJ5EwIPu4J1c/lx2Q8pgc
04zzlWQZzHbJkD5JXXiyi0DzaARPZq8kAihBOwmaCHSZcPe83dfrC2Rx/bi1
rRW9tHIPxksXWk4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q4xnQdmvp8nY9r/47ZmGsjcTyJLtfpvUiCyzan2WHaFfAUUIAhlcmqixrVjltwh2yPyO0c+1ozt3l1MlXQvGI4nEAA+yF9pAqBOW9noSQMP6bsQYR0cfrNTLLO1Bt4bWfXMllL2Ed4mKzYJV6zIIKC63yH4tUNx3+FMqCSNT9ZRC6+PIX4PyjN0yT6LemuQ4HFPrSBYYa6meWrxHk/lbSe7KWX7S3AwX+RXunf+yyLgIfTRW5SRJg/kfVIyaDyyW2XYwk+DbWDaa6kf5dmDfVIzn2fT68jJcYiYPgQ6hUQZ/c/keZz052tyzo9LCHikTVtEur30JjAAc9+jaEo1q56IG9EyBYpboW0akMXjozGNvx5PN0nOQuyVaJegO0SKRyByFWkc8KL+zZcqnZT2N0M3QIl5x+0eORa09ibI50oVbUj0+MeD5vqX/98oqYvrCDBSPr4xfl/X47AZ6eR/tV93Z7tepjqHcN0B1YI5O/siAhVImbNZlIYxa76eKSp8ADoREV//ZhsO5RsxjuLzmHXtJmJoe7rwzH2uOKtJU7Maipsrjalab9iKT3LJXZ7sCtU0LLQcRkKzHh+uqHERC55LgDrPVwzPzfTtMW0FqzAU3c7PK00X8CJJ7hG0AdLq+WeKKQMgdSSRe6nmg5br5SzLBubiVbzPSkFXCVyGreDcN74reiR1KhSAAb9N5bz5Ah2QK4d15Y2BRYYsHAPp3iMUwdnjpMIxffNCy5NjAkC2q3zwn5WVaspLUECczkBzciH7BlhG2w753ATHdedWtbPd"
`endif