// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AE4jvtBshDF4sLTc3YMEmP0tO/3Auhtzzrg0oHB+mnkUrlXQMaBppJChLyaK
BDAEINGqsvhuVZ111Mkxwp9Bo3orJMXXVHXwjFfQGPBeDHopllair8PPGF2v
mk7F0ug+0njSAmyKHa866umvV47t2Auym5SHlP/6jq2JtiU+E6AJBDfO68E1
PdiGeeaS8m3CaJW2rofIazF53SLcOHFcij4wfhf/ymaHq8AqRzLJJp3LN1iS
qjWW1ZVSMHV1DuoUfRRAxAK5Xo35RU5bh2J6GqYc6kxDOzXyLpdC1FD5ABpu
PsPYJ813SJayAmkBbu/6ByJFGuAMJCVhmbsfvhvMiw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bhbrhtFgVQeLMa8lYYY32eWNAYm9qRuKUoQsNLZPvpd9Wf9eCRoBIlMD3EW3
p3nbT1atzKe80+bNBgFxmTa1SG80SOa5y0NozJ6sMtBRc9GblaUMwo1DWr+C
4ntTPQBRVUEhwPY2flnO75uan2Fgb/UgUpKogxvAlOe+3W9asdtDUUItbTJB
hKouqTI81cfQop1NaHKXcs3/z7zxaYe6Pe7sTtDLEEMM/wcs04Z80ik31HwM
t+HXc7EFWavlczb9ErEUc+CyDkAoiXGcJnZXpXcO/lbWyW0vZrdpNT18h04x
trNapQop9yHMSDmiacPDOIFAD40rggHzVpOnCpHAnA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nyHCtzxcLwdPmBwL+Wlez4bybF4Ev1LIelu29DuVJLAxh1bKTikffmowx1br
czSy631Rih7qi4GFzOmq2GYNOWWHdlR+UD4WqXaR9qfg1C0VEQWbe5wBOlK3
r0p5xIBzy2rwAZBJ0NKvwOAj4lyfbWyoWiylWbD4VpX09xuEYqqAVLu7DOfE
FuPPjdLajh0R0BnCbZJJpLflfTebe/Z+f56Twf15rdaRn3TRPkHAaClgYUES
go0HFDbKMy5ZyhGo6cIZLdftUlDsNqgzfaOBNw2YuyRGNYBvnH64txdTXG5U
3ajSgHTwJj7eaHxscKt/iWRlUPOClkATw56nNw9Uzw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iGPy3kjOXjGuFJcW3l1FoUEDC71mBXZmC6PoqXt6Q6VJlLt80ugZO0vELqkD
XwtGdSKoFk86xvItqNUuykAPPSqiIREqzrpwZNw9g2/QuM6I1jz6g9Fk6He9
TeTyZ9+DDLOIGC+IBVXPgxBleZWAb2lgbvdnL8G9B81mjkYmrwY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
PIDpMOLRbPqR2s1/zL0Bi/+Fiyfa0wfg6g6Rq7jBW7cRJtxQpEXFVR3JgzWK
TmBgnhfdvBrXbSsSvyrIQw1wIUDmoEucraSFxYH8pjtYieodM3/KWCnsIYhL
SDbmV0/JiEMCdInKenrAQqsgYUaLIQg71T0xxeKNqzpIZUTBf4slluTEgpFf
7CIMOz4qlBA2HfDP1TvFkwcn2SOqDJxhSbFhsq0CoDocEbDA0DJfqhOUHRzS
deZFc00d+29SRVE9CFFb5YFTjBcfHzIXQTqnmo1HlYl3LOOphnMuUwN1PUbx
094d1sMnSJ71PN3Jj4R5DoHsU+YoIsFwj+vePUDkddh1/4jddEPcYJ9bJhEm
h0qSj/ASH2PabjgozsVln6+HrWiX1DcwVhYg0REG4OptOLcJfrrQP+LuugOn
XejEV10LR8Tf7yh37szbfp5J3+05+qhULGGZBn/KwTgSlx7xu6dJyFYP4Eur
JGh0Y4oH9TvYM8jb/GCVhOZWis7emnjR


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LnE6xlFMLZqhp4bmizphJ08MhZUknj5tfRmQZ0UWZkQ/O+e9dDKtl9uYPa7w
vLgUWyosb+WTV4oVuvgTl4++lH6ICJ7yd8vTlWkmpNnZ7DA3bdf+/dF5oAI3
KU6btOFwp0qH7xNO9BxGnGStCmvNiSSbpPEvXmr9hNoQ2nnGk0U=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jiuF+Q785+xwwjPLmvLrcgBFg69EOhig3SYbGkYNNxrIDJqzBiAMOy1avCxY
YBop1BWKildu2QAlsYzLOWzuiEtxzmggkb0LxUiKzeAIDQiXZi93hbvtZk9C
LjL3aYuFh56FovN3RH/0WbmBNkNcIltGMQYM5mUeN5TndLza3G4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8544)
`pragma protect data_block
PkIP7ssV1wSHeBRkKlDPUaOSrGyiZWO5n6mWnnVK7eq6LDCnedHp/y8GXnBT
Qv3F9U49QqmF4t1BDvwBKwombOtb143h4xI0TPWW+IqthKjiQWDYGUYbyk1M
Td2VGcXjc5XOD1JkaZOLKsQhg1qlL+dhEAQ+XIe7JhGHd+HjFzvyLfnUqdEK
Jboz4fZ6+xA3Vx8ifkSrMOYXqndBjKd74bXxo4bEJXeDafE0GXjhxghE1lyJ
nfgVJf9G1i9N7B6BnJe8QncHWmGUwNuP9cZWw7NRjQDf+X7X5cUaDYNs+R80
pgJIXkTmmGJwUCPrDXsRoddMuelCqI4rfCxdTZc+CB6/SY483UZUa2ip+zAb
PLn7RzROZ1SHhGBYjFFOqNRWRcxrOI0u7CLWGJvUoGKgPeynnqsdCjFfVJpx
Lym8+bK7Y7rz6sG9VsVKgOA5ZZ6+MuDUO78v2SF0y7WADS5mlhaIk9FkD6IJ
ONPuFvEbT9x9FjH1lYirBldDyqYE6I3US+QvQhjFUBgTtc5oYW8F+AiZ7XFS
fpeusb3JiKOijTvSUBoYB+B3nZ99+WtpCwa5UKi4lCkR1M6/Twegba6BSXkj
/a56/TdbCSgI8/o/ee+F/FzDHofwYP2y5ReJeWuYheIlEfI0UsCEQJW0ClF/
as7eEX+cVfGa1GfuA0lczaYEYDM4i7qYmRA8siXrvX/vmndGZOQ+kIQoJF+5
GtzOsoxEataDS1/quLHAtZgVP4zjiyu3fEz8REmT0RasAUbLaATDnOfNSW1b
NWARb6lH4248PKS89xcaIOIlqyCrT0LqYizCFZyx7SE1VC/vlfadyJemGx5/
zopNbNKslRZ+PDeJXCAAanmL642rUOot7L3h0MFHi54cPVCZaWiC6EMCMrrg
kgWQgi4ZsX96MxYfq7rULPs3KlBgPGGjqDEdOqKIe5Elk5ZZ91U3/E7qSQI1
vumlBdjN4rgfdeObACsC65AYM+fM5GVebA4jEaphyNWX9+BpG5Yxy1MdDUnJ
ijr7C5qjEkaJBRVyh5NRDidWV8ofypQpKktQLAfv+iWsFhwsXR7ooKQKkvnr
EFAy9P5DdlTKZMP6etiFU7gLJnDTs7XMMsHYIDXESxaZcUbO/DdDEMPznwn9
PBhIpi/xhP3NjvYPLNZD9Zt9QmjGbz8JDmzg+fq1jidWY8v6HgJmEUCI5mmH
iFCPdg1MZkqQUaFQb86MWlIclTZ7k/wrrto5+QYsyPk0gLse138/pqhzry2Z
Qqe8lFXbHdRPnarvvBQKfT80/rc1lMDlCy/II/Zr8eCKLQfAYhjtPPawFbQ1
KyOfimka2BhQtNJp9RbP59u809ZSVWZTX+io3XTAA5aZLzgDKUmonhbPfJv/
6qnqz4BxJdyUAZ3XsUaVXAvlo6OZCM8wmCJIANL/NHYxafbnBmZ+D1TH2PNu
il3QP7OYtqF72HAAN/ZT5mSc1C234UJfeHB8JYBsiq0w934UDDRjKq2RVaZg
ofVz3Edj6zpm1tbGjO/+FbGOcUhSAlFJu8KkMN2udPiHW8vn++3ocGQ9skfE
pxGy/P8C0SvwthjtDgq/m/IbEipVCaq62trHck9+Po4xdpIA91hCJExOw6pQ
huihmcCBgwxH9N6QiH988mvqtluNWwdhvITJP5/4ZPd8MiVqLXY3wOUHoyez
Kx83EpaxNPe4NO9wyWQmK9//fAg7ewH7/VqbaFLhpdDlWhe/qpw80Cok0GAq
wYG8o+KUw9vvHqaTBxmChczPqi7lpplipx5BiV078pFITDKSd9sjJIdJrPM0
DGdFa1ZnOkCeo44edBKF3IBTQm6Jfolk6sxpJf6LK7LqBUYBrHSopO1vAON6
tzWtTIihjaxgYukHDT5fW7D/e8B4diTfSqpaSGXgGduWqYFCIg6w6xSDYUqC
owtnySqk0//GgpOgRJYiJfQmg8Dhli5FBtOxaZfT+GvF73wmKilrHCKOm3dF
8n731m1MYb+9ZHnoCPb2eIeU09x+o06stL45iU64ohpw7hoh11NrxG33q4Vj
XOXqkRM2KG9sqDF7KtXXJx64K2/tbAPmxt19neIIyYTZXZz4novrwevxk4g4
sd+7K6O40vV7RbrAw6wiWiXLuHSWkn7hAoV0txas5fm0n5CfrYrFNijIuznb
Z18NF13EDrD4fn0z/pTr7fAP9YmJ4cLHmnlYPjYDqFIKWTEhYN5tc6zZLxma
14vGkU5Lg5X2Lq80SeCKnZG06rcmOMc1CYyKg2hwUQHYceq+ES3uIUBX/rW9
anPWsggD65sUId/xejc0XfVNpH+p8uSoXi42tFurydV/v60CdX1etzQVaLIC
9rLecHoHMWxbbfBZATxHtheAQmfxo+NzwAKWqYZUP0eDDIWQ2WTLnrkapedr
RcseKPkP8xOwohozONk4mNSb9Qo/Y/QwP8mFM3amSPr+CQ0BubAhUL9D9pni
zgsM3Mk2S3iAjc4fQATnq1s4skTRjraHn745F7S1uWu0wM/pj2LAiQ2JtZJK
ZKyTe9d3UIW5x35LrwDkOC2chaJBpWT0QIKAr9xQTe9FVzpo33O9aRvVQ55G
2T94ACdJ2vsFy5+LeL53qCtS77F9NYnrorG+ptadxWYrB1pmUM3b7lCgftbl
7gY5wuUuu3KoEQtMHG23SiXgqDnvxI0xk83xaGxOyglIMw3l1Q0/nwjJE5mZ
5i9liRoFOkB2nNzIBJ5s66lwz9A++00sjHDful1fS2g8+2mY+RasCqaVGbPO
pObFPMrCS3nFmrfr0vgBXDzYoMVq32QJhS0ZB2m0HuAvJIaBNAelPf0j0S45
E/jDWcj05TpglsS0pywdgIJnYonFBoQ5b4MLUwS+obIFI9n2GCJ8rSFUZ8eO
kB0Wwe+6zkOOxY841Z3yByy4YYWEX3P1/8JnJRjcQ0LM1tP5nA/TdgIbWUkL
vBpCQDMInxQFpAwcazE7eHj0kp/b/H+ARTvyLNIWO/4YJf8gdi2cW+7N00ZA
Ht7Ro2OSjMLajp0g9nJ0utiR4xEnt1AxLItZBTRKyKzZVhURXFvenKWYtyWW
JFuCAEVS3oKWy7hucS84ps6BuDjeshfsRdzgPueJoGt1iKDY9Wh3JiJgfpzB
22orontWp8Ry2n3D9qoO2X2T6g5PKAG/RKH6tBvokvXbBDCTChTK0Clmrt6X
bKUCG7/UlcJWmbFCmUbaQjcan8VcXxoy1qz3XN9QD6TT0gpLdgOQ2SD0FG2s
7zgLk+yYczj+CglRzP3QYfpG2+kmhPN2XMyLeNceowx7UwT0jsLqvWIJzAcp
Z3tGsiHDk8eRkyMvlInI+C0Hjfvtdl5lY7UUyJ+AjGcY28uQWDF4KIeKcdw4
W3zr05CP5p0Lpx1WPIWhn+invr4dVpoxFYfPDFYjYQfW5GR/eWxf0vmb2XPV
npMva3MsGmfhSiZfneypyur8Eps/0XVNXsE2y6yRNi4OioZN111qX5UaOcnR
FnyCgSRr9Zz+u7rtocb0p9DP7nndde9nKpn6e2cyzrF6sJn5lD38/9DuH6wN
qeFVL1MljWqCHzCT54tJbpGxuU6Hk+81Wmg/qO+dij2pwN7wAbDLfjNWOCCQ
TR5AoBNJFCIRuCA+YsN/l+QJJOUm5+yqbUkN3hRoPvBZCDgyebWLUYw9Rq/n
xFhNTpXHfQZhVQUNE8UOFTa6bbQTi8wnbKAtxe++4EkkXdCfxc28SUho5R2d
HC6aVJav7+I9TBJri7bVtZht1WxeTAndqMvLLwH9oyDw+EZsxecIT97Pussp
dqlWSX/oLAI/IUv1Y4OPLR0hMffCl2f7VRG+mWxMfLC7Axca1X1o4GwER1EW
ic+DDnXyyxJuNrAsYzYRl7R1uJa78fmAJhqiU9a5x1ZuhlzKYFkd3nHhe1tE
NCvFwwS4hhATuA+6A4+JU23e1lXeDycdTg5kh1mFYOXuozQ0ddE+i5M3lqIU
R6hSMXDDKf6QrEHtiY2dGREb9YwcHTkLadywWnhAgueXmJeg5UGQyjO5kyM9
dY1zqlfS9FqRZmE4LLoFgQbEw4urb6N5Du6N8zHiINrkNJz0YV+Od7PJDBfT
5fZsUVTtaK59/0VysoTAFW5M5fKqdHcnS2gE4JjBhNC9dQPqCpo3kPvgwOqj
Qvy5p9s0cfRlTDjOMNLh8aOGWajKITnAs1ejd36GV7LUWTp3aMkPzSUTLd6S
gzotPGtzmIJCOl1R53Rc8XTpcjN5Sc60gbKU2ZH8fCkvQRid0cAyC6knIZIR
sawNXuGUT1r1syXbaZZ5GT6VbAbHSVV/pAL15FhByVGD9oEaWJvHKioJz5Uu
u/geRmpX59mVmjUC+cRYFKR8SEvrwPUavSWNh7mlfrTrxOdnAtiFPGkIlL4G
gd2f9r0rfFMwFbfprrY3HwxUj+ZPeUZWo+X1BQi5Xqx0yI6zn/LuwCoCOzNp
oDNtiwY1JIw5Lm0rIIN1SP+xE4/sR5zl7VX4wubHl41JmQCzuAZb8R5EEx9I
/LJ9P+PEmcEtMqPEZE7EMBuNsApmTAv9UghFl1w79LP3xGUXQLl1vi4wf6AH
4LRYlAAkgABECjhVC8dnv25MY9r54fFMLA88r3OWNx4nk2mt00OhJ+/9VCea
0rK9A/HDlIabhREd4MdMGiRnxdOQ7sxR+atmvmbEbOBY8hT2VByODKy5onHH
XewzCNwHEYL81lelQkhsxHTUY59XES6Xo5fyuxg4b/hwdnGElNiei/OvJFAC
uE4H3aqTz8v8YPRB5LGJ/1SaTNtn5gImCIbNql9xOr3VhOIMXA3uCu+Ock/2
kZpHW7jWuR+eOcZs2QCOmU/wjqWbxBlnR+/PNIqCexAYP3oWUD4wYabNInXA
b6j3KITGdYQX4v6RM/titlsNcP6HxV/1Ot/3eAoduAXpCDMvgKTY2Iw1o4wp
SbhUv1rffzVmZPusYKBHT8TTMljC4LQ1Xh/Al/9w28kmH5IYGU0svx0s1XKt
PvFr/OZmm4Civn2upEZv18jRroav/vLKskkiNjTCJajxnBKS4qa8zA0Lap2E
gToDxIlHspsKmeQw60isCSc4vN+VES/qthWpwC2S2SARfNohhFtW372xd6HV
3a9mjz/lY21CSolpqx5stA93fXVgwWbETVyELicWhpaC7IxzvHBjD1vMkUZu
FAejMbPIYo90bTmhb6sXBsKw6JVNnfvtb2pkXVmMamgPiTjyEGKTO3CT1Sww
aZb1Jj4+Qo8oVA/TCjoD65roXS/UTyK+dqhChHPpZ+kQvdLD/CB/dHkXzpPh
CVltbA9EsGtca99zHJ9W0msiRy89IeeAxNu7hpPxd5yBIY3SX4MrtYlpLhad
k8Uy79fsy9mhFYezjUn7nk1uNFiwxPv19N6NSj8h5kKc1gMEBe08PevtRW0v
9NpieHpRiWxECoGDqtCxrSsRMEsPkUcmFZkSgWVl9Pj6jGAk3k8fqye4aRXs
nMq591qAiTVq48JVHCG0CpEm7SG2sbHJoQWlfAmBMchauI5QyOKs/0ZpNARu
R1NalfWGW7L4QIemPyQdwh4i+4gTyfp4odARrYZEaUay0X1NJ8dZ61QNmPDE
w8YlM8taLeZXr8Lf0DE0UY4QOEQMTP6Ov5BeAr3siHuD5Tg2qYYfw35u9Z9/
kNJv/tk4i6h6lxu9FO38Z2Nnitqq668q21IziMpXX40kD9trx59LmlCPKTFl
C6STzv35+0SSh2NPq/6yU2y3oeinjIAVhjnr8dUZhfBRcx2Syv2sGShKQg1/
z6QIshPmZycSZ4kWPOFRKaRujFduPl5PV3aWaGeR3OF2cn+HLId4V6dpHIQ0
jxDkXge5BVVdhULM0bLtHEdnLWF+UmgNpiUZ6n1WQQI8pGKSBVg92mwDULzI
wisWJjmqJWqQMg0QqG0TV5qHGiW4rHwud78PaJwM5K5BUGbW1PujRmYzb5KW
pIRYGeSaLh+yKBfvHYtxAr3mLB4sqGD5XgNiR3uiGpQtOi0L043vs8Va9RJd
tscC8fnJIYfjjFvO7YFcpTKnmrEUmVWUbFs/zncq8nc286d4jQbfQCOI8wNc
dHtctU5rbMBlGIqLAWA/FXUl4moJPDv7EF7heU0uZduTvDMvx/Yt+klhu/AS
TAAhoaZpBoJ1KO62Cb4Lfo3pW9GIRklWEaIYiKPcZ+KfZtAJCXuJSQZ4YUHC
0hWJczDG2oNY4jz0vSpnwqPQn7vmKA/xU+l0tKR95a/OkAQ/9v6kIkYEWLtK
bNQd5RCI1Ebuq1r08bRdZHuWPemdG7rpTNbmmTYrkWmA1sLpP1NyQyFuqd/K
QN8qgMjhcF86usCFPvsyVszp8qsj1C0LHX7ZayY7K+wz7mOWAQF5WFx+2dkk
XFwLfXdxMX6h3b9qu34ms4/GS50Q1QuTZ4qWl2PXAzYtmsNKFQSMvYRb53mm
ANinQre6CMyORpNSIXTXnrPNa8oPeEUNnOtGeXODpMv5NxTpCtY98MLYubUL
Jvd2HgToMizLO+yYN3rR4Fb8KJ7ax60TaBFWpZJNFK0s7B5rnr4YVuZ4RwGJ
hWukl9ZEDOaXARbtSd969UrvPuyzg0GPoC2MVIp3T3ncyX5yICgrWlD1nlLo
DBpJ2GBwoSZkjIiLGMrIJtw0zLRHvU9AskJfPdFvn3lJgMpdaCABLYoPXwmn
5XtrDLWoCNaMvJq7aFM5nNqrUSNURWQKNymC3xRhYxZkI97BzF1CglStgBka
pbh6k2KQ9NU0qjorCllXtaSPGyfNN8oZay4A1sdqoy6/fs1Ay8WILrAiBJIJ
cHwv1OPaYPV8kxGb5wcYvEFXwyY0asjdP2ETGVqBJnlNw0LLZEl2Pkm9R9+p
lknkVyTzcf1v90DHc/m3ZHpxCz9TidqDBz7RGR6goZ0ByBHkKD5p4+aUD+cC
GxbRcQKDCjVQ8a2CVM2yObESe0xS88kMI4g5sbHT0UgWKxhgrGk1NTfuchPn
J+h5dEYqk48vOPvGk9Zg370hiQE1XBPf/vGcepcAjmJ380g/Jr3p9qae5VG4
tPrZGtYBEYsuY0VW3XchGQzz+qOsHXuL6d6TxU9YE7ZBfwc1O89ntqIsI8DK
ItD1ZmGsj8Rq3mOv4VOOJgoIlladhk/PDON0SlB3ZF3ESy2LrfRjOs4g5V3K
zJZLKg72K54d543aJ4zbeTgxA/DK3mV0fmI9QlYEvkx428usvl6w3hPG3pAK
PCKrQT9G0PHWi1ly3P8sr3JdDHkw+cAqbPUltL9cDRBn+OoiV0J/UadL0S72
BMbhm5YBwUELmAcEtlEZhZpPiuxvL3acOAq6fPdTocBW0dvOa2zi6okIHKeO
HhX8S1e/B/0BoHchXlrr3Kc2ViKlujKw6bColOVYsm5hpSscCeCUQe42lc+T
wLY1qfW05erlGEO/eG13VD7r6dHTcRDjwtEomExcGfAGZ2w5xZ8wXFYh7YXe
ER0K6zNF5Rqc6XmkzVKUu0GoNE+28jNGJwkXH/0DfrLbsOOeQLVOLFw2YKPe
7snvylUAeDpQjvlJGsbtOaMU93St15znIosL1MDB4b54taIxaxFFpcVydmzG
/wHNLB7ujRMjxbR4ZLq4fnVy+LqZqp53FPAuJqqYPnpg8xevMyi14u8n+QBa
Xa/iptPa2eUMui+lC+EfHDfbXaYiEsgIBbTwDABYXLhektBl4SvJS2OaGu6w
BPozjFMJnnApXK/Wg5fBNetJXugHmKgahkVAaeo/vfz2142+aqyoB7osOlvG
/TXHSExztA85IwmCDDYtuM1JK4smBCuK/91GNPhux+mHmZ2BacIgT0YYzFYq
7dyq48bE1rzaKIWVUGkHpwZUCDBUC+ZKDB4vu5lWi9N4Qyx6XaLCgQrJdbay
MlT5vkZCLVST+OCEa4aMbMjwdq1HNF1ljk3Rz5JlFQ601F+Jf+8qGS1Q43Cj
eC3B7wlaKWo7XUH6u5AkzhVZ1rDqAIZ0p6svEly9N9zJKZpzCa7wX1U7KEeZ
xv7m3++nGn2MaI0ylxplAwh+vQAhLqUedPpgH960JkUpto4/Vh61F4JQB9y+
HIeASR5vgl/lMMQSf1JUNte+Q7yFxHyOay1eRv9aM3YTeP2VD3TsV6YM3gnz
Kpb/vjpwDm0bfXlAErrlht50PaA5rB5pNHOFldpkMh1HO59l6RYX8vHMkp6/
yG2l3VoKPcfU17C4xG6cLYf6z75IDbzJsgcWvZ1Icop+b9vc1DNXQlSWd2we
79FZF+B41EHzxSG+qKqsQelG1XTXRabMsstrOJgGLLUMbnFFuBIPbDqWv7Lj
xWEXVzo7cKZ2rlY5BLRKv/Oe3OxhVoAk1HoipGQE+r0Pa9dTA5TDrNvI0eR7
88/ESkq28FNL3+Me2oCttlGYyaZYkBe2Cya0zJv8Zf/vjYwrTtkavR++Hbf4
+2io4QZMQWuk9PJucPOxDkCsz3dxlzsYEDr2Bz36zrIfngYnCzFRZp/lfRJv
Ev7KYQ3gn8Sjm5XiROWlRAR1NRIT+FgzmuOFooNRlU9M/VhCAsRb1nGLYGNb
Ku/rybGmQTzw+y65NiN2un/EuVgzpleblPDbVgmrj/UdUV1dzv1b38ZoUaBV
2blNrDAfPkx4p0nmyHojH5jgZlnKKh71UQ8j/m4ptEdTY8p5MZ2dd5OjH+es
/ojIKyde0sG8LE17/wBFe0gHlm5k5B6Pyh39tQ5T7fTRkD3uaGlWSog3Fivl
Kom1cziIuXLGVltWh21tO6oW8TksG5aLDYJvRYTG61SAhNwEJYpxUChpeKFI
Clfox1TyaBdAu4fKv1+aHyoxaJ3863kIgeOFoelwiXhtiokWjvsfMWWV+mas
XLNDId8jWpHb9wgPO8l5ARjILWiQh9KU75QU1hzmeVW+lt5N4JfsngNLvOT/
fUVROpxQXwKWDHd93igiWOzXmykRMTuMh+FstGaSEWKK3uAr04Yr90lTQTHW
LCjXGFi71ur8mUVoq/RlDxNXVnRfP8DOl1SfUwkvWVis4ImIdPfZssvl/5nl
PcupV5zAxmlEgyHkrXWuPvGRM+Xfy0rlJ5PxzifUSekRZn+AkLccIrzoUn+H
yI5jbpuoSvfZOTjMof7y7GJ1QUbJvEmAFAvcNGvBQextdeBR7IPownMgXBIa
tq8Qp7c+oAJbqs2t+cLlWaOFClYbNlJo07Mg573yPa1iRRxj5yf09hJG80BW
h+FOZhuxMJq2ojRtcYo8bdqdykVZ0ASjxSCzSA5PGRqh+QF0e2/rFl5tE6O5
mwbC7V5upGOpKTnD3Zly2mdyx10ZPK1D7Z8iT0VCupHR5xYWDYoa6NiJg6qs
0eUDA0zKSco8yfO+8n3m7xVmOvvTG+oQjLoOCS8PNjMSzMKrsLY1IrYDGZrA
bGqhoWLWCKHgKhjxH2IZsAwUIvxklhsWGE4PqkpGGhZNarr78kVOR41KFaul
QtHzTNacJ03eJ2hfbhvYvs4YWh8n4egOIPzue0a3NWwTEvLWLFNEogeo9l7k
Fd6jTJZeyH4qnZVAaELejVIlw3S55xfrk5ND6YoJwKaGcfJ3RXhoBbmfusal
nu3dPKn4QBwQoLedLl07lfFIapNPb9g1mpR4iwzacBWu0XpjB4TwjX2YbFLo
gjD9LN5OWZc9x9rSsNuWXA9G5lA2V+qqM7mwTY3JBg3GY/TFjxirt7OJqvBg
dM9pHk6dcTWsPZhMS9c+smAZhIvH3C+3VPA22+XsMnE76HUopAk3RqDROl8Y
GtSyRxXR1KqxO/cW6LYJPgJgeMUXroSVPI+c13fA9Q8KRwYGLxW7Te9dXk1L
fO/aWYuAmqZIZ6jWyyI+dlvobKESIawejZTR+X8sAqD3ZCfzwXM/80mPzPkH
c1eg4ivTCJCadh+mjG3hbCrGyzGLfNH4idcctqVH6a5rk7TybZoYC52uErnj
mwL2StR0Plt5WgznoPRDeQ7Bw2nWT3qVAQN6etcu5cpJgIZ4T4OeMOoDKX1L
G503e/RLei2xBqwSaqTHRVF3LeXzMW2YzBraBOgwOwwbqSTn+KMHrE874916
eme7gz2mz6OgKIqn/VfwsBCz1gQHJWagGu12GaUQ/F5iseO9c1Cn+BphR2XR
gDQSgQdDifAAfTQF0w2P6uDO3amxrMOZNdIMOcaWhd23OreV95pTcvkz/cXC
R4wR4E0bLQkXAPxJYwA7wpZYDBotC59xu9ZXpVwVJv2LfD3NTDMyBLBVv5t+
ZvxX1OvVGiMy2qF7A5QpSJkyam+6IobgGkSHwD8hkt5wVd/RkNbk6QIBzRkL
XrrhoQBvT/mnU1SwhtJQiNYX9qjdAdrJa8DzF0RB3bCFF9wPPXaTQj4K85xB
gkGX9BHU8ry7B+I+A3fVodT7zn0jUxrNrqq5q+smVxD5Gm2o4oKmkRYnwEUA
ww2pa8B0+nXxFcd/+i6nqux/JNvtkCeGI5yuMvbVOz90CnXSVODK5psl7yU8
S6R6FSPcvizKlCItdYSSjzwGIIbIy9MwEsuqxLIknjiEkcNfi/pffqhcgE45
34S/zrGURGFEZEVpbTxjs//iF2UQYSpXny7UOzu4YRte1ELtoY1ML8j4Y2j1
mD0Id+2UxJBvNno0dLZowTK21bLO2aeAk7vP+va74Fllw7nc4nstQlS0J/Rv
lJC+TJ1q7+ntk8nvh7dAeGp+JJs1AXGB+t5cnSRrlFf2BI8Yqn9LjYpSk13E
EfInSElPgoRZBQT6ECVJU8+wAz8AUmWjhPSEXfs84LXDy9U1b21Ccplz0sk0
RH8lRmr0dfDt4vZCO+NFK2dFQ0/+zX1jfrFCr0HU1c7po0Badw8jBAnXJkA9
AJhoCNPMvtQoiMw/Ol7s7xkyCuPgUPTxDZjebjwxeojoLKVAwqAeZpQh/WUR
wnIRAMS0O+HAuKdxp6sjEu0AYbvOG7olcXfWmTZQXHmBcfW+581Ecarz2w40
KxGGj8q7xuOrwY64v77O4Y7xKrWp1rOz2H33KwhsbC5n/hLem0b9Fa+5BQ8H
dcrVEeclOpEI/ih1RNnCitFuLqMQLq1YHnGuG6ExDFciEmgxTUdZwHMnQi/5
hZkQ7pGqP0iAF1KaiU7cFPdz0mvo2rpMNp9+Zc4bmLlan/JHvOzys+EiB7c/
qMkthwy7oKgJngs4LxygpfXl45bCatewc5GsLRj/b12udcRAE+0rdvR2mDzR
qOpw50c+WsAM3vxlXUGIp/sCHKiorOG/7oUo4s4RQVrLP7u362cTJW1i78KA
2uKVoPSoteb4aM1WYkfQleQxjdXTxa418Js/YwVROtVcsZEm1FYHW3qB+WMh
ONImjyq018P4Ay1HnbSvaTNxbVvQNSGuGeh49FPFA+DwIemeArFtqM1FpoHg
54MjA0ml55qDcazrOFVjGnDiK9VB1mDHeFz0H8/pZ0TzFJQjPsO7

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q77kCzkJRt5T4Dhw86+8zKNmkFlBGX5dbKk8DYPE8NsDU5xCCMCWheaNTmmxIHHrevbNDUTcZFURbQznuvvvqQFfjKFA+Y5x7HG9OhJaOgYdQEK59RHnZ8w1WcuiqPbDZQs7ez7AaTltKhICkIWt15h+Ru3FUAQpBL/VweG3w+CpkC0M6o7gngtRSmQW8g01d0ktZL1XYBJIj9MluekYktxhlrVfoVw37RQu1MaGBPKWb+HBYtvzXYDDIBVmNQTKwFrZDa4OOqehC4kqb2ahk2Tjn5YrMxm+DiUNYDDT98RZPSBmk7C60vHdh5CWGBykmX2cbfq4wflQtF3v4l2mAZOXyaWYImu7ltvm72VECh7apU/uitCVQ3R0HV//Tn6qeptbL7NLD58cfFlYj6d33SRd9SvGcrB6gx9i3OgNM07DXfkosYWVrdzWSczg1gQODYVg97u6fEnAWGMLxMdmg7jWpe6G1M7nfeUBCJ6inHU2JJwRBoJUoetFA25Y6FEVbQCeRMzClT0HFQ1MDtwMKErHsxFIdeuM9fwWbFKf9/Osmg9lbw3zaSfnRqX1hQpgNyt4Z5sgy71/kwrWChBGeKMjrOOGtVWAmlNEit3wLnIafvU7/t76QYTVf6Z+BihSP8dZh+ila/5ZSVy68z68Qa6dcOX8VuzfkHJX09Q/MUfDVje3HZ5Xv8AU7CvzopsuyELaiKYeRRI8SBPN9dagBDoGIcrjGavnG/DC/cs7aYpmr0YyXekmiubjdZSm0mzDwJLzt0cHHENFBdn2CGw6Ffa"
`endif