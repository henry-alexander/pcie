// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


 
module system_intel_pcie_gts_0_pldif_hal_2100_7x7kbai
  #(
    parameter ch_pldif_l_tx_en_atom                      = "FALSE"                           ,
    parameter ch_pldif_l_rx_en_atom                      = "FALSE"                           ,
    parameter ch_pldif_l_duplex_mode_atom                = "DUPLEX_MODE_DUPLEX"             ,
    parameter ch_pldif_l_tx_fifo_mode_atom               = "TX_FIFO_MODE_PHASE_COMP"        ,
    parameter ch_pldif_l_tx_fifo_width_atom              = "TX_FIFO_WIDTH_DOUBLE_WIDTH"     ,
    parameter ch_pldif_l_rx_fifo_mode_atom               = "RX_FIFO_MODE_PHASE_COMP"        ,
    parameter ch_pldif_l_rx_fifo_width_atom              = "RX_FIFO_WIDTH_DOUBLE_WIDTH"     ,
    parameter ch_pldif_l_tx_clkout1_divider_atom         = "TX_CLKOUT1_DIVIDER_DIV1"         ,
    parameter ch_pldif_l_tx_clkout2_divider_atom         = "TX_CLKOUT2_DIVIDER_DIV1"         ,
    parameter ch_pldif_l_rx_clkout1_divider_atom         = "RX_CLKOUT1_DIVIDER_DIV1"         ,
    parameter ch_pldif_l_rx_clkout2_divider_atom         = "RX_CLKOUT2_DIVIDER_DIV1"         ,
    parameter ch_pldif_l_dr_enabled_atom                 = "DR_ENABLED_DR_ENABLED"          ,
    parameter ch_pldif_l_ptp_enable_atom                 = "PTP_ENABLE_ENABLE"               ,
    parameter ch_pldif_l_tx_user1_clk_dynamic_mux_atom   = "TX_USER1_CLK_DYNAMIC_MUX_UNUSED" ,
    parameter ch_pldif_l_tx_user2_clk_dynamic_mux_atom   = "TX_USER2_CLK_DYNAMIC_MUX_UNUSED" ,
    parameter ch_pldif_l_rx_user1_clk_dynamic_mux_atom   = "RX_USER1_CLK_DYNAMIC_MUX_UNUSED" ,
    parameter ch_pldif_l_rx_user2_clk_dynamic_mux_atom   = "RX_USER2_CLK_DYNAMIC_MUX_UNUSED" ,
    parameter ch_pldif_l_sup_mode_atom                   = "SUP_MODE_USER_MODE"             ,
    parameter ch_pldif_l_tx_mac_en_atom                  = "FALSE"                          ,
    parameter ch_pldif_l_rx_dyn_mux_atom                 = "RX_DYN_MUX_UNUSED"               ,
    parameter ch_pldif_l_tx_bond_location_atom           = "TX_BOND_LOCATION_FIRST"          ,
    parameter ch_pldif_l_rx_bond_location_atom           = "RX_BOND_LOCATION_FIRST"          ,
    parameter ch_pldif_l_ehip_lb_tx_rx_atom              = "EHIP_LB_TX_RX_ENABLE"            ,
    parameter ch_pldif_l_ehip_lb_txmac_rx_atom           = "EHIP_LB_TXMAC_RX_ENABLE"         ,
    parameter ch_pldif_l_rx_pmadir_singlewidth_en_atom   = "RX_PMADIR_SINGLEWIDTH_EN_ENABLE" ,
    parameter ch_pldif_l_tx_pmadir_singlewidth_en_atom   = "TX_PMADIR_SINGLEWIDTH_EN_ENABLE" ,
    parameter ch_pldif_l_ehip_lb_txpcs_rx_atom           = "EHIP_LB_TXPCS_RX_ENABLE"         ,
    parameter ch_pcs_l_tx_bond_size_atom                 = "TX_BOND_SIZE_UNUSED"             ,
    parameter ch_pcs_l_rx_bond_size_atom                 = "RX_BOND_SIZE_UNUSED"             ,    
    parameter ch_pldif_l_pld_channel_identifier_atom     = "PLD_CHANNEL_IDENTIFIER_GENERIC"  ,   
    parameter ch_pldif_rx_fifo_wr_clk_hz_atom            = 36'd0                             ,   
    parameter ch_pldif_tx_fifo_rd_clk_hz_atom            = 36'd0                             ,   
    parameter ch_vc_rx_pldif_wm_en_atom                  = "VC_RX_PLDIF_WM_EN_ENABLE"           ,    
    parameter ch_pldif_l_stmux_tx_demux_sel              = "SEL_ETH"                            ,
    parameter ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel    = "SEL_ETH_OR_PTP"                     ,
    parameter ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel    = "SEL_ETH_OR_PTP"                     ,
    parameter ch_pldif_l_stmux_rx_mux_sel                = "SEL_ETH"                            ,
    parameter ch_l_xcvr_rx_preloaded_hardware_configs    = "NONE"                               ,
    parameter ch_l_xcvr_tx_preloaded_hardware_configs    = "NONE"
)
(
    input    [79:0]  i_hio_txdata                         ,      
    input    [9:0]   i_hio_txdata_extra                   ,     
    input            i_hio_txdata_fifo_wr_en              ,     
    output           o_hio_txdata_fifo_wr_empty           ,     
    output           o_hio_txdata_fifo_wr_pempty          ,     
    output           o_hio_txdata_fifo_wr_full            ,     
    output           o_hio_txdata_fifo_wr_pfull           ,     
    output   [79:0]  o_hio_rxdata                         ,     
    output   [9:0]   o_hio_rxdata_extra                   ,     
    output           o_hio_rxdata_fifo_rd_empty           ,     
    output           o_hio_rxdata_fifo_rd_pempty          ,     
    output           o_hio_rxdata_fifo_rd_full            , 
    output           o_hio_rxdata_fifo_rd_pfull           , 
    input            i_hio_rxdata_fifo_rd_en              ,     
    input            i_hio_ptp_rst_n                      ,
    input            i_hio_ehip_rx_rst_n                  ,
    input            i_hio_ehip_tx_rst_n                  ,
    input            i_hio_ehip_signal_ok                 ,
    input            i_hio_sfreeze_2_r03f_rx_mac_srfz_n   ,              
    input            i_hio_sfreeze_3_c2f_tx_deskew_srfz_n,                    
    input            i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n   ,           
    output           o_hio_rstepcs_rx_pcs_fully_aligned   ,     
    input            i_hio_rstfec_fec_rx_rst_n            ,   
    input            i_hio_rstfec_fec_tx_rst_n            ,   
    input            i_hio_rstfec_fec_csr_ret             ,     
    output           o_hio_rstfec_fec_rx_rdy_n            ,   
    input            i_hio_rstfec_rx_fec_sfrz_n           ,
    input            i_hio_rstfec_tx_fec_sfrz_n           , 
    input            i_hio_rstxcvrif_xcvrif_rx_rst_n      ,    
    input            i_hio_rstxcvrif_xcvrif_tx_rst_n      ,    
    input            i_hio_rstxcvrif_xcvrif_signal_ok     ,       
    input            i_hio_rstxcvrif_rx_xcvrif_sfrz_n     ,
    input            i_hio_rstxcvrif_tx_xcvrif_sfrz_n     ,
    input            i_hio_rst_pld_clrhip                 ,     
    input            i_hio_rst_pld_clrpcs                 ,     
    input            i_hio_rst_pld_perstn                 ,     
    input            i_hio_rst_pld_ready                  ,     
    input            i_hio_rst_pld_adapter_rx_pld_rst_n   ,     
    input            i_hio_rst_pld_adapter_tx_pld_rst_n   ,     
    input            i_hio_rst_ux_rx_pma_rst_n            ,     
    input            i_hio_rst_ux_rx_sfrz                 ,     
    input            i_hio_rst_ux_tx_pma_rst_n            ,     
    output           o_hio_rst_flux0_cpi_cmn_busy         ,     
    output           o_hio_rst_oflux_rx_srds_rdy          ,     
    output           o_hio_rst_ux_all_synthlockstatus     ,     
    output           o_hio_rst_ux_octl_pcs_rxstatus       ,     
    output           o_hio_rst_ux_octl_pcs_txstatus       ,     
    output           o_hio_rst_ux_rxcdrlock2data          ,     
    output           o_hio_rst_ux_rxcdrlockstatus         ,     
/*    output           o_ss_ptp_rst_n                       ,   */
    output           o_ss_ehip_rx_rst_n                   ,
    output           o_ss_ehip_tx_rst_n                   ,
    output           o_ss_ehip_signal_ok                  ,
    output           o_ss_sfreeze_2_r03f_rx_mac_srfz_n    ,     
    output           o_ss_sfreeze_3_c2f_tx_deskew_srfz_n ,                      
    input            i_ss_rstepcs_rx_pcs_fully_aligned    ,     
    output           o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n    ,              
    output           o_ss_rstfec_fec_rx_rst_n             ,   
    output           o_ss_rstfec_fec_tx_rst_n             ,   
    output           o_ss_rstfec_fec_csr_ret              ,     
    input            i_ss_rstfec_fec_rx_rdy_n             ,   
    output           o_ss_rstfec_rx_fec_sfrz_n            ,
    output           o_ss_rstfec_tx_fec_sfrz_n            ,
    output           o_ss_rstxcvrif_xcvrif_rx_rst_n       ,    
    output           o_ss_rstxcvrif_xcvrif_tx_rst_n       ,    
    output           o_ss_rstxcvrif_xcvrif_signal_ok      ,       
    output           o_ss_rstxcvrif_rx_xcvrif_sfrz_n      ,
    output           o_ss_rstxcvrif_tx_xcvrif_sfrz_n      ,
//    output           o_ss_pcie_rst_pld_clrhip             ,     
//    output           o_ss_pcie_rst_pld_clrpcs             ,     
//    output           o_ss_pcie_rst_pld_perstn             ,     
    output           o_ss_rst_ux_rx_pma_rst_n             ,     
    output           o_ss_rst_ux_rx_sfrz                  ,     
    output           o_ss_rst_ux_tx_pma_rst_n             ,     
    input            i_ss_rst_flux0_cpi_cmn_busy          ,     
    input            i_ss_rst_oflux_rx_srds_rdy           ,     
    input            i_ss_rst_ux_all_synthlockstatus      ,     
    input            i_ss_rst_ux_octl_pcs_rxstatus        ,     
    input            i_ss_rst_ux_octl_pcs_txstatus        ,     
    input            i_ss_rst_ux_rxcdrlock2data           ,     
    input            i_ss_rst_ux_rxcdrlockstatus          ,     
    input            i_hio_pld_reset_clk_row              ,     
    input    [11:0]  i_ss_eth_fec_rx_async                ,     
    input            i_ss_eth_fec_rx_direct               ,     
    output   [6:0 ]  o_ss_eth_fec_tx_async                ,     
    output           o_ss_eth_fec_tx_direct               ,     
    input    [13:0]  i_ss_eth_mac_rx_async                ,     
    input            i_ss_eth_mac_rx_direct               ,     
    output   [13:0]  o_ss_eth_mac_tx_async                ,     
    output           o_ss_eth_mac_tx_direct               ,     
    input    [13:0]  i_ss_eth_pcs_rx_async                ,     
    input            i_ss_eth_pcs_rx_direct               ,     
    output   [7:0 ]  o_ss_eth_pcs_tx_async                ,     
    output           o_ss_eth_pcs_tx_direct               ,     
    input    [13:0]  i_ss_eth_xcvrif_rx_async             ,     
    input            i_ss_eth_xcvrif_rx_direct            ,     
    output   [6:0 ]  o_ss_eth_xcvrif_tx_async             ,     
    output           o_ss_eth_xcvrif_tx_direct            ,     
    input    [87:0]  i_ss_pcie_ctrl_rx_async              ,     
    input    [7:0 ]  i_ss_pcie_ctrl_rx_direct             ,     
//    output   [87:0]  o_ss_pcie_ctrl_tx_async              ,     
//    output   [7:0 ]  o_ss_pcie_ctrl_tx_direct             ,     
    output   [79:0]  o_ss_uxquad_async                    ,
    output   [79:0]  o_ss_uxquad_async_pcie_mux           ,                   
    input    [49:0]  i_ss_uxquad_async                    , 
    input    [79:0]  i_hio_uxquad_async                   ,
    input    [79:0]  i_hio_uxquad_async_pcie_mux          ,                    
    output   [49:0]  o_hio_uxquad_async                   ,  
    input    [99:0]  i_hio_txdata_async                   ,     
    input    [9:0 ]  i_hio_txdata_direct                  ,     
    output   [99:0]  o_hio_rxdata_async                   ,     
    output   [9:0 ]  o_hio_rxdata_direct                  ,     
    output   [31:0]  o_hio_lavmm_rdata                    ,     
    output           o_hio_lavmm_rdata_valid              ,     
    output           o_hio_lavmm_waitreq                  ,     
    input    [20:0]  i_hio_lavmm_addr                     ,     
    input    [3:0 ]  i_hio_lavmm_be                       ,     
    input            i_hio_lavmm_clk                      ,     
    input            i_hio_lavmm_read                     ,     
    input            i_hio_lavmm_rstn                     ,     
    input    [31:0]  i_hio_lavmm_wdata                    ,     
    input            i_hio_lavmm_write                    ,     
    input    [31:0]  i_ss_lavmm_pcie_rdata                ,     
    input            i_ss_lavmm_pcie_rdata_valid          ,     
    input            i_ss_lavmm_pcie_waitreq              ,     
    output   [16:0]  o_ss_lavmm_pcie_addr                 ,     
    output   [3:0 ]  o_ss_lavmm_pcie_be                   ,     
    output           o_ss_lavmm_pcie_clk                  ,     
    output           o_ss_lavmm_pcie_read                 ,     
    output           o_ss_lavmm_pcie_rstn                 ,     
    output   [31:0]  o_ss_lavmm_pcie_wdata                ,     
    output           o_ss_lavmm_pcie_write                ,  
    
    output   [2:0 ]  k_user_rx_clk1_c0c1c2_sel            ,     
    output   [2:0 ]  k_user_rx_clk2_c0c1c2_sel            ,     
    output   [2:0 ]  k_user_tx_clk1_c0c1c2_sel            ,     
    output   [2:0 ]  k_user_tx_clk2_c0c1c2_sel            ,     
    input            i_ss_user_rx_clk1_clk                ,     
    input            i_ss_user_rx_clk2_clk                ,     
    input            i_ss_user_tx_clk1_clk                ,     
    input            i_ss_user_tx_clk2_clk                ,     
    
    output           o_hio_user_rx_clk1_clk               ,     
    output           o_hio_user_rx_clk2_clk               ,     
    output           o_hio_user_tx_clk1_clk               ,     
    output           o_hio_user_tx_clk2_clk               ,     
    input            i_ux_chnl_refclk_mux                 ,     
    output           o_hio_ux_chnl_refclk_mux             ,     
/*     input            i_ss_tx_fifo_clk                     ,     
    input            i_ss_rx_fifo_clk                     ,  */    
    input            i_hio_pld_rx_clk_in_row_clk          ,     
    input            i_hio_pld_tx_clk_in_row_clk          ,     
    input            i_hio_det_lat_rx_dl_clk              ,       
    input            i_hio_det_lat_rx_mux_select          ,       
    input            i_hio_det_lat_rx_sclk_flop           ,       
    input            i_hio_det_lat_rx_sclk_gen_clk        ,       
    input            i_hio_det_lat_rx_trig_flop           ,       
    input            i_hio_det_lat_sampling_clk           ,       
    input            i_hio_det_lat_tx_dl_clk              ,       
    input            i_hio_det_lat_tx_mux_select          ,       
    input            i_hio_det_lat_tx_sclk_flop           ,       
    input            i_hio_det_lat_tx_sclk_gen_clk        ,       
    input            i_hio_det_lat_tx_trig_flop           ,       
    output           o_hio_det_lat_rx_async_dl_sync       ,       
    output           o_hio_det_lat_rx_async_pulse         ,       
    output           o_hio_det_lat_rx_async_sample_sync   ,       
    output           o_hio_det_lat_rx_sclk_sample_sync    ,       
    output           o_hio_det_lat_rx_trig_sample_sync    ,       
    output           o_hio_det_lat_tx_async_dl_sync       ,       
    output           o_hio_det_lat_tx_async_pulse         ,       
    output           o_hio_det_lat_tx_async_sample_sync   ,       
    output           o_hio_det_lat_tx_sclk_sample_sync    ,       
    output           o_hio_det_lat_tx_trig_sample_sync    ,       
    output           o_hio_xcvrif_rx_latency_pulse        ,
    output           o_hio_xcvrif_tx_latency_pulse        ,
    output           o_ss_det_lat_rx_sclk_clk             ,       
    output           o_ss_det_lat_rx_sclk_sync            ,       
    output           o_ss_det_lat_tx_sclk_clk             ,       
    output           o_ss_det_lat_tx_sclk_sync            ,       
    input            i_ss_det_lat_rx_async_pulse          ,       
    input            i_ss_det_lat_tx_async_pulse          ,       
    input            i_ss_xcvrif_rx_latency_pulse         ,
    input            i_ss_xcvrif_tx_latency_pulse         ,
    input            i_ux_tx_ch_ptr_smpl                  ,
    output           o_hio_ux_tx_ch_ptr_smpl              ,
    //deskew signals////                                  
    input            i_deskew_rx_ch_clk                   ,
    input            i_deskew_tx_ch_clk                   ,
    output           o_marker_found                       ,
    input            i_marker_found_up                    ,
    input            i_marker_found_dn                    ,
/*     output   [2:0]   o_deskew_rx_source_sel               ,
    input    [42:0]  i_ch_muxed_rx_data                   , */
    output   [42:0]  o_ch_pld_tx_deskewed_data            ,
    output   [8:0]   o_ch_ptp_tx_deskewed_data            ,
    input    [7:0]   i_ch_ptp_rx_data                     ,
    input            i_ch_tx_mac_ready                    ,
    input            i_ch_rx_mac_inframe                  ,
    output           o_ch_tx_mac_valid                    ,
    input            i_ptp_rx_dsk_marker                  ,
    input            i_ptp_mas_wm                         ,
    input    [42:0]  i_tx_pcs_data                        ,
    input    [42:0]  i_tx_mac_data                        ,
    //lavmm signals////                                   
    output   [19:0]  o_lavmm_xcvrif_addr                  ,
    output   [3:0]   o_lavmm_xcvrif_be                    ,
    output           o_lavmm_xcvrif_clk                   ,
    output           o_lavmm_xcvrif_read                  ,
    output           o_lavmm_xcvrif_rstn                  ,
    output   [31:0]  o_lavmm_xcvrif_wdata                 ,
    output           o_lavmm_xcvrif_write                 ,
    input    [31:0]  i_lavmm_xcvrif_rdata                 ,
    input            i_lavmm_xcvrif_rdata_valid           ,
    input            i_lavmm_xcvrif_waitreq               ,
    output   [19:0]  o_lavmm_emac_addr                    ,
    output   [3:0]   o_lavmm_emac_be                      ,
    output           o_lavmm_emac_clk                     ,
    output           o_lavmm_emac_read                    ,
    output           o_lavmm_emac_rstn                    ,
    output   [31:0]  o_lavmm_emac_wdata                   ,
    output           o_lavmm_emac_write                   ,
    input    [31:0]  i_lavmm_emac_rdata                   ,
    input            i_lavmm_emac_rdata_valid             ,
    input            i_lavmm_emac_waitreq                 ,
    output   [19:0]  o_lavmm_epcs_addr                    ,
    output   [3:0]   o_lavmm_epcs_be                      ,
    output           o_lavmm_epcs_clk                     ,
    output           o_lavmm_epcs_read                    ,
    output           o_lavmm_epcs_rstn                    ,
    output   [31:0]  o_lavmm_epcs_wdata                   ,
    output           o_lavmm_epcs_write                   ,
    input    [31:0]  i_lavmm_epcs_rdata                   ,
    input            i_lavmm_epcs_rdata_valid             ,
    input            i_lavmm_epcs_waitreq                 ,
    output   [19:0]  o_lavmm_fec_addr                     ,
    output   [3:0]   o_lavmm_fec_be                       ,
    output           o_lavmm_fec_clk                      ,
    output           o_lavmm_fec_read                     ,
    output           o_lavmm_fec_rstn                     ,
    output   [31:0]  o_lavmm_fec_wdata                    ,
    output           o_lavmm_fec_write                    ,
    input    [31:0]  i_lavmm_fec_rdata                    ,
    input            i_lavmm_fec_rdata_valid              ,
    input            i_lavmm_fec_waitreq                  ,
/*    output   [19:0]  o_lavmm_ptp_addr                     ,
    output   [3:0]   o_lavmm_ptp_be                       ,
    output           o_lavmm_ptp_clk                      ,
    output           o_lavmm_ptp_read                     ,
    output           o_lavmm_ptp_rstn                     ,
    output   [31:0]  o_lavmm_ptp_wdata                    ,
    output           o_lavmm_ptp_write                    ,
    input    [31:0]  i_lavmm_ptp_rdata                    ,
    input            i_lavmm_ptp_rdata_valid              ,
    input            i_lavmm_ptp_waitreq                  , */
    output   [19:0]  o_lavmm_ux_addr                      ,
    output   [3:0]   o_lavmm_ux_be                        ,
    output           o_lavmm_ux_clk                       ,
    output           o_lavmm_ux_read                      ,
    output           o_lavmm_ux_rstn                      ,
    output   [31:0]  o_lavmm_ux_wdata                     ,
    output           o_lavmm_ux_write                     ,
    input    [31:0]  i_lavmm_ux_rdata                     ,
    input            i_lavmm_ux_rdata_valid               ,
    input            i_lavmm_ux_waitreq                   ,
    
    //missed out interfaces
    input    [10:0]  i_ptp_tx_data,
    output   [9:0]   o_ch_ptp_rx_data,

    //adding interfaces for muxes
    output   [79:0]  sm_pld_tx_demux_0_o_pcie           ,
/*     input            sm_hssi_pld_chnl_user_mux_0_i_c0   ,
    input            sm_hssi_pld_chnl_user_mux_2_i_c0   ,
    input            sm_hssi_pld_chnl_user_mux_3_i_c0   ,
    input            sm_hssi_pld_chnl_user_mux_1_i_c0   ,
    input            sm_hssi_pld_chnl_user_mux_0_i_c1   ,
    input            sm_hssi_pld_chnl_user_mux_2_i_c1   ,
    input            sm_hssi_pld_chnl_user_mux_3_i_c1   ,
    input            sm_hssi_pld_chnl_user_mux_1_i_c1   ,
    input            sm_hssi_pld_chnl_user_mux_0_i_c2   ,
    input            sm_hssi_pld_chnl_user_mux_2_i_c2   ,
    input            sm_hssi_pld_chnl_user_mux_3_i_c2   ,
    input            sm_hssi_pld_chnl_user_mux_1_i_c2   , */
    input            sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp ,
    input            sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp ,
    /* input    [42:0]  sm_deskew_rx_mux_0_i_ethmac                        ,
    input    [42:0]  sm_deskew_rx_mux_0_i_ethpcs                        ,
    input    [42:0]  sm_deskew_rx_mux_0_i_fec   */                         
    input    [79:0]  sm_pld_rx_mux_0_i_pcie                             ,
    input            sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie       ,
    input            sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie       ,
    input    [79:0]  sm_pld_rx_mux_0_i_pcie_bond                        ,
    input            sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top   ,
    input            sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top   ,
/*     input            sm_hssi_pld_chnl_user_mux_0_i_ux,
    input            sm_hssi_pld_chnl_user_mux_2_i_ux,
    input            sm_hssi_pld_chnl_user_mux_3_i_ux,
    input            sm_hssi_pld_chnl_user_mux_1_i_ux,
    input    [42:0]  sm_deskew_rx_mux_0_i_xcvrif */
    
    //r9 additions
    input [42:0]     i_ch_muxed_rx_data,
    output [2:0]     o_deskew_rx_source_sel
                
);  

pldif_hal_coreip 
#(
    .ch_pldif_l_tx_en_atom                     (ch_pldif_l_tx_en_atom                   ),
    .ch_pldif_l_rx_en_atom                     (ch_pldif_l_rx_en_atom                   ),
    .ch_pldif_l_duplex_mode_atom               (ch_pldif_l_duplex_mode_atom             ),
    .ch_pldif_l_tx_fifo_mode_atom              (ch_pldif_l_tx_fifo_mode_atom            ),
    .ch_pldif_l_tx_fifo_width_atom             (ch_pldif_l_tx_fifo_width_atom           ),
    .ch_pldif_l_rx_fifo_mode_atom              (ch_pldif_l_rx_fifo_mode_atom            ),
    .ch_pldif_l_rx_fifo_width_atom             (ch_pldif_l_rx_fifo_width_atom           ),
    .ch_pldif_l_tx_clkout1_divider_atom        (ch_pldif_l_tx_clkout1_divider_atom      ),
    .ch_pldif_l_tx_clkout2_divider_atom        (ch_pldif_l_tx_clkout2_divider_atom      ),
    .ch_pldif_l_rx_clkout1_divider_atom        (ch_pldif_l_rx_clkout1_divider_atom      ),
    .ch_pldif_l_rx_clkout2_divider_atom        (ch_pldif_l_rx_clkout2_divider_atom      ),
    .ch_pldif_l_dr_enabled_atom                (ch_pldif_l_dr_enabled_atom              ),
    .ch_pldif_l_ptp_enable_atom                (ch_pldif_l_ptp_enable_atom              ),
    .ch_pldif_l_tx_user1_clk_dynamic_mux_atom  (ch_pldif_l_tx_user1_clk_dynamic_mux_atom),
    .ch_pldif_l_tx_user2_clk_dynamic_mux_atom  (ch_pldif_l_tx_user2_clk_dynamic_mux_atom),
    .ch_pldif_l_rx_user1_clk_dynamic_mux_atom  (ch_pldif_l_rx_user1_clk_dynamic_mux_atom),
    .ch_pldif_l_rx_user2_clk_dynamic_mux_atom  (ch_pldif_l_rx_user2_clk_dynamic_mux_atom),
    .ch_pldif_l_sup_mode_atom                  (ch_pldif_l_sup_mode_atom                ),
    .ch_pldif_l_tx_mac_en_atom                 (ch_pldif_l_tx_mac_en_atom               ),
    .ch_pldif_l_rx_dyn_mux_atom                (ch_pldif_l_rx_dyn_mux_atom              ),
    .ch_pldif_l_tx_bond_location_atom          (ch_pldif_l_tx_bond_location_atom        ),
    .ch_pldif_l_rx_bond_location_atom          (ch_pldif_l_rx_bond_location_atom        ),
    .ch_pldif_l_ehip_lb_tx_rx_atom             (ch_pldif_l_ehip_lb_tx_rx_atom           ),
    .ch_pldif_l_ehip_lb_txmac_rx_atom          (ch_pldif_l_ehip_lb_txmac_rx_atom        ),
    .ch_pldif_l_rx_pmadir_singlewidth_en_atom  (ch_pldif_l_rx_pmadir_singlewidth_en_atom),
    .ch_pldif_l_tx_pmadir_singlewidth_en_atom  (ch_pldif_l_tx_pmadir_singlewidth_en_atom),
    .ch_pldif_l_ehip_lb_txpcs_rx_atom          (ch_pldif_l_ehip_lb_txpcs_rx_atom        ),
    .ch_pcs_l_tx_bond_size_atom                (ch_pcs_l_tx_bond_size_atom             ),
    .ch_pcs_l_rx_bond_size_atom                (ch_pcs_l_rx_bond_size_atom             ),
    .ch_pldif_l_pld_channel_identifier_atom    (ch_pldif_l_pld_channel_identifier_atom  ),
    .ch_pldif_rx_fifo_wr_clk_hz_atom           (ch_pldif_rx_fifo_wr_clk_hz_atom  ),
    .ch_pldif_tx_fifo_rd_clk_hz_atom           (ch_pldif_tx_fifo_rd_clk_hz_atom  ),
    .ch_vc_rx_pldif_wm_en_atom                 (ch_vc_rx_pldif_wm_en_atom  ),
    .ch_pldif_l_stmux_tx_demux_sel             (ch_pldif_l_stmux_tx_demux_sel           ),
    .ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel   (ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel ),
    .ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel   (ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel ),  
    .ch_pldif_l_stmux_rx_mux_sel               (ch_pldif_l_stmux_rx_mux_sel             ),
    .ch_l_xcvr_rx_preloaded_hardware_configs   (ch_l_xcvr_rx_preloaded_hardware_configs ),
    .ch_l_xcvr_tx_preloaded_hardware_configs   (ch_l_xcvr_tx_preloaded_hardware_configs )

)
pldif_hal_coreip_inst (
    .i_hio_txdata                           (i_hio_txdata                           ),         
    .i_hio_txdata_extra                     (i_hio_txdata_extra                     ),
    .i_hio_txdata_fifo_wr_en                (i_hio_txdata_fifo_wr_en                ),
    .o_hio_txdata_fifo_wr_empty             (o_hio_txdata_fifo_wr_empty             ),
    .o_hio_txdata_fifo_wr_pempty            (o_hio_txdata_fifo_wr_pempty            ),
    .o_hio_txdata_fifo_wr_full              (o_hio_txdata_fifo_wr_full              ),
    .o_hio_txdata_fifo_wr_pfull             (o_hio_txdata_fifo_wr_pfull             ),
    .o_hio_rxdata                           (o_hio_rxdata                           ),
    .o_hio_rxdata_extra                     (o_hio_rxdata_extra                     ),
    .o_hio_rxdata_fifo_rd_empty             (o_hio_rxdata_fifo_rd_empty             ),
    .o_hio_rxdata_fifo_rd_pempty            (o_hio_rxdata_fifo_rd_pempty            ),
    .o_hio_rxdata_fifo_rd_full              (o_hio_rxdata_fifo_rd_full              ),
    .o_hio_rxdata_fifo_rd_pfull             (o_hio_rxdata_fifo_rd_pfull             ),
    .i_hio_rxdata_fifo_rd_en                (i_hio_rxdata_fifo_rd_en                ),
    .i_hio_ptp_rst_n                        (i_hio_ptp_rst_n                        ),
    .i_hio_ehip_rx_rst_n                    (i_hio_ehip_rx_rst_n                    ),
    .i_hio_ehip_tx_rst_n                    (i_hio_ehip_tx_rst_n                    ),
    .i_hio_ehip_signal_ok                   (i_hio_ehip_signal_ok                   ),
    .i_hio_sfreeze_2_r03f_rx_mac_srfz_n     (i_hio_sfreeze_2_r03f_rx_mac_srfz_n     ),
    .i_hio_sfreeze_3_c2f_tx_deskew_srfz_n  (i_hio_sfreeze_3_c2f_tx_deskew_srfz_n  ),
    .i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n     (i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n     ),
    .o_hio_rstepcs_rx_pcs_fully_aligned     (o_hio_rstepcs_rx_pcs_fully_aligned     ),
    .i_hio_rstfec_fec_rx_rst_n              (i_hio_rstfec_fec_rx_rst_n              ),
    .i_hio_rstfec_fec_tx_rst_n              (i_hio_rstfec_fec_tx_rst_n              ),
    .i_hio_rstfec_fec_csr_ret               (i_hio_rstfec_fec_csr_ret               ),
    .o_hio_rstfec_fec_rx_rdy_n              (o_hio_rstfec_fec_rx_rdy_n              ),
    .i_hio_rstfec_rx_fec_sfrz_n             (i_hio_rstfec_rx_fec_sfrz_n             ),
    .i_hio_rstfec_tx_fec_sfrz_n             (i_hio_rstfec_tx_fec_sfrz_n             ),
    .i_hio_rstxcvrif_xcvrif_rx_rst_n        (i_hio_rstxcvrif_xcvrif_rx_rst_n        ),
    .i_hio_rstxcvrif_xcvrif_tx_rst_n        (i_hio_rstxcvrif_xcvrif_tx_rst_n        ),
    .i_hio_rstxcvrif_xcvrif_signal_ok       (i_hio_rstxcvrif_xcvrif_signal_ok       ),
    .i_hio_rstxcvrif_rx_xcvrif_sfrz_n       (i_hio_rstxcvrif_rx_xcvrif_sfrz_n       ),
    .i_hio_rstxcvrif_tx_xcvrif_sfrz_n       (i_hio_rstxcvrif_tx_xcvrif_sfrz_n       ),
    .i_hio_rst_pld_clrhip                   (i_hio_rst_pld_clrhip                   ),
    .i_hio_rst_pld_clrpcs                   (i_hio_rst_pld_clrpcs                   ),
    .i_hio_rst_pld_perstn                   (i_hio_rst_pld_perstn                   ),
    .i_hio_rst_pld_ready                    (i_hio_rst_pld_ready                    ),
    .i_hio_rst_pld_adapter_rx_pld_rst_n     (i_hio_rst_pld_adapter_rx_pld_rst_n     ),
    .i_hio_rst_pld_adapter_tx_pld_rst_n     (i_hio_rst_pld_adapter_tx_pld_rst_n     ),
    .i_hio_rst_ux_rx_pma_rst_n              (i_hio_rst_ux_rx_pma_rst_n              ),
    .i_hio_rst_ux_rx_sfrz                   (i_hio_rst_ux_rx_sfrz                   ),
    .i_hio_rst_ux_tx_pma_rst_n              (i_hio_rst_ux_tx_pma_rst_n              ),
    .o_hio_rst_flux0_cpi_cmn_busy           (o_hio_rst_flux0_cpi_cmn_busy           ),
    .o_hio_rst_oflux_rx_srds_rdy            (o_hio_rst_oflux_rx_srds_rdy            ),
    .o_hio_rst_ux_all_synthlockstatus       (o_hio_rst_ux_all_synthlockstatus       ),
    .o_hio_rst_ux_octl_pcs_rxstatus         (o_hio_rst_ux_octl_pcs_rxstatus         ),
    .o_hio_rst_ux_octl_pcs_txstatus         (o_hio_rst_ux_octl_pcs_txstatus         ),
    .o_hio_rst_ux_rxcdrlock2data            (o_hio_rst_ux_rxcdrlock2data            ),
    .o_hio_rst_ux_rxcdrlockstatus           (o_hio_rst_ux_rxcdrlockstatus           ),
/*    .o_ss_ptp_rst_n                         (o_ss_ptp_rst_n                         ),    */
    .o_ss_ehip_rx_rst_n                     (o_ss_ehip_rx_rst_n                     ),
    .o_ss_ehip_tx_rst_n                     (o_ss_ehip_tx_rst_n                     ),
    .o_ss_ehip_signal_ok                    (o_ss_ehip_signal_ok                    ),
    .o_ss_sfreeze_2_r03f_rx_mac_srfz_n      (o_ss_sfreeze_2_r03f_rx_mac_srfz_n      ),
    .o_ss_sfreeze_3_c2f_tx_deskew_srfz_n   (o_ss_sfreeze_3_c2f_tx_deskew_srfz_n   ),
    .i_ss_rstepcs_rx_pcs_fully_aligned      (i_ss_rstepcs_rx_pcs_fully_aligned      ),
    .o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n      (o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n      ),
    .o_ss_rstfec_fec_rx_rst_n               (o_ss_rstfec_fec_rx_rst_n               ),
    .o_ss_rstfec_fec_tx_rst_n               (o_ss_rstfec_fec_tx_rst_n               ),
    .o_ss_rstfec_fec_csr_ret                (o_ss_rstfec_fec_csr_ret                ),
    .i_ss_rstfec_fec_rx_rdy_n               (i_ss_rstfec_fec_rx_rdy_n               ),
    .o_ss_rstfec_rx_fec_sfrz_n              (o_ss_rstfec_rx_fec_sfrz_n              ),
    .o_ss_rstfec_tx_fec_sfrz_n              (o_ss_rstfec_tx_fec_sfrz_n              ),
    .o_ss_rstxcvrif_xcvrif_rx_rst_n         (o_ss_rstxcvrif_xcvrif_rx_rst_n         ),
    .o_ss_rstxcvrif_xcvrif_tx_rst_n         (o_ss_rstxcvrif_xcvrif_tx_rst_n         ),
    .o_ss_rstxcvrif_xcvrif_signal_ok        (o_ss_rstxcvrif_xcvrif_signal_ok        ),
    .o_ss_rstxcvrif_rx_xcvrif_sfrz_n        (o_ss_rstxcvrif_rx_xcvrif_sfrz_n        ),
    .o_ss_rstxcvrif_tx_xcvrif_sfrz_n        (o_ss_rstxcvrif_tx_xcvrif_sfrz_n        ),
//    .o_ss_pcie_rst_pld_clrhip               (o_ss_pcie_rst_pld_clrhip               ),
//    .o_ss_pcie_rst_pld_clrpcs               (o_ss_pcie_rst_pld_clrpcs               ),
//    .o_ss_pcie_rst_pld_perstn               (o_ss_pcie_rst_pld_perstn               ),
    .o_ss_rst_ux_rx_pma_rst_n               (o_ss_rst_ux_rx_pma_rst_n               ),
    .o_ss_rst_ux_rx_sfrz                    (o_ss_rst_ux_rx_sfrz                    ),
    .o_ss_rst_ux_tx_pma_rst_n               (o_ss_rst_ux_tx_pma_rst_n               ),
    .i_ss_rst_flux0_cpi_cmn_busy            (i_ss_rst_flux0_cpi_cmn_busy            ),
    .i_ss_rst_oflux_rx_srds_rdy             (i_ss_rst_oflux_rx_srds_rdy             ),
    .i_ss_rst_ux_all_synthlockstatus        (i_ss_rst_ux_all_synthlockstatus        ),
    .i_ss_rst_ux_octl_pcs_rxstatus          (i_ss_rst_ux_octl_pcs_rxstatus          ),
    .i_ss_rst_ux_octl_pcs_txstatus          (i_ss_rst_ux_octl_pcs_txstatus          ),
    .i_ss_rst_ux_rxcdrlock2data             (i_ss_rst_ux_rxcdrlock2data             ),
    .i_ss_rst_ux_rxcdrlockstatus            (i_ss_rst_ux_rxcdrlockstatus            ),
    .i_hio_pld_reset_clk_row                (i_hio_pld_reset_clk_row                ),
    .i_ss_eth_fec_rx_async                  (i_ss_eth_fec_rx_async                  ),
    .i_ss_eth_fec_rx_direct                 (i_ss_eth_fec_rx_direct                 ),
    .o_ss_eth_fec_tx_async                  (o_ss_eth_fec_tx_async                  ),
    .o_ss_eth_fec_tx_direct                 (o_ss_eth_fec_tx_direct                 ),
    .i_ss_eth_mac_rx_async                  (i_ss_eth_mac_rx_async                  ),
    .i_ss_eth_mac_rx_direct                 (i_ss_eth_mac_rx_direct                 ),
    .o_ss_eth_mac_tx_async                  (o_ss_eth_mac_tx_async                  ),
    .o_ss_eth_mac_tx_direct                 (o_ss_eth_mac_tx_direct                 ),
    .i_ss_eth_pcs_rx_async                  (i_ss_eth_pcs_rx_async                  ),
    .i_ss_eth_pcs_rx_direct                 (i_ss_eth_pcs_rx_direct                 ),
    .o_ss_eth_pcs_tx_async                  (o_ss_eth_pcs_tx_async                  ),
    .o_ss_eth_pcs_tx_direct                 (o_ss_eth_pcs_tx_direct                 ),
    .i_ss_eth_xcvrif_rx_async               (i_ss_eth_xcvrif_rx_async               ),
    .i_ss_eth_xcvrif_rx_direct              (i_ss_eth_xcvrif_rx_direct              ),
    .o_ss_eth_xcvrif_tx_async               (o_ss_eth_xcvrif_tx_async               ),
    .o_ss_eth_xcvrif_tx_direct              (o_ss_eth_xcvrif_tx_direct              ),
    .i_ss_pcie_ctrl_rx_async                (i_ss_pcie_ctrl_rx_async                ),
    .i_ss_pcie_ctrl_rx_direct               (i_ss_pcie_ctrl_rx_direct               ),
//    .o_ss_pcie_ctrl_tx_async                (o_ss_pcie_ctrl_tx_async                ),
//    .o_ss_pcie_ctrl_tx_direct               (o_ss_pcie_ctrl_tx_direct               ),
    .o_ss_uxquad_async                      (o_ss_uxquad_async                      ),
    .o_ss_uxquad_async_pcie_mux             (o_ss_uxquad_async_pcie_mux             ),
    .i_ss_uxquad_async                      (i_ss_uxquad_async                      ),
    .i_hio_uxquad_async                     (i_hio_uxquad_async                     ),
    .i_hio_uxquad_async_pcie_mux            (i_hio_uxquad_async_pcie_mux            ),
    .o_hio_uxquad_async                     (o_hio_uxquad_async                     ),
    .i_hio_txdata_async                     (i_hio_txdata_async                     ),
    .i_hio_txdata_direct                    (i_hio_txdata_direct                    ),
    .o_hio_rxdata_async                     (o_hio_rxdata_async                     ),
    .o_hio_rxdata_direct                    (o_hio_rxdata_direct                    ),
    .o_hio_lavmm_rdata                      (o_hio_lavmm_rdata                      ),
    .o_hio_lavmm_rdata_valid                (o_hio_lavmm_rdata_valid                ),
    .o_hio_lavmm_waitreq                    (o_hio_lavmm_waitreq                    ),
    .i_hio_lavmm_addr                       (i_hio_lavmm_addr                       ),
    .i_hio_lavmm_be                         (i_hio_lavmm_be                         ),
    .i_hio_lavmm_clk                        (i_hio_lavmm_clk                        ),
    .i_hio_lavmm_read                       (i_hio_lavmm_read                       ),
    .i_hio_lavmm_rstn                       (i_hio_lavmm_rstn                       ),
    .i_hio_lavmm_wdata                      (i_hio_lavmm_wdata                      ),
    .i_hio_lavmm_write                      (i_hio_lavmm_write                      ),
    .i_ss_lavmm_pcie_rdata                  (i_ss_lavmm_pcie_rdata                  ),
    .i_ss_lavmm_pcie_rdata_valid            (i_ss_lavmm_pcie_rdata_valid            ),
    .i_ss_lavmm_pcie_waitreq                (i_ss_lavmm_pcie_waitreq                ),
    .o_ss_lavmm_pcie_addr                   (o_ss_lavmm_pcie_addr                   ),
    .o_ss_lavmm_pcie_be                     (o_ss_lavmm_pcie_be                     ),
    .o_ss_lavmm_pcie_clk                    (o_ss_lavmm_pcie_clk                    ),
    .o_ss_lavmm_pcie_read                   (o_ss_lavmm_pcie_read                   ),
    .o_ss_lavmm_pcie_rstn                   (o_ss_lavmm_pcie_rstn                   ),
    .o_ss_lavmm_pcie_wdata                  (o_ss_lavmm_pcie_wdata                  ),
    .o_ss_lavmm_pcie_write                  (o_ss_lavmm_pcie_write                  ),
    .k_user_rx_clk1_c0c1c2_sel              (k_user_rx_clk1_c0c1c2_sel              ),
    .k_user_rx_clk2_c0c1c2_sel              (k_user_rx_clk2_c0c1c2_sel              ),
    .k_user_tx_clk1_c0c1c2_sel              (k_user_tx_clk1_c0c1c2_sel              ),
    .k_user_tx_clk2_c0c1c2_sel              (k_user_tx_clk2_c0c1c2_sel              ),
    .i_ss_user_rx_clk1_clk                  (i_ss_user_rx_clk1_clk                  ),
    .i_ss_user_rx_clk2_clk                  (i_ss_user_rx_clk2_clk                  ),
    .i_ss_user_tx_clk1_clk                  (i_ss_user_tx_clk1_clk                  ),
    .i_ss_user_tx_clk2_clk                  (i_ss_user_tx_clk2_clk                  ),
    .o_hio_user_rx_clk1_clk                 (o_hio_user_rx_clk1_clk                 ),
    .o_hio_user_rx_clk2_clk                 (o_hio_user_rx_clk2_clk                 ),
    .o_hio_user_tx_clk1_clk                 (o_hio_user_tx_clk1_clk                 ),
    .o_hio_user_tx_clk2_clk                 (o_hio_user_tx_clk2_clk                 ),
    .i_ux_chnl_refclk_mux                   (i_ux_chnl_refclk_mux                   ),
    .o_hio_ux_chnl_refclk_mux               (o_hio_ux_chnl_refclk_mux               ),
/*     .i_ss_tx_fifo_clk                       (i_ss_tx_fifo_clk                       ),
    .i_ss_rx_fifo_clk                       (i_ss_rx_fifo_clk                       ), */
    .i_hio_pld_rx_clk_in_row_clk            (i_hio_pld_rx_clk_in_row_clk            ),
    .i_hio_pld_tx_clk_in_row_clk            (i_hio_pld_tx_clk_in_row_clk            ),
    .i_hio_det_lat_rx_dl_clk                (i_hio_det_lat_rx_dl_clk                ),
    .i_hio_det_lat_rx_mux_select            (i_hio_det_lat_rx_mux_select            ),
    .i_hio_det_lat_rx_sclk_flop             (i_hio_det_lat_rx_sclk_flop             ),
    .i_hio_det_lat_rx_sclk_gen_clk          (i_hio_det_lat_rx_sclk_gen_clk          ),
    .i_hio_det_lat_rx_trig_flop             (i_hio_det_lat_rx_trig_flop             ),
    .i_hio_det_lat_sampling_clk             (i_hio_det_lat_sampling_clk             ),
    .i_hio_det_lat_tx_dl_clk                (i_hio_det_lat_tx_dl_clk                ),
    .i_hio_det_lat_tx_mux_select            (i_hio_det_lat_tx_mux_select            ),
    .i_hio_det_lat_tx_sclk_flop             (i_hio_det_lat_tx_sclk_flop             ),
    .i_hio_det_lat_tx_sclk_gen_clk          (i_hio_det_lat_tx_sclk_gen_clk          ),
    .i_hio_det_lat_tx_trig_flop             (i_hio_det_lat_tx_trig_flop             ),
    .o_hio_det_lat_rx_async_dl_sync         (o_hio_det_lat_rx_async_dl_sync         ),
    .o_hio_det_lat_rx_async_pulse           (o_hio_det_lat_rx_async_pulse           ),
    .o_hio_det_lat_rx_async_sample_sync     (o_hio_det_lat_rx_async_sample_sync     ),
    .o_hio_det_lat_rx_sclk_sample_sync      (o_hio_det_lat_rx_sclk_sample_sync      ),
    .o_hio_det_lat_rx_trig_sample_sync      (o_hio_det_lat_rx_trig_sample_sync      ),
    .o_hio_det_lat_tx_async_dl_sync         (o_hio_det_lat_tx_async_dl_sync         ),
    .o_hio_det_lat_tx_async_pulse           (o_hio_det_lat_tx_async_pulse           ),
    .o_hio_det_lat_tx_async_sample_sync     (o_hio_det_lat_tx_async_sample_sync     ),
    .o_hio_det_lat_tx_sclk_sample_sync      (o_hio_det_lat_tx_sclk_sample_sync      ),
    .o_hio_det_lat_tx_trig_sample_sync      (o_hio_det_lat_tx_trig_sample_sync      ),
    .o_hio_xcvrif_rx_latency_pulse          (o_hio_xcvrif_rx_latency_pulse          ),
    .o_hio_xcvrif_tx_latency_pulse          (o_hio_xcvrif_tx_latency_pulse          ),
    .o_ss_det_lat_rx_sclk_clk               (o_ss_det_lat_rx_sclk_clk               ),
    .o_ss_det_lat_rx_sclk_sync              (o_ss_det_lat_rx_sclk_sync              ),
    .o_ss_det_lat_tx_sclk_clk               (o_ss_det_lat_tx_sclk_clk               ),
    .o_ss_det_lat_tx_sclk_sync              (o_ss_det_lat_tx_sclk_sync              ),
    .i_ss_det_lat_rx_async_pulse            (i_ss_det_lat_rx_async_pulse            ),
    .i_ss_det_lat_tx_async_pulse            (i_ss_det_lat_tx_async_pulse            ),
    .i_ss_xcvrif_rx_latency_pulse           (i_ss_xcvrif_rx_latency_pulse           ),
    .i_ss_xcvrif_tx_latency_pulse           (i_ss_xcvrif_tx_latency_pulse           ),
    .i_ux_tx_ch_ptr_smpl                    (i_ux_tx_ch_ptr_smpl                    ),
    .o_hio_ux_tx_ch_ptr_smpl                (o_hio_ux_tx_ch_ptr_smpl                ),
    .i_deskew_rx_ch_clk                     (i_deskew_rx_ch_clk                     ),
    .i_deskew_tx_ch_clk                     (i_deskew_tx_ch_clk                     ),
    .o_marker_found                         (o_marker_found                         ),
    .i_marker_found_up                      (i_marker_found_up                      ),
    .i_marker_found_dn                      (i_marker_found_dn                      ),
/*     .o_deskew_rx_source_sel                 (o_deskew_rx_source_sel                 ),
    .i_ch_muxed_rx_data                     (i_ch_muxed_rx_data                     ), */
    .o_ch_pld_tx_deskewed_data              (o_ch_pld_tx_deskewed_data              ),
    .o_ch_ptp_tx_deskewed_data              (o_ch_ptp_tx_deskewed_data              ),
    .i_ch_ptp_rx_data                       (i_ch_ptp_rx_data                       ),
    .i_ch_tx_mac_ready                      (i_ch_tx_mac_ready                      ),
    .i_ch_rx_mac_inframe                    (i_ch_rx_mac_inframe                    ),
    .o_ch_tx_mac_valid                      (o_ch_tx_mac_valid                      ),
    .i_ptp_rx_dsk_marker                    (i_ptp_rx_dsk_marker                    ),
    .i_ptp_mas_wm                           (i_ptp_mas_wm                           ),
    .i_tx_pcs_data                          (i_tx_pcs_data                          ),
    .i_tx_mac_data                          (i_tx_mac_data                          ),
    .o_lavmm_xcvrif_addr                    (o_lavmm_xcvrif_addr                    ),
    .o_lavmm_xcvrif_be                      (o_lavmm_xcvrif_be                      ),
    .o_lavmm_xcvrif_clk                     (o_lavmm_xcvrif_clk                     ),
    .o_lavmm_xcvrif_read                    (o_lavmm_xcvrif_read                    ),
    .o_lavmm_xcvrif_rstn                    (o_lavmm_xcvrif_rstn                    ),
    .o_lavmm_xcvrif_wdata                   (o_lavmm_xcvrif_wdata                   ),
    .o_lavmm_xcvrif_write                   (o_lavmm_xcvrif_write                   ),
    .i_lavmm_xcvrif_rdata                   (i_lavmm_xcvrif_rdata                   ),
    .i_lavmm_xcvrif_rdata_valid             (i_lavmm_xcvrif_rdata_valid             ),
    .i_lavmm_xcvrif_waitreq                 (i_lavmm_xcvrif_waitreq                 ),
    .o_lavmm_emac_addr                      (o_lavmm_emac_addr                      ),
    .o_lavmm_emac_be                        (o_lavmm_emac_be                        ),
    .o_lavmm_emac_clk                       (o_lavmm_emac_clk                       ),
    .o_lavmm_emac_read                      (o_lavmm_emac_read                      ),
    .o_lavmm_emac_rstn                      (o_lavmm_emac_rstn                      ),
    .o_lavmm_emac_wdata                     (o_lavmm_emac_wdata                     ),
    .o_lavmm_emac_write                     (o_lavmm_emac_write                     ),
    .i_lavmm_emac_rdata                     (i_lavmm_emac_rdata                     ),
    .i_lavmm_emac_rdata_valid               (i_lavmm_emac_rdata_valid               ),
    .i_lavmm_emac_waitreq                   (i_lavmm_emac_waitreq                   ),
    .o_lavmm_epcs_addr                      (o_lavmm_epcs_addr                      ),
    .o_lavmm_epcs_be                        (o_lavmm_epcs_be                        ),
    .o_lavmm_epcs_clk                       (o_lavmm_epcs_clk                       ),
    .o_lavmm_epcs_read                      (o_lavmm_epcs_read                      ),
    .o_lavmm_epcs_rstn                      (o_lavmm_epcs_rstn                      ),
    .o_lavmm_epcs_wdata                     (o_lavmm_epcs_wdata                     ),
    .o_lavmm_epcs_write                     (o_lavmm_epcs_write                     ),
    .i_lavmm_epcs_rdata                     (i_lavmm_epcs_rdata                     ),
    .i_lavmm_epcs_rdata_valid               (i_lavmm_epcs_rdata_valid               ),
    .i_lavmm_epcs_waitreq                   (i_lavmm_epcs_waitreq                   ),
    .o_lavmm_fec_addr                       (o_lavmm_fec_addr                       ),
    .o_lavmm_fec_be                         (o_lavmm_fec_be                         ),
    .o_lavmm_fec_clk                        (o_lavmm_fec_clk                        ),
    .o_lavmm_fec_read                       (o_lavmm_fec_read                       ),
    .o_lavmm_fec_rstn                       (o_lavmm_fec_rstn                       ),
    .o_lavmm_fec_wdata                      (o_lavmm_fec_wdata                      ),
    .o_lavmm_fec_write                      (o_lavmm_fec_write                      ),
    .i_lavmm_fec_rdata                      (i_lavmm_fec_rdata                      ),
    .i_lavmm_fec_rdata_valid                (i_lavmm_fec_rdata_valid                ),
    .i_lavmm_fec_waitreq                    (i_lavmm_fec_waitreq                    ),
/*    .o_lavmm_ptp_addr                       (o_lavmm_ptp_addr                       ),
    .o_lavmm_ptp_be                         (o_lavmm_ptp_be                         ),
    .o_lavmm_ptp_clk                        (o_lavmm_ptp_clk                        ),
    .o_lavmm_ptp_read                       (o_lavmm_ptp_read                       ),
    .o_lavmm_ptp_rstn                       (o_lavmm_ptp_rstn                       ),
    .o_lavmm_ptp_wdata                      (o_lavmm_ptp_wdata                      ),
    .o_lavmm_ptp_write                      (o_lavmm_ptp_write                      ),
    .i_lavmm_ptp_rdata                      (i_lavmm_ptp_rdata                      ),
    .i_lavmm_ptp_rdata_valid                (i_lavmm_ptp_rdata_valid                ),
    .i_lavmm_ptp_waitreq                    (i_lavmm_ptp_waitreq                    ), */
    .o_lavmm_ux_addr                        (o_lavmm_ux_addr                        ),
    .o_lavmm_ux_be                          (o_lavmm_ux_be                          ),
    .o_lavmm_ux_clk                         (o_lavmm_ux_clk                         ),
    .o_lavmm_ux_read                        (o_lavmm_ux_read                        ),
    .o_lavmm_ux_rstn                        (o_lavmm_ux_rstn                        ),
    .o_lavmm_ux_wdata                       (o_lavmm_ux_wdata                       ),
    .o_lavmm_ux_write                       (o_lavmm_ux_write                       ),
    .i_lavmm_ux_rdata                       (i_lavmm_ux_rdata                       ),
    .i_lavmm_ux_rdata_valid                 (i_lavmm_ux_rdata_valid                 ),
    .i_lavmm_ux_waitreq                     (i_lavmm_ux_waitreq                     ),
    .i_ptp_tx_data                                      (i_ptp_tx_data                                      ),          
    .o_ch_ptp_rx_data                                   (o_ch_ptp_rx_data                                   ),
    .sm_pld_tx_demux_0_o_pcie                           (sm_pld_tx_demux_0_o_pcie                           ),
    /* .sm_hssi_pld_chnl_user_mux_0_i_c0                   (sm_hssi_pld_chnl_user_mux_0_i_c0                   ),
    .sm_hssi_pld_chnl_user_mux_2_i_c0                   (sm_hssi_pld_chnl_user_mux_2_i_c0                   ),
    .sm_hssi_pld_chnl_user_mux_3_i_c0                   (sm_hssi_pld_chnl_user_mux_3_i_c0                   ),
    .sm_hssi_pld_chnl_user_mux_1_i_c0                   (sm_hssi_pld_chnl_user_mux_1_i_c0                   ),
    .sm_hssi_pld_chnl_user_mux_0_i_c1                   (sm_hssi_pld_chnl_user_mux_0_i_c1                   ),
    .sm_hssi_pld_chnl_user_mux_2_i_c1                   (sm_hssi_pld_chnl_user_mux_2_i_c1                   ),
    .sm_hssi_pld_chnl_user_mux_3_i_c1                   (sm_hssi_pld_chnl_user_mux_3_i_c1                   ),
    .sm_hssi_pld_chnl_user_mux_1_i_c1                   (sm_hssi_pld_chnl_user_mux_1_i_c1                   ),
    .sm_hssi_pld_chnl_user_mux_0_i_c2                   (sm_hssi_pld_chnl_user_mux_0_i_c2                   ),
    .sm_hssi_pld_chnl_user_mux_2_i_c2                   (sm_hssi_pld_chnl_user_mux_2_i_c2                   ),
    .sm_hssi_pld_chnl_user_mux_3_i_c2                   (sm_hssi_pld_chnl_user_mux_3_i_c2                   ),
    .sm_hssi_pld_chnl_user_mux_1_i_c2                   (sm_hssi_pld_chnl_user_mux_1_i_c2                   ), */
    .sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp ),
    .sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp ),
    /* .sm_deskew_rx_mux_0_i_ethmac                        (sm_deskew_rx_mux_0_i_ethmac                        ),
    .sm_deskew_rx_mux_0_i_ethpcs                        (sm_deskew_rx_mux_0_i_ethpcs                        ),
    .sm_deskew_rx_mux_0_i_fec                           (sm_deskew_rx_mux_0_i_fec                           ), */
    .sm_pld_rx_mux_0_i_pcie                             (sm_pld_rx_mux_0_i_pcie                             ),
    .sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie       (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie       ),
    .sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie       (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie       ),
    .sm_pld_rx_mux_0_i_pcie_bond                        (sm_pld_rx_mux_0_i_pcie_bond                        ),
    .sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top   (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top   ),
    .sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top   (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top   ),
   /*  .sm_hssi_pld_chnl_user_mux_0_i_ux                   (sm_hssi_pld_chnl_user_mux_0_i_ux                   ),
    .sm_hssi_pld_chnl_user_mux_2_i_ux                   (sm_hssi_pld_chnl_user_mux_2_i_ux                   ),
    .sm_hssi_pld_chnl_user_mux_3_i_ux                   (sm_hssi_pld_chnl_user_mux_3_i_ux                   ),
    .sm_hssi_pld_chnl_user_mux_1_i_ux                   (sm_hssi_pld_chnl_user_mux_1_i_ux                   ),
    .sm_deskew_rx_mux_0_i_xcvrif                        (sm_deskew_rx_mux_0_i_xcvrif                        ) */
    .i_ch_muxed_rx_data                                  (i_ch_muxed_rx_data    ),
    .o_deskew_rx_source_sel                              (o_deskew_rx_source_sel)
);

endmodule

