//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HrWoS4XOHP9aIEJCIJUGnHSK8E2rNsoKME3JnXmVifAUYj/USPMEpSN10JOG
Gugkj3omWU35NlijDsnbeW1pXxWMpOyMDwO9YaeoA/4F9q8rdr7Joks+A67d
31IY00nNcwEi1JAxBgyzh7N9/IZfvpkFjUWLR7LoWtksQqflDcpry6kPTHEl
KF2z+ENCOaG7omgYbVWKBhwiyKlQmUluqMUkz8zugBin50P90Xxi6ItOYYTB
LnYbKYgAB7jVUbBmkunK9p9Lo27GaoN5qGwjf9LrN2hdTwGamQmcSslO/dy5
Bj8c6uhMt2sfZSpcmTNqq2xgXS5BxJN3Yvdq+FOwDA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lB7x/G/t7SpXV6n5y6kjlKZ9ltXlF7uizCda0snJrIadqmveYKGKwc3m5+mQ
PdV5Izo+KI9mHbTUj2d+Cr5sNbSRgZCdz1Mh1rt1Syc0tSPelaphFGB6Lndw
Mz9N8TgvWviTbpocTsNLpJ/8DN1vts2KLRrBFO+JR8XQQLWcFgAg+yZcTPzx
Ld8+TsJbXhcY2xQuD66tKR1s+qtyN5OWFH/lVpUO5cf2imDhzilTPFBJ0FFu
Czbh9jNT7Uz5Up3FdoetMfoMoFp/+i+7ewZP6fOvkqrkTMLI/EutxrvAMWIL
PhglIMpLbJfCzuTDOJ69wK/JLDUeNovWyKeQwt1S4Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kFkewgwFhOBgM3QkYJmmoJcYXVJu/qDY4BHkjm933J3H6IHZ+CDgL8OOnKtF
OHbbtpx3FAKSfALOlzt39au34RmYL8Rs2JZthnPNQm+Z61kqW4gqPtl/gVKu
VW436QLA925u599eUV0/DhFC23RCicHyPkEumrKYrlBIcU67OSen1a+Uyl11
N7jS+LpiTGrqHBTmdecwMIlS+itG8JKZoIWdxpQIXQRSJZ+qZ06p0Rt6jtUy
2OJxeeNLY3Ac3mxGvJ0eDdc2tes2aENKEHACCQ3zd1lO/5qX+etlWjJ/PInb
qh/HQRzshydS3gbc0GWYwiBwCDGC9OJjd7q18NE4Ng==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m2QOVfoqey+Pe7wBZXiaD3EcrIZclg5Is2l7D0icz5T3mxOhP0PN5uoybqIH
ANmjjfJ2sjPoKEz5TGfNutFPaj6I+MYseNY5FYlqbK1SdBLZ9zJd9rlXaY3r
y5PSRucKK+AN3kIEZppSRRAtXZNE8LUOlPqKKgDCicLz5iRac0w=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Q7Rys4di3/WkPm8iSvEdzRNj91BcU4A0mNseemZrK1YhIYNfE8Z8YZGIY942
EyZOzKon5IX5pddfGJBo45ixF2MV83DHg9eXUOfNRytR/wA/M+61IC2zW8Oi
O6Mx5Lsvk2gQIDbqzV1/RhuTUn2IKwDioAtNdcZo+Jif30hCP8lok6CvvRhb
yRRfIjsQm96BTDcERJXsbfODvEu7FbeWmehsaHpDPAyOCyvvQscTT0SvlOQd
zdlLW1hmrjkoX0vQSxBuRsp9JrJzFY+fuDwDMfEvnpj2VcOFT1tH7JbUWW2P
EyQOu7AauK3DqySpjrzUG+puoykqHpZq1l0qfU0zjRCNipuQ7WvJ3Els5cZS
ekBHRhRHCyEV5M+/NVucPsrTCEMGFcd42w0K4o7iA3EAbvzieTma2wj2omPJ
9cxpcsuMe136kiQhBKhy9EB4XvfpK2aADkQz+55jCFA6tc74yRAPt0tD6Qrr
ffOQBPpUaemMp5XkCFHQlMRs1z4bS0Sm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BudCsp6JOg/BomEQuSL3bZXoxoyQBrSo4l+6/281JVrZUQiJHV1R9OOLx3YG
BKfK/+wPFiO0ftIUmSiB5WSXCu7nrVkq5nTiIN1YxvUR1BOhieG6NPf7022g
7M51J6SSI9Hm9rXdn84XX7nHRI6VH62UR6Os1LgrpHfrlGYUVuU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
r0HNU9WMBa8XXNX647tKqd5paO0+m0O/MupIKtld/OFyOrbt+U+DCaKoqGHZ
ZQ3+Nru8Muf11HZxEd77QObUlLh9ZxcV45ayVazdoRF97cAG6PlXkjEI/AU5
8EAtbFIW7Je5SUMpQZL6L3Br3OagLdMZakmL6H2DSqCNjrCw/BQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4592)
`pragma protect data_block
JuPyYKchnO8/4Hr+Vv2r2Z9QjkDpIvDm8nCqXBO4AAEalpddOAobjnzGBj9U
Q8jY75J0v/c8jcqGgHWihKqTnEXvzRA8jY3E+AzkY9HYO67qx2f5PB5YsFXV
75yyP7VRxGEjutlUezKaLDlgDuLqSdBgMxRCcLB0RVobkJoW+lZ/7QX8W3G0
NhVpIQ/Hae25bFeovyFnc073LGkTEZ2XqcTQxpt7NgBeBOwGNjkpWZYpFjXh
TkuIlDEoGdqTY3pxdIh7tM23Zu8HStukfeyw5Y5+ER1LriARwD7XciGS4Quo
iQoXzZeVuAJJbxtDHG0+udWyWsYnyObugvQ9Y3QLlzZIi+qgkblHesWWL3j/
2hF2J1hWOmT9lAJRkGSfgwSTPgL7/cSVotc/OTnEwx5ev+jfV/ykRFuGmJxV
Mq0RKi/mgcMG+Ic4LTlcOWbQtds0tvk7TC6OHrT1w/MK4GBFSZgKZIcUR+FV
GtAV+E46bLB2ubDCfDQBFJyR9kaE+rW+xoxU9d/LOAU5HXERILWpLcRDHBT0
LCqvMW/gxvWoDM5rz0U2wJi5t0SwpZCS2cXG9NvjoKglyh15Kj7jWKB6z/pR
NeQBGDZ9FiHV6CscC8tYVpDiweuWgeo0cSQPl2yuRGO6oGfThoelxxqeGspu
Z1Zh7ne5iDFEhJ4lYlRugwN7+yxsnkTgY7EjYhXoWJMFLqWI265YdrAmiGGm
W77gfGcG8V+0qHSMH5hZVIUUJy+uDplkDDYdk/FB1acwD2fZhSP0kmsU3WnL
qzOAUWkXUwJlvMVAmQzM7g4ekfTib6k/odVm55G4tb+E4lN+jdYGyq7l/26G
EA0JZ4+23/Sh7SlWCINr9Jg5ZgYDnkg6qW+zGwD87ZIy2rQX0/mvYpolcIse
JJBenJJeBTu7UUsAoSU09IyCWQUcGxpetYc0Em2iIH18KhISgmdlrQGBubhC
l6ZMfP1hzzgiF9jqkID6gXsaNf5OSU/ec1UCsp6zV0UsG+6iQ/AcoYA8ajUA
URE6yb1hMr/PtPSuuINPwxULcmS+YfTcq2SYIylWAfKE3CfFuBKImbn7FXgF
SH1vh9mDsn2fBLbau+Sf46TGjjmrciRuqswvPWYK6oMGwRWWDS5hatD+vYGd
r1DiJgZoizeEGILZtJovx1Sewgt8WvBIyLqmgDZeXeyDoOECYKTSH0sdvNtP
XURfYxAUJnUwgL5RhdHYwVcuO88pgmPxvfx8L+g0sp+1xM6WT2N2IlUYrUUA
Nfzkz7hmu/20xfERFbE5wy3/WWVDmkQxnH3pleWyVXYpZ4YxC/Mhi4L06Km0
st9uKvcyrjTsNeH9qwZXzA7l3IyWmuemxu9+5+0vV9leyUNSRxmiDjLUt8mW
gUEE4BVP63GC8zFTzyMURheB8a8xiqd+3iCGKVJ4synyL90h2kN97CbLhZjH
UJmYskvWDL1kln0xNgm0WEiHakG8b0xSpOR4WNI/aVWaWGJFExj9+S/Bh1pQ
vyieliqnmSBc4ayEEOu2fkixe2OZKdMP0uzE5XeIUf5PUba2V68+NqAv7IeB
wsbRjv4i7l8gNqsH63D3cRT1h7klFhIJ/toP/rl5VRcwO5zAsRflqXxmqlsX
M9r+lLKwDk8S0esWGq/7lkxntIhOeA0ZHPmAyfD8XrkY2ne7NAu2usBeiuLI
yPOfJ0rK+At/obOtEd91gchZXnWBTaTUPFb45mQVGLgSaCn42+frKgwaUJwi
k7yupUPBF1hl4n6xAJNB0kFVfg38atEyw5aOL1W6FCtdGJ5loC7NbvzvWU/g
bSrpu1h4BX9tk7B0g62FxXQz6jNb/faiYTzKcTDZnotlugQKdIWaVHRAKuC8
TMnjf1DhlcMNQiTjaZpSLTtg+qdNxrQs1wd+dzS/9BJEx0AJ8zRjqKI4NqKb
PcZx2y9egPAZ5UFoS8BRqPoqS1wSP5A5I7Yz/kZktdMDEnkhXRf5PIaDhWVn
mr/YeIbxsCOIdQ3Ad22o7bmJJEqPdoIPaqTvJ6+fc9en9VqLAs81FBpFr904
1VwjSUai1J00F49jrqB8Gy5awNq9W4i1A/ckSNw92Ulipq66KhFJYKZSxVJZ
EVfstPO86hpBHYqYnvpHtg5RV+MWf8KZo8cGqBaMQ4ksrou2YLwi0o69FI2j
KBUnHaIs1ZrM/npd3vu5JbNcnmSj4Eprhzom/4KvfobNrxLpNLK6PHQenl8F
ITZxzg83kWNbDtTWJIbBNsbSMpu7VDlKxo9ZHbrtXOXs5YZb+wjZcH508wcK
BpeOTOPcM30aKZgVAUbc49wUuXMQljQPBG76vkd7rY3TLAcQ2EVP+8CLojD/
VQeHIRsjxxnMXWmhHg48dc+d03NhLgXSxhc1nRJllPn6SNQ4T6u1lYVPNrC0
o7nm4lTiMRD+MJiTwmNw/tED1CJ9XZIs2cemrdEAXWh/A6VbcItzfogtAlYx
+/Bwpa16Hjen6qm3POYNRN3S1oA5TGqK5Kk1tFzDqAln9zutnqi/tFmmxdkz
yWp9g2exEoUdPALIkerXVGLh+5NBSqPobq3/sBcdznLP56g1QEpi1G3RVoQR
wI5qb4Z8SlVT8NXCrX2TL6cOnLGsofFxLS0bxU9BII9vWhZdUWQR3QFLnmJd
o0f7/59032ds6yT4UNzhXhgTrWlJJapX+CavYLXBiTtT8ij++YLh1UQy3wHf
PlHFYSMFebwAdr3xLiqNAANeOKmN7A11r8lV7W0JNbW6jHt2bF9vvg27n4c6
jpFeN7RLi3wm27Qt+ZFUxixAYCfP5mCnWVzldboGWPk8x4RJ+xBD9TZ14O/A
F0nw+SQ8JNCv1vw23mtIovcBR1FptPH501PZ0adWYaMKHRye3ZbcCV0EsTPa
QZQNA45WXQM7Ay8Xaj206840s0PpZo9tSmRAHHDi+ivwEai/4Pp7R/S3WTiU
y7jD/7YrFDYmaAG03j0ti8GghwhfPCQao+uNMf2M4/bsh9HDv9VTFzaYFRjF
xW4BWisoZALNtqbh1lK+hM7xVcmniTWlO252I2iNkwap8H4qAWLBdGV89mL5
ObELoSrs4Y95Fghne4+JFLEqq4YCyic9LegacMiyAqsZ/3mYRJ4fOxz/6+ZY
v/RC1+0fCzZenlJqV+mwy2E8Kd1tLFGC+lqcmzWJoNK5MiY2NSZlaRV1Vew0
cod5DDsFE7FYK5bhfjcHzSeBtq0KK7SJQITB5QBdMtaA1AKNUS26Hk9sgUkr
lGySzqs6XSWg2lVhERBkAyfWXM+XuDbQmZ/OD0bzZIW4uJeYUZDEKW5B8OlX
3hdx+CM8o+QxFtLHgEjQeADgbA6JIC+SlOQ1hO0uEN14VSo9/n1S1U9lTkAT
x1nVHHlTluQQAQirwQfcjwab+RNRaEIv+lOHzf7fmb8dXUS16ah3fhiaPKCZ
W1pR9euLpUhY/lkd88nJn/Xm4Oe8fPNO7XQhdEdzry4Ag1epslTid+qsuGbM
x5Z4rhOiY5VJsgK7i01KvEdt24tLwnIrRUe/9tMbA3iSUswGod8TvtRLtuW4
Qb8HgPTSJHAIJ+uWrZdZSHjvWpxeDlzgjDsjAmGtTXqv1WXkSp0uM+4Uta/B
iCVl6UfoagzsoejhGvv60pnP4iZ+kM3h7MILzYzbooXazHIsgylnefQz0gap
a7BDAwqkXM17KLMeBpLKAQu1Fm+iE4+UH/s31Qr8y4G+d63/5wNep/dAL+7P
apsDFfxNvMKgPRE5lIJU7orMgcZnCZf78o71op9nL5gkADuRWP3x9IOtrCuP
22DitRe+SI76vueGfN7ZtD0K0hwCwCRA/zM2g1dUYMi5ZT8tvxEmawXloS9j
VCwXsxD35FYXQuodMWUDgUj4auT6myDX22zraldI36MqrGqUzkG+zSZBIwQP
ry+MgqmaAzI1GNxPj8qaoS09qpefEfei15TVezVyGM9EcE0ox6+Q9G/HIqcj
bMkWgpvnfL9m/Ysy7aUAHXMBtgvTWMnJvseiqH6Uhck8dyEUoPCQsKw7zioq
BSEgG+63u3rv+xZwILiW2+LEtlhgkARV9cgfea5LqWqu93uHhBNZD9ye1XEv
awDEgXlHuiVIe2JQhV1lhtbzuMtnv3IWXey/Y5WjBgxONN9jnYl3Azw4Adn0
tFKTqjlvyaqASD7BjV+LNPGUm+yjOuy4/iTP/W0hqo3KyucK/tQ4+NE4LcEt
EhAPWh+fTqhsgTXKJXLbz5ylpP9VgYuUnfJBPjvsrSDfuB5RohGKLreJ+pH5
twkHtHwzjNtqKz+hqqempRaSDrJEghEpH01zIdqdMc05RU8dASt2rCQTSbx3
6xF18c+z3dHSQcZT8o2RTPx7fAbPRmn+oeRaxX2KEygD0jve5Wi4Ph1d5HTd
CFWhLvGf0Lh7ZfiiGxozM9vKXLDdqdJvJRCowBiONRQEzq1fVmHS5ARxegJv
HONT7Q/fOryRUcXvcq4FPD3MLZbWa5y8zPeYJBrNQA9iWzgqq2l1v4HtILlx
vPaTVXwO/8+F5lh8MGezsqRHhylwvxsO2YtdA8HRPKGXRNIeBxlrnTUz7snI
116kOxPXD1Obv7MK5l50rY0a58ruN9Zxbsz8FILuMSfWGz/zl+VVl2yyZJ+D
aJeRcI6pIS1hlqpNkqEJ75IEZsVotXKLpSN9t6Ysc0fDnJg5AH+432GAFRV7
IEx4XRrmyjksVJP0uVefBS1QWgbwncTsBhpEYcWw1lfvbub7rhot9/WHVtvT
1ZnoauDjmc4QLWq6f69QpB5HcxILYJzr+gsk32n5Jhqif8Z0GRHGj9SNVjse
/ZPK2rhKQXw96HAGpzqYttNRHT1kJvMXgrXd5N71nYLOIZFk4c362bEyZebb
PESzMwGr7dxmhg1grWDWQthZKr7bJ6FkLUJuPvA/afitGa62/TPzkefs+vQ/
Z35l8RshRrNNNIoWi9gYr3HNcVrSHpHJT6cAOs0wuAf9DXUDj/i8xPrnhipk
U+BwLd3wsKu4LdvGXSikeKIbEB5q7dB/9ASfx+637aOxHBcDg1cmFff9mtRL
zIPwNV9T2X6fOndlkT5KXB3YvBwSx07t4U2OWDx97BQv6pYEs8+wuhdtMNaD
S2JJHijrs7anXnKPKect9WXi3sj+Iq55Yofgi7MlTMLB5GTSSNMQt65twCak
CLp2pKfTvvY4xrp2SXPhKfqK7XT4YM51XX+U1BAI2l2GDE3qvVUt+vmhpgbe
TfEtZx39i2I7/31kDz+IC/c9V04I7ejHk7jtU1i6UA6Tf7uFzT549CHVpTE7
3TV2KwLAcH2KgV7N511j3C+4snfIwQhKV7qDevOrfksXUla22rVz///dfQ5f
GxQHjNstzrVNclbEs2uqGSIw4jQ45elsWqiqpY97HjSfAd2vEI2jnYCPaN4H
oH6z9QB2bSKzGATMlfTYhoSPmXbOYiKS43wI/J096RaWTtBCVwopxGlv7DC6
JuuRCNFyERK+KGzfdstXAQcWKTRQ+f00a9msOg9bhxnY7YwtCbGEQAAfUvQQ
DPWiWwJR78VPcmmeLpAp8zo1H39Y2l1hZ2QltER+9wi149t5ns8yz64sftQG
tugLxX6W1u1MPTqxyMj5XNz+b259dKGFv7KzFOLI0tswdPy9P2BtkFwbxcIN
7FJXaZOmELHHfv+GVIiZGei3P81zoEaHudDWvUj+EtJtuQ3PV+M7d05vvDtm
NL4qRrkD1pvj7xJ89XHRpz+mtt2Ht+51Y9u4oCGy4y5tVm0gHhLk0SLqPkdT
LXr7/wiup5IInqsREcIBtPGuv8hgr6hB+NwxESv0nRuoSCcFfB8KsqVgD3Ye
W6Qh+ioApmJYIlwwRaSRaMI7HLNdp/vM1jr2IKv817gqfWfQ09rPyc134eNV
T2i42T/fgdk4RJj/KVyW7VWO3JNFZzKc4Xf2jOwrk/U78+eVzTPAY6S5RHj4
XlI2pjI4OJxi5dF6KuXA0SuMKWRqaa0ZJ66smZRnHSXaoOYDIN24IvHZbons
zQsgbplWTs5/PQVVPez4cRk+D/HyHDO1bheFIqBsx1PT2S+0bfdknt4hHMiv
0eTl4JbSvcW0o3xpL9B99/nVs4AEi0+GTYpIJ/A+Vja1vpQRuzAxi6NlpNXG
Ibo=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mLkFRQ37LQsEpWjQ9CnNEw/wJ1iIKzGtFMFSALmEnPAxDCenJ4fPktVHwav+1KtCj+4La90664IMCB58IxoZKCgLShC5ZMdrtGbim0cltFZ4VFQRH6trxSBINH+yky44eEMQhXw72GDES6FCRM6mTQOnWIRsar0JECf8PeYWvc3Y6aeC6QSgALrPKnGMhVM4cfxqkGIDFY0IMldAjWI7FX1ODnUHwfIOircISssSz5EjtOE4p1Abnj0P8KrioV+9xw0ZQNKHLFQjIpGsWHaWR0ytS+inbQZdZ3uIZqY6MM57VT4QtCoG+V9nxsWIB/kzER3QJMm0Sild/RGwsKmFaJGkLtIaoooCvMbW0fQTOYFwf/ISFm98WXU7ttX6MtfODlxglXHWNuEQyMsNE4AXyWEAwvUiFZYE+iOWFFdWWnlNQ/NhBI5nW/36Rr49DhryadDwJDOcayXSTRhn5IQkJ/IHYL0t9RMy30LwRPFY6jtYIO/ARuWHU35W4g90ORe7fNNWBxqyqewvEMPvlW7KmyHXVagibxIu3FjMbp72MQLpUAZThmpfSIJ8u80/mzWC+nfsvWd6l4TkWG6lToL82yKEbQE9fzr+hvDMyu04WLVN945JDJItpVc8xB3pcOaJl4gGgGn/EZoamvLfBmz53aj670apqlWrxFwvSfQDN9GkG2IQuoRhjeG7tQo/zT6jCOjK33q8u8oFO9G6+TWzn68Arcs0xZgywIqwFjhJvv8+akKzFhvO3u68oZqe1XHUkNKEmpMjU4kYXgVJgZX65c"
`endif