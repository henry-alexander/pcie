//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n6OYkRYNPvbOqjdOtucM/Teuz6IKluhfbu/Uny4uHfAJYGOBJ/jg8Hl+VeM7
Qm48QEKIGGWjIdrheRuMb/dAT976E6W+W0Ap9Zqn7raiVDt6ty5mhVtjBDpn
0/NkkF0+dWygIbfRnMYS74ITEYWGgP5IZ80PiHS7GQSOQeh5Uj34gnuq5e5+
2tqErHj/jzSxdHyCgHJf1p9dia+KUVZwGCjWcY3REFhRByuyieq70Njo4ZpH
f8nMSVUUduMFBA0keBEfMzGoyAA/dDCsiW41WmgDBWFAuqjNZUM6359rLjac
A0ppuTurj4LijoZPTFLQ6u3YcGkkXVYNuwvjJ58vDg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NO60d1kdQH2WkjUnwanAUcTvOb0rt2J46mA3Ag7h2/kxkRN3Hn8gcgj1/G7X
4EBnQK7kDgXF87Czwk4PMUvqyxnWaodJzuzdiD5TA4Q4JvE697ifG2d+EaJV
bMIsNAL6I0pSEnQSYdHoIQ9b6A4qtbZUapUGVobohXdWKyYv8hMip88WxxAi
RipbJCmjSMoqSnuvRNWDWurHTo5J8XpXMrpAeSOQ9+lopn3IoDfsw/TWRtBb
dO0g7JxmUoG79Cw+I0pwwMfaJ8vRSb+ZEV29KTCmRuHlb4HPLH0U5Dt3WAOf
XL6GuT0uimSW0CfcwWm+aZTtI1cnCT91IfV0SQi15A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NcyQ/Q0DVl0GxNgbvKckgeaqZGgIhlKRzNpl8ZPwF1hhmOwde8AZlhqwrghg
6mbwvppaj2N36hwlAXIMQLxXQPMEu7V3yH7PHvd5rrpJryAfs74BaRIQLgeT
3Q3JGLv5AAw3nYBdvTUUeFpuuzbrItF9ZvczEgvqtCh9xjV0q8vQvPmaaHfv
tZB2mdJoRuMhRda2ktWHjESAjVomz4B4W64MK8/P5V4ZH0D1eewwmyMhZ0ed
ew+r9TwbpDd0vCU19y2eqfWQTpRzIJzfUfOEr+xiOBXjVMvYHEex3i9cQHKQ
HCDtwn4wmAihbKrNp6KvyhsZWlXRCu7JUmdwzLtEWA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
g7UGnOYBor7hoKdHIQtSijMHUAtAYJh/SpnCWFEe7Ws8v4Yr1CdxLwptWMDP
Y+KBqwY8VeQGjVjFgGIotAktcGzEpJEcm98WxzpYWyiSHxqe1l1IZY7GWoSZ
xyp8rz6UtPfimxT+gEBoomHVlS43JYhV9z5r6g8XAtAEC2dzJus=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KVTmAlcvGFS03cWo5PGA7rPRu6tMv5064h74006p0DtP6C6kLifeghU2etqz
ABY2HM65yiNOPBV5OIiE2G7YgtjcGORNYK+B3bE0whqF684E6VmyH0UtiTXj
yIoSDcS4tnyg5PyB+jbTD2wPVRMV/dmHtxFFJAOo86+ls2/JNAAueyKYFJzl
CYrJ7sM99p4xK08fNyM9LE9XxN78TkJHPzQlKkaDOXSrsSb4LglQWMRqpoJj
EJ0dclONtCkU77PKGlzgh9D9HD6VHSSArm59unh5YVrfJhBIOeFrdYn9i0Ud
spFxH+SP0t8HciaMTX7WZqLbF3YCeRcYO+A8itYEDhuLv6GT3RPVFoYjD9RN
W2k+c0Y+IESU2xbco/9RFV66S4f1CjHpPI16DQNpt34o8fvAQFLbdSq5JevL
W9PfpA8Rq29uApvI2zPPrPDcQv1HSDWbQXVe98KweHyM5rTKxchAtP5cS84S
pVjiwpS2vn9Qjd1JwdfussTOgirAYs8W


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VGZDFoSUNgpJhlOP+l+WQ5lwYajtky1A1VFdSi2LWbBw7/kg7FzhiKr9tFwT
RbU/XQn/FiDhIlBbyQHM56dti2LOugPWa1K3tCMvZm6Z0sxUjQHomG8lJT2C
x1SBd7LLUH9PyqZEdYvnLN+nOIylv9EmyBUmKHmo5QUsd/xcsvg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uBfgvKiTYgEWYVXc4ZvMbe3Z9Z2ik20vgobKC2F4EbumDttjVoLkJCuE4kRp
Q3aEu5AaUWPoYcqVo1nocGtjELxhu3Dod9QrgGGONZlucbG0ZhrxvN1DAbah
HVFDpYAiRtCWrINO+oVxILFO7pWy96SXOh1Maf9a6rvmhsTefd0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 19648)
`pragma protect data_block
74h0uq+lI7ReWJe/hGNH0cBg9SgcqozjlaKohenWeKBdDzmtctt3P0csNNRi
7iJeKX+o0kjZkBjgZWLTK5CnGxZOtK3nxJrCzyWH50Y8xozNc6Z6VaTA2ecu
tBkn9uf/bZKLaCGhzjYxll+wLwXjUwF4UfBw0bRCXzps4MunUAaqGnoOf9a1
E7YyhOAJdzzg4wvUL/xLMZfFPvdUY5LWS65AjtHB6b+0p7IHzEo6V153Mczg
yyW054ZWyjJCSTniuiEB/ihrzCYeaPeqkv/+r3FPmj8dVZxaORR9wGavarEF
ObG6OPYgSzNOMAmmm5yg2Q5OzLoxgpTyNmCFHD/laceVz+Tz5SwrTKUjiOfI
JOzAN3a7Fp3Dy7o3+Ftt3DlE78VbMtHGmpz8pUe4Sr4l6+styDGg+my2McnF
r1gDFwRbBdRb8hAdRjlEFkqh4EiymmN2cl5WpEHeVWGrLJrO0V5wAlNlwvLq
JzO/x17gzYuyLTErOMWTX4kCOtvcVpfNb4qN+lETnaFgZMhPbVlxTGXMZUim
VEip/rvrnD/sREdTtW30vNNe8dDPK5tGCcxkIkZE2kVHafBvMicDO+CygNLz
UkQ/Gu7qJdsBG85hzc06QdAOtKSB32dVPoTd9C/Z9e00JRlPSPvMiVzHEDOq
MJ1zaw2KxTE2ogvMcHEjMapFDrrpsS8YwAUQeyblEtsfQVY+WjKbsw5/u+er
BnStcJ69zvPM3ZOvW+jJkskCtDmsqUnOZdVvJpnagJE7M3dQlPRpmVl/ssmp
jRqmqMZWkwFgD5y7msY5a2/bilcs57YfgMTXkoQ1VgOaLaE+orLRbTvreC9I
vLMsbMtwNVRpbKrjWymWqxDiRobTdrB/fw+yR406Yza0pIfobeyXkITDybBM
z5Q9HxF7Pl9bcX02aWrpBIJ3rx0IJqcarJkPGUy9hFDdlh9dUUxIULu3SDED
tMRCOwPADHAorxdiP3j6H95zHfRfWZgaX5gMnEsdVDYXuiSTF8NiJKkeoQzg
ZAqYaodeYB3+kirnsmnWQElYlrXXSwfKGUoQE6g7iHAw6Son+EKejssi3dD2
gHnGh3VOo+k/H3FJNRUMAZO+oFEZTdZ+qTUuzn9/w7qL8u75Zgi/75b7SPa+
I9ImrXNiEz98eJBHEp2RCeHJlseB8mkWJYyXaMBL9F5+U0kg8E31+c/mCQc/
/ChaBuWIKERfrwCDmzLwrdr0WChxM/uXHwnKGLNeLpPQH/EBsgs/OPpibAEB
XjmRoxuevVj+Ky4v6oZWQoPdadq673bGy56XwQBtImpx0FCUboZr9tdUh7/t
F4bddz0/sLyoYaMFOXcRO5x/Qj1msvQjtHLvnaKhg7phAjN/l4PYWfdKFRko
6P4VncTJorc/c+v7H8wOdbCImbvVWS7d0aN0Oh39hVJZQfc+2ovW16fYysYo
LQHuyRUPWQdNQthudArmXzlt1xk3Tvu8/GPuh7JZ8C55D5j4GtG0WlkCNo4l
G6q885aqHMDGVd7XC5V+QMCuXfMDTzSH1Hl0/+XdWnNudYo2Mc+ZcKDP3ZNx
iooIrgFxKDHkMXSY/RLWvoxaTvoN1ZJZ7hckzW8uaWu6VQtCTYAaTcXuPJLd
oSuvGzyg7KGUh9tFRPJYC/rN2fQ4PAepD/V+3nD3xSEpvSll48o/jeQ+j3pk
DhQFVu+QNgPOKkmvpXxrkLz3nIeWsZbCzH5xqoFBj80XFKUUxIwyW0Y0xqSb
3XnMM8R3vCpVPWwYZLeaVAdpVp8NiMT1ovGB6u2RQFNFurvR82sFaswPK0wY
wBP1YIRMmXu6H2jcwotF2SknTXRihlxJWI4AGqhof5HD/X/Cgb+xi0lKoM1A
0HVpo2uYYDmSkMT2kc3+Hg3WQ5z6MG0dSiUwQfR41wQD6RVOOgyJo81nUa9L
RSk0LUGQlEEe2uo8y2ro+x2dq6cQK0l3T5ePLV3s3jCUeVc7ZbX272tMolN4
0GVwFSmfSFyLm+iyRfnNUUGRPYzBL6U/8oVI1m5G15dieoHf+8Uu+A9nR0v7
MMlpSH8NjB+vSMSlVNe4QtUH1W470osWsb3Mi4ukwXmBbTQ7MZ+WfxO1knou
smqJkIIucH4sc2KgNPSO8kxxJOuQ6ume7UEHa7j+S+t1GtOCu9GXdRgVuhAr
KQbQkNv0P2h7kTDUEdvsajX4K0UtuwfZUiqZpuSvfw06TKkXQtSt998faOnf
kQdo9XCzjdTf0DstPSZ94gyX3q6+pV75dZgBAULjtKCMyA9yMgAPddQQOSxT
Zuqv87YJkd5HDMyinmZ4fS5WBOyCcuFdoEfmQ+hTaJNRCJdDycM+ynG6iXOh
rEmBVDS0BjpUS7W2uzyf+MsRxy4bGWokEAG6so/8vs/yKNMcQEP+iUDfiND2
dZEgeqQXBznV7y7ELYi7RiPElUk4i3OsbHeghoAN3+a9a2tema1+YR4I89pF
pAhLWpGICU7uxmDDwjjRWEBgMIpVRYUsrhpZwnY/5iNnw+gOynb8oHpCmMCP
MMTW0mFdPHibjEXsncz2zOUa751O+LhfnsFwIGct6rufNLrMF9JsplJPN922
AU91Ka4w1Aqds2qU5bXsft62K1IhnIYJi4pgesM/CREhhbVrZ5eSabdupHUN
muAXSjEH7SpG4aXZCuHTlaOiIlb3aGGUW7z7URVFHnS+DqLTdBDx0W89EGUD
1ekEIfklQ+8oO6Yb2jW23tOg1WFui0kzjn7sxGBreqp9yCgtH56K7gpzTR4C
fqIEaQXhWMDz5BXooVL+0x3Nu+cEsWt/jXFUlZIw8sxVXJvQGjWHObKN67K4
TSLhbTZPOwMu6udNRRKYnWg6rYzcl/XgEicxU9+8ft4nEtTE+aUs/2ubmYLt
2zVpeWNkFRO6QXbzGLJlpYoWVj9g4xMvU4L+khMfUrxrTRVf+bqGLnyQ52U1
ctQMv1dRT3QovEbfDp//z9wzGx6a9yV+3Qux9ln+xUD2TI8NljD7sX6ZDQvj
CBTd4xHEHVjomsp/WyUBS0vzooYFfYzeqvyPJ0qATqQ7+LH8k++T71fm9v0P
7Y6pP9kX17+ATwPmba1HUBP2dJXIvAxq1EZGTkUWTTSIX/NBwL/BYeVJiJoe
2HWASL3ExFurjUgRl5m4fDKrNj4F98BS0IpVvT7KSmca8zS76XuWmH1DXHz6
UPrQTU3vo5mRoIFPK8K0a4Fcx0ZMfYKXdIU0qQjaHvT3mv2S3NoGtFnjKpgZ
GzybuMEB9xzZHz5vbbK9qaugGUNT+0MHWz5a/mL+T3YrR1eH1zw4wS1YAVu5
x4VBgoXmG6GrascdKYRx2JGZ0FW53k4fb2KcZdWjpTY0TQy4DZidXCHmARSf
Aozth1XWWfemGV3CpvrvdDrogjsevSmQMLne6HqW1CPQXO/3U5EDftntep+c
QYm/OFKbIQYLr7GpvDflNsy9D+TiuNTMjWF5rVawzFVdXXbdxXiOH3gWf6j2
cfi2NrDlXApGoaLPxqvbtuqK+mOkTHaDCzfPRNHWGAZsDwQ+zum8H87Pr/xQ
5p4YzxUWdjrIrg5r0DH4Rzxl2bY26Sx3AB1bOX2J62V+FuOW6nSYSE5tCl1F
7IdU6ueGtDupvkiYygyb+kkAPuWI4IPxehgvqLvSVeykPAH5Exy8oSoJ9MT8
g20ZnSJLHi29tdA0Njn2YQ4RpF5V+T1AW91W9JU/RbubwiWJV+Hku9sG4Nkh
VyR4Ux8MIVpaPvTmv/UNflY8Zy4XAk1Bh9AxKF/+Ep/whWlqMAlvUgbVQLCm
o0OZdLPIwf0PNG0sKGJRDBMXIsACbCuL42cnprRSFDmW5JVWyikwIF+EQq2g
ocO+5A3W0iLbseDwoLN91dnFpYLN17rYjyWZB8s7hGh1+gmG2Y4T/OAXvAj1
eHdFSXW3b9a70SWT8wl+3LQ0Fv7Bk1N+hj5u1dLWgzaorNR7Ac9xDITKCxPc
9dZPdWcIO3uYrzHtdGwjpTO8QYXJgl9QTkUh7HjUiFRwBo+EkyMd3IHKfY3e
EDJP58BFs33CgdXLm8MkKe3TDWDnZWyQs4Ji7RCK9eDkSsuSuVdKc5fDuh5z
V2iv7juaVTva0+Z3stkpm7VXqVj5Lr4wtdpr75uI/ICEQWEbf5lj52wWPwPY
CAVMy2CscBvJZmXyfpvCjcujQkpeH2urCJPHnVoolLbj2i1yniYaAx/osOF4
DUnyhED5MSq2MR4alXijT6BwsbJ6o/ZT/zy6FFmHFIFFpk+d5xC4AX0mU7cG
R44D/b1VAxgwDywcr1h+FoWFzgy72q7E1iJpWcjkRzhqh3lWT8oyIHpteTKH
6lJO5PoUOF3dt3/JkKHpClX3Kr77qXsVcaYXv8PnDWw8Ko25g5+JIpNg5JlS
0W96+yCNcj9GY9FBM6ru8fbiLUiJJxqhKDUxdY1WPAFzu9MoyapAk6rL9p4+
H0jFFbrCrvNES/uFi9l80wvoW7ttLqOoVU804WxzGn9XTpcTdeThudKh3yFU
c3MnrQq24kfO6SKLbMZb4E/hFCGPz4usmHJt0pyHE6sDpYSiajA0c1QsbQqw
3kXlj+mzHG3ZK5UcGALKM+lVaLUDICdMOlLXA3qCcOqdd/pgks9jD1m1II32
ijaE0OZCXBC/ly8Zr2sRMwBjSxbJBG2FWltlWxjR7zs5vxZxdvSCXac9xUsp
aQXUcrvmfSyfPqXjnoEc7l9f2rOo9XDyHuGu+d2jU4A3WYE0q8fjG5NTk0/y
kafMDce0+k4oy8WeXCZb4XTzexlFffQXyqDi6NdSR71KuIUVMoTulpXL8z5B
x0ufWsPXP2yc66xZcK1Ye18EybcVDxcmpU4fvIfoMeTRnGYhHsOfuPclPNcI
vlczihOTGqexPId3fMntA7Gw2t/Rv5MgXUrT+Y1xc5N4a4633zDbgnXKAzAm
bUajbIUmyfF3Qf3Fy6uqlfUTkoET8RCkXULS+ehTxrqzcTIvbgipvwaE4QwL
a7b00P7RxQ3jWgWM2sQo/rVlhbmRJa/1RvVkSh+Dg4jjD38gxxXBi+l+p4jG
qrvFqWbO67p47SFmv7+1BqfhJOuoymLhv0kMZmNA3v1ujW3KPoTDibuIODD+
wtZ+NfFgnAVZkVouid3+4Brhg6Yi2KPnu7kRdXugRbs2vmXvSM1Eo70AY43z
XwHlhcORzF3ATPbAij6OyA7ESGH5o/p1E8jE3e2WDcL3vycO4HnjIF9nKGkh
5R+CBYd9ZiZmkDxa9H4KrOlxZMs0OGmjNDFFd6tH06rPuLuFMPWgMT1l6SUd
GqXJ41839l3cDbeGSUJPPpxjYQJf/5W9lQCrW8SCrE3rl0rBp9bQzsYFkrZH
z7/KOtwhJXbzzOwJInaYOe/4IWgOfHLTh+3oCjvrDlDK4rTkOlGQM0+mpWy9
1VZTzinp+ZaxtSKZiZlwAf2vqo47ExRBofauo7IEVkLcfItgvdLPVC0fOGBE
zDxgryfRtJkTZLLxS0RrQ31OUSr4BxZTuuG5QsJU+K4uzQt+UdryAqkiygEm
m4NC8SKtX5IlZCTZe5J+Z7PV/gPELmUNRkR5aAs6E/wrorrij12sP2NM4+mb
NUSnbjljKbjchujHhxvvk+qLk53VEr8HquOJRZk+wGblvu8sheLeUvrcnGet
hzUVAtPmprOPdiKYTOeQ+B7cLA7at4Vx5qmZe8J4VeGSJ/1MLORTq+NxpZCa
gf7fEKjekesxMynnMtc0yYnNTsnK1F1KWi/0mtDYTPK0akZ+k/nIl1K6M6DV
flvPtxWj5E9N6Yxix6ephexem9WOpWcQ9V97gTmYzAjIEf4dbRDxEJZRyeA7
4Sh0Uw7baPSsGtga/VWGwQ7EpEWYEJjvdAsGXq6jvS+h91A3B5YQv6pbvAZ0
MJkgFPBaZ8fTft44j6ECM0KlZQlh5xzYSyKkt29h0NSBjOqYS7/BJXroMDBR
s4tuKmPwT00e5/zIgNKX62wC7Q+8qQS6mN4+cpTiv+EPkJRhScGhhNZ71tNA
h+J3QzBay9YNWu4B53I50VxJBKw6okB94GXyhHUoedJxJOV7o7eIGDo1JUr+
WkZ+T+SwO+bLTGm6AIylmvPV/zyw4jYVLYGTd+76s0OoE9VEjpDGcZvrXdjK
MHp/nTBUi6zUMdu8j/NKBMxy6zYSgxi45nIhiazXVQ6BFFDSPIcf7eFyqjY3
hDylnolc8WV/Cj9xGwLuz8wx/TMxE0rPBnhMBgUZWy7C0HdpQAj+ebJxBwbS
jXtNpKisqrHEMEyzgtOsCdX9xo2C2S3qzmjPg5HKBOVVvWpT4JZlqaTeAc3v
8bqFimw+eMiMJqZcPWqq5zk/YBvjpi9kukh5gBCYUk1f6DEX8XL27igHZ3T3
E3oZIWHlvLLV24xGV5JpHBh5A0xq7206lkOdPWDFQ/n4JNTTuMb1jvicQBDh
PPm4t7D6TKEzQe6Z07VPHa0eb56gleNKwUf2PM48fWLe2dJ9C6pZrPlsN8VB
SPlJ1xEr61GjWHzacMhzjBo9iv3k/Lf6+QzoX0P9WEiUCtqnqcqcg/Nf9Fx6
81R9J7xggFznt3O0uAnPvIKYaV4NvUN/0bCwQDZBvEPcIZYweGn9rJobLdjs
2PyAmGnsjq0KP/+zdHA1K1Rv0s50WPIYg0zGSyrHV5aSt9QApPlDy4PFehV+
UOlcARfAjFkomuAfJ0Mk/180LC0PQbE7S+W0zTucMkfCL2ttQsdk2jgBL1/e
Ug/kIAngoYbLyZeXqBOO6bf2ytM/89OmZULShHN0k/Jf+LuQsWmBZguFfteG
Gekn892WKGoIV+bEitMujrAzyA47k0dyPKO87+YapJhXKCWPueIaik+c3nJr
8GJBrLKkj0cYQiO5pZsjcEOpDQKTcjHaCIuKPVAR0nvXNtkp2iVhME4Nik6L
13ZCuJI+3vLdlah/j81Wl4/ImP2qD1WVySxkbwGrQ0353Xp5cEO1ZlzMYkNY
KPi4QQeIU1mGISXHgWsbID60uX2JIM0fMfWK4Cz/EK+e2EWvTj94//1A6SPo
xmQhLGFLq7lSUChhAdsKj4mhvWF4hv13SIpfgw/ceSgv1tfsCzf0v0hXT0J1
QFeshMAiWNKMFITtc6tovo5zU0W3/KG2I0I0tpsliA3NSSIRiCN09S8ETUFI
yCvkcByY50bDBHAzwaY/s/YMq3YncpSEf/jpLncFFmDPGtYWllLckfe/siUt
4UPC23LCwW8dkK1V7jBInOJtIpz6eEYqE7HMBsy9o/RQD8CpP1jayMa7EeUq
95TV8RxYbJ1sluwy44suktUKx1DUhaq9jveGlUiOw3hzACxgjAxh5RNijqYa
01ktnYiQ1SRTKq5WzjcIi8PX8kTGjjW/foGiibCW642zlB64xX6DBFNZ/DhA
GUPAdP0uGW2SPvNqyV1QZYTOxIOS0YMTQ4tyKcdX9/Gtt/JcT6O9BgxNkOwE
cym7BSLfEDNM5kTMXp1Yal7AZTJzskz+0g06lZbPR+VwfhuRsDNm06QqKR6O
iQbkmhLxPtEfg7GQoznrxFyIaeV91pPEdyeZa3ixVrcUIssQ3/Vwxl/E1qPm
TEx072bKYySZjiM/Zq+hDvLNNbnk5O8+gOe2zUOiSqVimTylv/Dq2Q7J+Kqy
hTaPliTD3LrCF+3RTPCAjD51uicpn7+rOZZHKbhprpwdo0HN5SEtO01Rp1yS
KxkPn/Ms8rtKQhXKLI1VuNRQOgvRGxR40laX2S+EvBIzoVnzb3O2Hu3+HDF6
GXbZ3oAzdXvMe2YTcpK5CN0OHeJgEcEn+okmS0/iSdHc4iWoOf+lHTmqEpcX
/ivFcaotNA3F+4ajjGJz58n/2vFTLJWyxUaerRTv/QJUGWvl4jOc5L0ny1fk
mswXc9Cr1zlI50kDpy2/biBFEEp5t/YiSeipfSBIf1/55K9uDlOFxS8RWrrn
VVzWOlNAolhcKnTcvxvWrjatyuh8eU865RA861UWmCnRu5NEaUNgv9OOptMn
eze+rPMrsYYDFTRyDc6zgc5wLNZ8s5x1TV9R6a+X/qypicOW7Fg3DmElfmRB
Q23r/Q/W/Z3Tcn5weeBuPL+leSNOtG7SyuS/LjiPC4E1b0LdNEyVkA6NDZ/I
vomq+VnzVzI5vf7cwytAXdfhqYHq0wzSFyahQRDDpQgUFE8URtzIOThNqrF3
oHA3GgJLiQcSV+kmUiP8zxc0aTrnP2adU8zRJ2Q3YOGmpN+8rL/E2zbFLPSZ
nkfmA7EagWxoSwHoFd+cMSCou0YcxvCOY+J7jLCtS4u78ihkBTHMVeABzhrb
SEsf7h9h/nUe7d89g+uEUH8FWnXssWKAxlwkT20ayL2K8SCnlqgRfziAwuK4
TNsDk1IWGW3BK+eiKI79RsU+8SjqiilrR6go7z1R5HcBlNutxbzukaRyV+JW
DNPRFY93beFOGg+adLHXYs31kPeqbohpyd/mRqXEN5bKD0kgsrVTZIsYPQut
UyVwBemtHfxul7HemDEl86+w+vZFBwPAxfbIUpVfLuTGz6UD9PzJHi9g+u0K
8f710dDL6q+hJMYqDEhTz+Eu5Yj3vBQhxGGobodIWtLbYi3/O+wJo4i8gNKn
ZwVWbcnUs3F5ynVYvLyrY5aegqawe0GE2rePXCV3YXY42BGWyygl1k9dj+0/
iYcIJQd+yvxiIMDEQl7oG3PTOqdxkCg7+MQmBpS2IkTn4ZNPuU0J94gxmp1y
D5ENzIEGZkPfKW68PbEiIj6aVaIce2rKVUnbvZQlrpf203rlH4pWj/eg/4vm
Vp/trMXi8x1Q6w0EVQJBZc6s2bzOfGtCFdoMyo3ALy6TGzXzkX6E2Y973eVM
QUDu5rceAOsXSTLiLHatrZNI7z8Zm1U1HYNygykbSe/PW2rl/UOS/G4qsD/l
Ba4ilMMpkBeKPn+SVY84PmsXPue/Md4RA09PoZ2M1rnipBfmJfYLaxCxEAba
juxH3i8prb183ik7N/9Lo6iBx5rt6i3bPC0sSPWA0gBavmSMHcESev9D3S2m
KWrvIZ/x0fF1kZXXlI4cOJfZ4qmDTDtcDT2/k3RtiXL1nK19lDSsa2E03zm2
wB+ei+mhz8VKHfeS5jTrfDQsFilMhHuvlWdFUgyF/9012QZmqF2/3Cf2kpA4
/MVSd5bp47RbSZKTTRsogzeoHCcuRzUZlhlDDdsEvd4x/vTtjV15LdwH+mAj
RntUSTNLzlGkeDdttTGdvMWvkh/V0JCMKviDx8GmIkcL/bychUuZM8VNOKVp
FS+kJ2d5WLQ8zqjKuGC4tgUtDFaeuDCa2vRBPxE+JHDXL65/mVTMrO911VhS
9FnXkhnk+BdQ2jcc8H075RMpEVWMoUap9gsda4Klyzy9Tv1tLYLxy781Lf0G
FbR5MULfDDn/UHQejZSyrVyADW8xVxjSpL3oKpzD2cBxx3BoIZgyFtLszqn2
iDsxkx8hoUNKdssCVKZRxs/JmNkbH25SmDVqQfX6u1x9xkIdtUYBCN2UbQMf
u+tyxYyIis9dfSuKQdkDJi10KIgWpHO2jaRMn0TzvHWKxxlMAef+l5ZD/ehr
/Eu6utpM5ReaMzsFwBDINDCV0k1BzWuFzUysiCFLqclfi0I4pEVp8tC8LR+R
wC4WPhVWY5uzy5Q03bnveB8F15591gv/BPvgaBUZOr4+cX+kb3yUWrAyQ50+
y1T3gvxM6FPGHR76YsJUM9qJGDHZqOgM16Ot2mKXwdeVjQzoux29T2rh/6ue
OMqUMWnF3XZvBjEK5uxqrh9KWWsHlrR/CwAOcx/F59cXpyjWNc2Ts4DyJSCr
TFP2u4MtxpiT+03+sRXnrTNXgvz7mqK5toc7egeGyiqHTbMZhqcsSpv3v+rK
wfH1imv4HRp7m4m7gkXXPaecK/x7l4ofhw1CUrv3X9tyNyBX30GhB2D+a8EZ
fpx9WWZ61QN1na35BL/YI0abicce2uYYmCIHboyD18BOnyed2ziy9pCer/5Z
iGKWfUhEtTeMXOeKhF3jcFxpovElL72+wMUnbuskjcBahU0Nm4crSw+TAHD3
l33KBnFfROOvX5+r1wf+KBQlfRHam/cnBAU8yXMKIZrOAJ1izAZ7QLWNrltR
JQFWGFecfCsjavLoNGYDdU7YFaA9H0kn7kQUkAgNmOVXtEZS4S2fiU3qJo7D
GVA/N4qxcHCSC5OnAkEg9K53S505Obi3XjzUFDW8ZA3e2gFeU2TCCRGfZwn8
fjA4GshxSmESXOL9uVgNFBIP8YZwS96pKCMyOIranOP//QOFmZVBAkYC5DQH
HLNHyx/8NVmQ4PFrF0qi90MGKKXhPPw6TxfeBQ+REC1Q1z7lyjma6R1KcPjJ
yiI9v+PI64OVb0IWyGSMlSbGvaA4iSH/ErTDvPIB6s0Sy27WOSHvOw8ydIPq
qwrywd4CsfAW/AWa5t/sHF8665lXounB3ucO2LzYUPjjGgGEMNafR/rWIiwW
BELsmc6w0exGDxyAJCz8SG5SA80tZh+wtWvgLPqA1anWg9V9P0HXWVhlcR4d
E9gIDdE2pjSOquT61x78BZvsMQeg2ICRhDGaIqGq+8UDjCSUODr97/4FwDx0
hJ9vtN5a/4DVRiX8oMciouZFd/E8zsbHivUTrEIPyrM2VqHdZ6RGuCY2pXl+
hZU1+LYt+ZtonTfn1Lwf5Q3nh1qLKEKkoPPusbq7HUW6Je7XSP6LxDN9JB1U
vda4Fyi8vN9Z8zbruyv+A0Wm5wMjDk4FG6DoigYQ4pipUIqMiAWVm/589aa4
WQ+tDtPElMznRWbbqSv7WvSz80aNlDa00TXSN1yhIjZEN0VIGSnrMumynt+E
LaLFxWNjRi3Uw/ZMv5WFq7/MXEhKcm3qIwsBAKchvVr0sknf+qEwrW96wM86
DW7rkwrTFZ5zV2KBjeDwCGsjYqYrTR2MimzqccU4wLEEJqZATQegT1UKP0aJ
AyJu8NRZQFeMV0eM2YKUHU3Jl7vkstfNws6SNOoxubB6ryzNuwY0mXzwJE1s
JAqnS3yENx5v1YzUZglzFVbVg4QZYZjFeW+8GMd25/Q4qYrss1PiUXjuZ0Y0
JhqxZcdWAwE0yOCdAbeaQivirfXcbj51DOIVOeiJmKJbH58emD1HiEeUxlHw
JIeT1YKpugMmQFbgxKPDmRAJKwDKSpGemhbtMXUdEgT6TQScPU+KDx+7bSQ/
TZ13mVeSc1aTD9dFRLdrNFBPEMcBL0hgfTwfWrVp4VN3Ff4dge7L4qeWKpg5
v5laUwdKUEGThqMzEYyFOlcJTOSfK3czjgfmczkOxdpALmKwv+bkeE/z2iSu
07ehMvaE3BteZgnUU7+9qGuWuebOrfmMMppLjPxjaSwoZbH8mOQlSBC2tIXU
gBlpf0K2P/vbSUqy3NLR294qOMSwlpzbtHuX7mrtXlMiYAl758qk5olqDaGk
pa0EtjMq0uPlbMR6T1rKwk9EWseoyvkF+ryuivtugTtjnO4pj5Tl6v1KdQkv
zpDkA+lWxYAD3oXayktqieTFFvVfGtZZemg2oVVLTo/997jnxnzPwyf4HVtT
Hh5YLptSAxlzgidH11QE8XU4tN281xVp2yeIjATEc9gmZmXDiW6Wf6bVfgdp
qvQuCSTiC9jQqngSroo5khyErKM9X30fzvU0ys+RixfqMiF5fbHKcG+MGVIa
POh2n3Bh/43OPPg1dXn5OdSVDNMawpq99ScLnIRUEeVjPJBqL8rkynvnNLjn
GUt5wJ8BscEHYe2AmETZHjfueHhhKchDXglhhC+i4pa6Mw6v46v9elftgFLi
GwVxqFw2a4IkuVNaignv2vFdWQ7vLOCpdkx3ckAqFiibnkDHVjzTIgUNSBgH
hDC/MjMuglB5z8w4cbPCl6Vb0wYvfl3zSjCBzxMwMDPoP+nlRipNySt1Bdnm
AKDziCItNUGBFciWUV1RzBPfcKb+K0xouGEiY/xxV8QWvixufrw8Opz0mkki
A4nmokFT5DlWn8KmZychwDgQwSrs2c6a6suYW0zXj/NB5IILfLtd4Dg+d0xv
Oi2L6pqR3cvqQraDg9YBIJ0d5CDCrT67jdOhU6W5K4vz5UF/xzBE5kzLdCLY
C/Z+AIXEkyWifzcwvXumbkvGWivs4107lMt6iRfuh26kvP6vQ0XZv2MfZx4q
OYA0Xnm2zxQ+rS7yLnRo3ET8RfwByXNCIWOOVAoOuWuA9fQ6smfi4kUXmwMU
Y4FPq9Ep++guqMLAG2/U/HlKRSIlWLymxnHVx6CzVTubhTaaHTInKkFsit6q
XjduPIcswlvm/8DobDHJ6lUull+rqGptMfMvLjOoz284SgrNAbFjWwRldPE6
n3C9JRQXELAEBx+VkG/hQcoknnZVmaT94Jw8/jNTiB1B9meu1ePCZTnTx9K4
pAYKUCV0qNRhSDzrdiVV+dudWsYIzv4coAxCpTtr6ArwtUu+4ect0tDuYeOi
RhsJBiUL4XUTnX8o1t7SS0cWjTgLrb20gapkcwxacerTJuefD8upTSw5wOn6
HDFPdHhSoWO4gHPzjfrmMTXvK5ageMSr/RMkm6RgY4rL0RHi6q1VT2HK+8Sa
f7EGCOG8zlC69cbKgpwYVYVKaTEkJ/4yIY8kD5Sl69rNQ5OAIPHHsAzrUpf5
ycM+qbTycsQwCTSbgzIkOTW5nt5yk2FiinF1dgM141NiMF7hkvXy9RR8W5cE
AJ3ZrUEgfGpTYrpeAQBRdouYN2M5tMXkZrZVthxnKC/ft6SjHYPwG+g+MFCC
QhB1HBW9srY2XxKUwUVtFflq9tLbDaeAuSUPK+hiDex5v/6NbhMwkxq5OO3/
Se2HlFt6Z+Dett/ViV1UFaOmQHjGy9bU8OB4LkB0uMzeAa47e8yrBnJZ2SoW
n9kLU2Ggcxa/t96RZ8df1QbS3sXM7DDJ1Katr3skW0j0syVFS/tYj3WUjzB0
4xeTHRN+5WX0ApPx4sG70v/rwrTCKx6KEGZ5RhQ+L2UMnHKf94JYyphfHGcy
ZLXO8ZQOAXDorQnSMsmZXAGJCKzWDnjX67orAXaYHFgM0EwUZgE/mXvIMOdl
pGwhvdQafJAam0mG6T4BBAMqgjoqHfDrYHzhYm07dIDkZtUPMz4pYpCM8e/r
Azm2/qDNW0lpZzg2ZjqKul09l25utkPBo/W3PSgjNR9bCxX1dqLtSLo9bBOP
mQOWcz5TF3XTwD8zOEpkmZ5pSLWjLuES2kPa1fsvhLkNdW246CikvhScVRLI
GVziw7AHm+Bb2TKpouGE722WXw2vV7EDNKq0zEKxr9wT8E12tAmX1uwcmC/0
7suoPGgbn4ZFTdjZWzHifjLlmhD3xmBR+vBhQ6rwX5d+z3huyPhUKoB9iu+/
OTGdJeWspTDZ9u0w3fVkF1AR7/yp977U9RKMA76BWPuuYZNvEfRyJlJ+Braq
ELLQrtIghIbTjsWTznt4oUYmBH/DWVXGKX5i0p8jkTxpOP5DcrvoaPMioNB7
Uz6q8WlkPMvugSNTl8mXzcJ0J86x8/VbUwmgZqYpmP2thssNSJfpQyRtaA6y
LZlWAitA5SON9eW//sqAEVN15z5RLiWvf1yclJKOKkCI1ub1qtEz7fn/CFgR
4vANB+PyVD1U963/irWBRO+hc35+5xXa959Pw23e37cKGFdIcwT/sWbA03po
qwQBSHLGp3GLYV0mGuIoP/QbR2G6IfzmW7yEzsT8TdleqUJgLwOn+qqLn3lU
hCe5S1s2zO1WROozB/0a5RAT1XbniPQEDve0ndObPspri79+xbOXTL3UWGAl
JOAiXuNvg7QCi1BpLboS0UcBmbO5r40K1/+AfHiHi4TMGF/jj0ih93P33k0V
hLUQJv5PZ7w8BsBI9peg7USzbs/53VvvgJ/FikT+qi2MHh6J04B+Cfza5Vif
71f7xC/+kwF1Op8Gt0QiMd92o28NwQNQvl4NUFhql+GwvS9zZQSUJifmaeaH
vWOIs6wCATXWPv239YUfHwv5NxTCUeflqZQePhGYrC/BiwT9aBn4q3CnPpch
Sw/xQRU83Kz2ZrZ/kYu800+jDk9gpGu5/q4M0gJaOi7B09yH2UQQIh0bUXNt
085L2Llyk7bHzP2hFDJYXn21vx3sP/OLC7x/uA2Z9ZXcTUc0itkjZVC19eGo
DUuI2bKTgYWXpiZ4k7IdSG4gLtuMIe47XLGzM3gGOTVKm68FVYd/oa925Kxa
KG6DosRSWSm6buDlbtl1QORMtCCK+Brh6gwJdFMfjMi83eZyw1rmN/v2d+Ch
bPEgSdPy3irB/4KJqvkTbjUzB/F1d4G31wPK3ng2FFblykVNalHTA9+dx8Q0
WbyJBsD9Gtpd3nfNWIseYwGODtQxVlhkHHkHx0tG3D85yD9pnbjDPLG3vru4
PSh4TgP1mORKM39sZ1t66jmcWMACW/RZ36FbYFJIIBm1dPwJ7FZ9hQxwK2JP
ycaMJxaVPHcY/5TwEfnOz10JDa961eLHNaFuAGvqK2SlG+QrMHhtTzD5Xl6A
WhDUe/BaWXWsqUFpAylgtf8qHrh4LqLTD9KgDG7yeBUod9SvuORzgPNQdye5
7fqjRIyRIsKjwZSk59oqDoaXN7H9CJGCsFR/WEclgMPREX0n3i1B3yrNygVb
Qsx5Kb4PBE/UeiyVc4YnIUMfVHugC2M45ujIGWNHUl3mdN3pFxlEOWUX9vXF
gx08IzmgrEfY4/5QDfv46Y81tNTTFAU2KYTYpN+gYuE+VNSmQaXtObIDfetQ
I1jEuMVAfkMNG4F9gcNKgBlBDKRmd3ts67wzTHBMJFQ4M6/oLs46SCsO2sR7
NnDRYxoOvVw+fUsqmKZcqhKv8i5KXwBGm+EYhGC4rJdYe89ED2bxEf820M9Q
A5j/+F0FoUcpbEq1lxki2pep+aA0sAfFChCj0YZoP0NDVckero/6ENRaMkbj
IWk2+t2KhQgTcR70qSSH1m4KZv9uezz4YaN5IK3TZnR2awV+ZseIO9tIikFN
SaCkLDxxg2RebPqiCuP/6TCwadUxKbXLVJo+3xp7MCOiOlmflV3ngUPxQQsE
jendGyS/nlhofmrMl1beTsgmkaCjhoLEAnNQWKseQE3T8vUrLn+gLQuRNVTe
nhwIcpcApF8gxgZOSfMS1gRw3SHJZPHeF3W9G7ifg3kTm481iYcw/r3H4MNk
MoI1vg0dYcQ7e1Hx73KQtpUhuAvIpi0HrFLMCSQWJ2yW9pJSykQfZhcdCHsL
xUWl2RePpl/54YzRvvikjHYleb2cJqq82HCmqrqzj/PMnCgUfCMF97/ayopD
8Nza95eP3s1XzEWdzbWzpvGw9Iy8wZzUW8N+C9JwfTyEyUl9vNHVhYFWL5BY
hyrwl7ClkwI3ZoK7/GSTOsJQTM/AGYvEY1HjnKJFvPxabF964huxv2gupuKm
7VR0d36r+e7g9U8jNuFKw0t8m/WLNhcL0qkUG7kdiDQlQH5TPMz+V7Vsa4Ae
1KKMKVSfWgv8y95mKPF82Sz5ENg+swZ2xlrTKYU3vJbMkzGAIHsG2G0HQSRq
yMPu4UE/HzEvmigxAAT+7H5PQPy9vXyypu2+cdpEioFO+qLAzkYDlL2GTr0V
kWladHUPysWLGVFHY7iO0dDs7r2hcnpklV/sH4PUAOJw3JmR7Tvz4AlrcCKE
xghuX2u3T1mdrN6LKsHh1VGJFzSZ1gw96WfCtsRnHpKoA4LUugSR0RqteWhp
+VQjlUabQE+avANvAzfe3YP3fnydFCKx5/4sYakIeekQMcT0SS3/CPlGoyBE
54E3SrzRJjFYWMrXfm218tVrRWb7JMTa1grlBxNqnI6T7NzxaNHwl1DVqEAP
NMp95ZULiqEGwgqLA6dteU7DyWo+PhYDCaGrnHFtzoiQ4Rt9AgsZZf3JFCjt
X38hMnKgFmP46cuT3E7uYhz9SSV8ZGgS5RjgTCtm9b7RE5NIV9uBRJMYDIyZ
+EpvfmRzlp7I18hw3nJz4kYzmrWgbt/54dXfANtf2EbwZdJo8DQ7NcPDo4AE
Xj7WJrt6lKnIVt6lhyiWoD94tnrnHlAly2N+trf+kNEpUSTtBOY8ps4hB4j2
rzOT5TxlxBiI4mhr2dbY4YNjBeFS/dcH98hcne0qnZId0NFRcoZQ1CUH1jE9
Q/C2+DXSW/fbQ66vj8KAJph3TjGxv9ctuzHGF3l/XdXYbqjlxpXD1SPPd1TW
SXBj4OR/kYiamF7YMupHFQvc+/bDmJdinf2piZo8H6f4eS7HwlSgnUDS7bLW
bUX6oMiNolgiKz8Zpl7F6BI+6ddrcfb6TN8Ql+3RYpCY9VEC3eSbDOu+uMuZ
8lF0OO2obMYNusTtkVSaZ+AolkAbadotRibfVdaulhL6OBxJjSDgaJE+rnP0
217U9wQewaPjd+VIUemQdX46zPyXFKhpJjzUur/EayU23dVJ4WbDptbuKlV8
KDpojtFXcYPFec6w4Oojp+/GkDTTDLzkn7hOzzcVJBLYzdSMHUl6Ki7lOMe7
UD6INviMdTUC0I48xGT6A0cHunFvrv33aVOSlns4LzY8WR/BYlMJP5+IcZfT
ZxF4rA/M9DuSmsR3Pmcn3JfvQTTWyidH5ChNik6N1jTz4srOYzQxuWyxDKN5
1oUb9l1TUMP4oRyBnbszaIi7p9N5FsC6ac0ICrVWHbF5sZZdKDwWi32Bb6fQ
A9GQDmvmRPXqPqQ7NoCSr1uZskidHmcF/UWnbSat41a82j8CwFmflNxYTm77
AQcLRSpGmokoxOC1h+nAv61eelMSpIEsdEc0xk/YmfLiz/x3yC37OGMpFVWK
Lm680q/FpAON8c0+HrIZh/yTzug3RLGLcXtt4yBiDTqKcHi5joRUVAAx+m2Z
rwBkMR4rGkhjxflyc2n9M9OpEDR/z7mvqhdjJY+/nZIOM2hySritR4sHjumv
SxDLWeJWTAcfneThZTJv43PzVKt8keB53orM2Et7kTQ/xGzJzEqRn8fgtj7Q
oOqZD5iK2jmAyl15Ec761f8jh0vwedzoX6BH2chKBooIMkZq6Yab5pUFl8IF
OhLJ9brb87fxzLrWdRhuweXPo51rwPBe9LEw+WB/XvmGRjlYCT00UkQgwItD
ZIAxvkMmWERmAhoDtgZr9sfw2frhU9TVPcWMlhOVmCIUMkzgcGGhUuNvRKcA
FgmiqlQebny4Apr9uJLdYOGRnAMCtKCinIuSCfNLH7C3KlCZFwQbZ6l80OOL
c4vUVNLA8dwGeP7LyukB6DPbp1DuJJx0tUsyRintC4jJGyOzukG/EGpx1B4e
UrWqNUdF04LnohueZb1orWyIl9wrNiB8EozBwv/KiqipZzGTHQvk0wJ2jHsG
btuhSffscRVWbKx1Vs0diylAz1idrCodobZLubXMPhu9ts9qXOWSPoHKQ/3s
DpVUV3YijLBlkhmgE6hzpCE+EBRN1GZqAbF8MCIyr86MseiSJ3GsPd88Lb+W
85r0HfHTwZ1BoswB2/Kv9+u7MWgaBarKoev0G9aQl09E+1q68VM/p4PgfCHH
n2FJ1bceREGcRcHdulMcZBTyxD8b6Dqr7UWKE7AdL9tDQmh/pAmJoLunQnuw
NXkLmJn1rRsWrCwUKFqENtVcddbjQgkObRzIMeQjWVHCp+amf4tQP98iq1+4
VxuzTI2cNG2F3jSirABkj/id8fYGOOSoyuVOixLOpWBxFQlCw1/zg291EJg1
cST53QgU5WTg+cAAXAAFdTxyuYnUr3A8hEU4iAZVLT2z5bqk589x/25PUctn
HkwNaKgROEMR68Jkv2fAZZsjteOcbbNjwka5gHOSImgPKYoZ5/oHezfxu4M9
EalrFDxCfAovvHRNe2HMU+MWu9VU9u/KrA4dHMP2TrlkCRdhLN6BDmQHnyV8
u3leoxFowv7NqX8oZ79lEhHIXFH12FEwooc5UFZyHYw76yIUqurQikdvYCHJ
jCNoNtgiLOWBf8dtYjcFaCza7dKzqcn8hcjYPmEJRE5iDkqke+hIAvUs+cxt
gX943A3R9ysAi0cs2LwQrzMeUEKiYPSHKHWFpGTq/E4ZrY2CdpOVOrOY7APp
uJN1kxzdLA4nPvVSM6I9AMH4/1jE9wPC8u9MTh/CdNIsR1lujBArOPe0QB/E
ETzkbbGhgQ4gLKNjW4z8VFW6xNXdqCK8kIDMUC3S7IZ5qbwhOjZIl3aBoZDl
xM93H2df7R1+4z8KWCfv9S8OejZRH1gbpzXVUVgye+2jL4LHAjN9qIkF3TFi
e0REgEplkhk0VRWSZxk82lvWlKCSmmP+4aKSv+zHZvoU8bGoq1LNo/hPRAih
KBx7Sx4PLCs9SaMvNuRAlY0NXMNtB/D6SgXXN/JPdTEFWlCJVexPkE5TdOob
CjQM219zwNtlpCrLW6Z4LbXvGGiS7bn2Zl0n9hydautPLSdSHI5/EbvUtrUR
SHa+MzA3NaesnRRE+7EfYaWg5TKhTOC8EPIE1sQCvgwnWLyHhuGZG/ziQdv+
3mWwu42fd6tNIixqRG1FXpWT/yobt0w6MZq4boynEo8QxaaHj9biW95eLxZy
5ItBXF+Qd+LM9PTM4RozohcIa3C1dGuky+kF1Dun0bB3lstzoeZe+SyXoBfA
jA03m+VvOtMUXKFi8JCZzGVDlpBg4fbrLpL1rAY7THnUob6hJ7PmBL3aAwvd
QLIJm0MlqcaTBhNw0czPfx4+em4KAl0DG3Hspl3JuVB5xtBgrvoNpnJppo2+
Wkw/5Jhyo1U0qBxo1CNl/0znVkVAPvscPhY0ei8tHyf+LcR8rx0C36gOxfkL
Q8u20VBooNuJuxiG5kAq2iaQ+xqOg8LELANcEhGY/14jpE2qvftq65hsqy4j
GE2jvYJsXOUh/JiPgchjQhtZWCBotYskh5Ub5+eptgopNLWRVrR3BBooAY6p
onNi+XEKGUjqEQn1nqDyIxlrgw3AVFbUifIlzRWWhfnM1QnY0FabNctc4wfx
jer57D2wNnlrU5FcOO0lk2C0LY8R7C5XVcCv8/HgEjIVVOTIZ9RjrVwShBmX
XB1RjSZyxc5L45UdWu/bNQKJDcNQ846xm+lL5BM8tnXohnO13uRSQfXGd6YZ
pqo0vmkxCfsfan2HMNNy/Zoo0ioGKhSEqVWiTQ4d/M6is2aN5CGto/kp6isS
xQPvsE3anIMXy4rMW3wIVMu2Vt8lnEsb0kuk5BvZ7jFa24pxi9coMVBDyITZ
KoAlb/7QdPdOtBJSNLunT7rGIZI5rvinksoiYNJZGXUNjxydQPxK8qds6Wtr
dUfrRZoQWjoUF0XiP0OfaEpyVksF3xTlh86lYxiGZln7Kd+aP96ytIr34k+L
OdpPvVRkO6MQqGWegn2GYT/qiFtMKiEHAx9AsibnYpibQr77UMryecT14DXp
ZF2EvEDDKayLo+zOhWkYSmOcmkrLZXRhiKlUmq2jXvhL0LfuefLjdOeBaZDl
p/Rcll+u0yEjGcz2a0tstaIEl4ZflTjT7akQDdO7exNipg33sysx5h5+ahvO
Bl/il5XCwS5nfSv15/7qvWXM3MNYLrNv0mkZu767QxkASSDB28hBM7iVnSbk
4cURWNkEr93xAjCZPzQkhtd1gB4v0YW0BrmV9+s1T9cQ3NNfYDxas0VHPP8i
G+wK+oC3wXdrS70cJR8ZGgKG54st+Yu0XmDlpxQW2+0jyXz0nMcetni/X6su
uBHNmsrHQYWhblDBssJmkhjAkRBMK2O0gZIQ6ncokjsDpINusxTBsP60ruXX
oYTcfB0R25YF62oJRYvsArrezUYujo77+aTMQw3rk260X/sBDabxuHhNxCZC
LrG+Mg6XpzC1GHU6JgM5ZaDajSvQdIaUKRnvcLI/tnNrM7XOQ0a77Ok9Elra
vMCHGN718Wwf0ZBdB5WduJvuP1XOxdVDrnP6hHrxD7F0RhhmILEvSd55A23G
HCv5AX3mnX5uguIQIyoI7/WBH9MZBl2AB1620fubfI7ISg6bTNN56Dwcy2Al
HYESGaZKtFWPSoJN8hKNqsxchhlP4W+N8aYgdxHkQk3jc7py2JXGxOVd/bhl
sMt0EJES+/hNmCtD00Z0MtxM6EcDb2TvNA3bca0p/fDw5bCsiVDDdXZ7Qpp8
w5B1CbqNbSL8bh1OUWkmE7QfgIm7N4i1FiNQSk0ibUU1kUMTsHLxv+wCZCP+
mOqc/wH49JnjuhZnJhJgTYQrMJt9vy3QZ7VVWC11V23whPUCz3L87SzV/jDY
TqlKxgZPt2T49OVsJvSmNSFJKxHJL24sWUbu2fNkTSnzTSNxnhbi8SbQ7I0u
iXODyY3Tz7iRkRI1+AjBjU7aWlE+UAObk6lR/TCwAVNSzKD3CjFzm7hh3DF6
qIw/cWwgcHpeXOHN4QPeJFPx92cZtqNixEfBmxkVu8UCqBK6SofxrfOkdjK6
bFQ4nNCkbD/oE3AecfehNC93XaJvSDGg7zfc7b7D6j/ie1vUxj91xBBRG7JM
oz1nHFP1odPxo8TWEpVgagwEiQW65ikNcde0oclg5t+QdMihW6CKFOWQmOsI
Q1zQK2Wp9Seq4In+AywYZB4F+tJVL2kNO8pU6mDYcF/TxjwXLxXRLO3hLm4Y
omjcjAd9alP/cHAZhf7iCPvA319ecBe6mJM+OvsKMxxakeyM0zQWOMGzrfBw
tHJqRYOLGd/+2BDllgWbLYROyncGo7YvFngy+uKbOfUFG3/2teMeI74XvtOc
yvGuDuggBoS4dSnrrTBhdLMa+wTULKTPqL5J+bSHvVwO+qmcebHXpTCW6Psk
yO2zsYFA5pGXhC8ZAAKhCeFyvpSoo1TSalbvsji1fk5EmPVf/F3ycN5P8OKi
/g5nFXiAT/zBlTHjA0DOSzP72umDxz6muxdxIMxaIBdPJJrG4pK7+1bpQfJ/
qo2YwtCsv08MV2nbKpf8Cpu0fODOi0fWUpr2CdL1P85oKboesSOaH7hmeWQa
TPCEptOvRelSt7r8Yws8BQKoAYOMN7boVIEbaftF1G7C1QrKR1Vban/xlIjo
JXw/Jhu4WR0wTc3e5SPIsjAOyQ8qsdKv8UlYxuyyvYqPoQLVGu/TaNjczMaj
bRLPAgsutXffgQb8/qxyrDwIy02HM69nTaCdkQ6ES4LpbJw+MliHCf2LRAJF
rz6YsZq68qIIgUHiA5ckgWQTvPXde7iXpHE2OAJYBiIfwPvavIubwxTO0IwT
G72h7c3EmpOHRrcYi8yItWHo0Odm27Xo2Rkpqll84XEwHkBkrFvi5LHTJLO/
RvRvwHPblbvivWDsEC3TAtaxWr+jUroxBVQ+yXVDxAzMjr74RwGFSrgwzjMJ
LrlD2rT1t8iFrVRvkCiAOrVVvm49upKFVZhtypyxbDvC+CJQWAbg6yJj63M3
4OhpKE/hZtqAOE0wCAGuMIyEFtspeQqJfsaCuvtjyCMJY8Bc8/IjCeqqcMYG
/Duzo8d5GpZ53UjpmHPFqEowoj0ScfoOtWjliB2q+GL2i0a8m4U88wnJjHJX
e+PLsroxx4y30i5CJv6bX0TjuXUX3Ds84xsJdanWb5iYguJsSUXlD95uqopK
Fx1kq6J83JrD+I8/S7Rk6ZQUYoeztKU4CriZ4Bk08q671U2GhHNyCf2i7qKm
e1P+XCHBA3A8mQ1T7xrPlzlt8CQQ9j/Wwi4rmKBZWRTeDrnQRRT5rtB/wpb9
FJlZy9Qculov5BHHaocsyoVzHWpIyHHKbP5bpILXlt9ryiZhiOJX27vzkN5b
Q/IChD623UD6KcjdAMOWxE2euzTZhI9cqrTdwpIPfsx0hjBlWizmt+MrjTwD
/FkZMMFxDa5+MOHJSyVwYODnDecADC1sB2FmP7sou3srRBHjb9ee6lfrrRU6
ieWsUd/UKTgErxXJrdZ4VFzjzm1bCXBDSPb84sZufWYjy0Jxr9tvzwtMO1o8
kV6hAfN6mx0PhZVJ1QpVFHRHVbE93xmNcofgB1zKxuoWtkn1JboWiIvh+pND
ejxwjPhljLXQyl5Aj4Bt198gTZzZAb/a6+EqCn753m9A225zD3yJUMsy0Lvu
QUWIYTEJzXhjPn/u4EI0wKJ0Gd9naZ6bzp9iL7O/UreBCmBRIV6xd7xhIHve
KnKr8yqR1qems2ndUAbpFEAwiPZaZcNDaku71Yn3y672jLP4f0FwXaKbun0S
ecbvk4PB7BgZUbz4MdRVOzjghASTKXCPsDoFq2G/CfoXROhMyY41YxlHTdIY
SKwY7JYRub3GaKMSyQsDSItxA+CazbYby4UXHQWi663ggfGjaehWlQSy+JQj
k9tRaPZ9/nSpfsVvpew9AdvS81I0Vu5teXJirfNy7V+7zpf/tM84dzmIx+rK
lTGc6Qvasjnm31Umb47vy/08RldtMOZCq34lyfXO1cX80fdcedbbGz4N7okg
Ek3eNjegRvwdtulnwoSn24USDc9QJxcwz7NU4g2RyB222rnLZ+aKFNga2IqN
R2IJvE8h7s7Bqv8clv1rp7Lg2PcemkgCn49qzIM+e0OklBhalRLsJn3uVpHk
ye8Ivzz/iFGXutVzViBPo5WMPD+efGp/uGI5h7T9zLd5a3SwUiHMHnZL4QHy
LT24Xf+FIbeyhbi6welA4CR0AXwcxOUwmoIIo25w499fAy/wlsiNSPMWAH2o
bUayIPwE63886Dl2MMSLU0xf8Bso5H76wq46j0j61M4ABTE8gv1je5/lj7o4
IszoPrhJuVKnd37L6p0DWXumpRFhJaaIZ4EMQMIzYssZpckAUrVPwKkXmRUz
+EILkcTZB2zPaT+n5O9FjjsCguzCBAvyc/TtuYhc8XNDR0taTL5TtqXkCAxq
K1CjluYyW/qCrU8ysCdimYWjdYgyFX6UigoEVjE9O6wxfK9KvJCY7ofTnqgu
hkjA4VtgFjnOqw0h65YqeLUPEWw7/jCnxqR6/86Fo2KqCqb3T7wDnM6wDy6h
YutFiCTXTi+hClL6lUuW/PUMv9ksqfBnfXNrzsctUpxnHL+/KBejybtZiMpx
gopIjYcKbVV3rDqoglfjFNExeFhpZoZYGU6VL9VK5h9qC16869sCcF6xWqTy
GXlNjOtxme/yfMaCoDkZAtCjy78JasW/mgRUPo93Aya5KcVUPuvjJewa0n6U
5tnlFTlyxWeTwo9w5oKanMSUo4Op2NTjQAHYSmpRKHxGMlr9irqgfKp97q9X
VZLAmRbKYphKMtfHFi+vTvnGFlYcxhqeqLJ/h2JHsCGmtFMiMEr3c1rg5gjM
SZebZaau4zz/GbCCDKLXnaRl4RBobIia3iopN+GIx1UgVcuMW9hoz53h3nx9
YWxjVwqmmg9UhN/yRuUR0fvBCm5KboL74u5qdJ+z/9L2rUcy2Hk5o2HHqMA7
4LOGW03F10sZTkvQ1dTALyCmLl8kiknCsccvI0FSPbsl6Y4ipqPZSsLpuux3
rNZ6E+jZHFUyTF80IZoz/wlzyBC2SN4o4zTzZdT6y7ez4A2sfkeWkI9tcv1p
/gt3M0CmrK9Ly5yM7Wkip9kt8M4Vc2GoW0zt9h2tJq9Pg3+fbc1gc+Sqo7f6
ueKW9CqnHrxasm/9AENa9y1sxc06P9QcCB8sp0fi9nqd7z66D2NCsjXymZg+
e9u9rbzat/1gsLR1TsQogjJq9AQ8pDMkZq4MROeglszfUM19OOzhbGaxUH6a
Csw7YKZXij27npCzcdKOv4VSdQhfHbXUVdaJyv9n7URE+UGAd3Cj/S4onbPA
R/LFNVDfAAR5nKWuKk7h6eqTVmfUHdvJhHjW3rnbHPpFyY2G29CSOJa0e0Rw
yQMzfhacf7wE2Vit8YHFFoWyAt2LthURP8QjV5B/O3xtUSzExdmeYCDl00fd
i+LMP1lDs5R6EwDtqDLKh9kJivNtGF2Sy8MP9eoOUqBzlJ6TQ1bqJSGqGNRk
wqRVQ1cT5n9bH27Zx6sVcIxtVdxk7qna4HR5OGm0W6djY+07uJoeCMUCtrzN
bqX/MVxJhbah8iQbZaaKFCYWXSZDkTCuGrBXXlR4eAwaqOuXHYC2ayT4ZxQd
iIu6mSOBtZRFYOzklVbcQ9BfMNAUbqmvhCO+MiZbwydaqqQwdxGjKQZfCvxb
X4DbF0DMxgxh9Gu+ZtmowFzQ5e54l8SwSeR19wXiWfkG5Nv7BpBoEqQyYoyA
uSWKYPNqcjCisEvzd8lXiUnmZcW3B1GtMG4WBJvh4/1mMi8TONoFKP4GIJrg
KFFa/wX60fyldQeLfJ8AfNBPodcccw8Psz37dTd5gqCy6Wi0ait5CsgTXjQk
RmNZS2zOV9MVhYbRQQgwpwAXrIQekbR4FrzViEFMhXxLtcjQ1wh2hiwiqOcW
/+dFY3Udpos00Uypmi52RW7ct85QxCgXXCo9DHmSoeaHHzpVAvlGVs9tr9oH
HMnJkLaWWFyLM4/GXENyiNlroGOP+PbEiQdCB/S1kjTDaT2aALhnkS/ghEkI
BX5bRPndbxu0VV6hUYIGZJ6xQg1hj7pDy0ajuo+lH47RfBD8Vh84VzNUwcWX
YI9nXCxO4MNNypMwiM+XX814HYB03XutNUhjrKUqyU9U3LfX1LIIzclXRvA2
vdKNwLVzwgNmYup0r+hmj+lOeKEdWn+3WtUCEBoMTren66W2OrKjwmT0kjwb
Syl4ELGKG49jL6ZmNqqurRTW9LvH118ovkjNOREqIGut/Xg0FP+a6KwJVoU9
6lmj87m24OD9UBH0b0r8c6LK64nkcnU4vp3ANfYOsag64nzcgaWIrU4gAf39
7zclIfcDJ9WCNwwh8E1UNGZG1yDAwspZRu7Sv9jPrrexdVS2URlf9OqTeW5t
D9odwL8GRO4Jql6eo8A4N/aASZH4wVSX+E1uAJXzucRaDzoXIqLgyU05zpZA
rI6LA8tFGKuTwA4qmv6LDqp+IirJHVXpLHlxX29CYenI7hYH/PndOgdsp2w7
AzUzPviZ4dVN5TYE1Zk7MaAg7VUHyAzB+cvmjhxO7TAE64y6tHz4y2ILD4ql
Ey3Yd6nrsY+cFgPHpswbNnTiEksOPV6HjdT4PTpBtwCVAAx4YAk5NkAtGXpr
OJ37IumiJe2EoQ2IYBvZf+1xhqj1dGSbYSSCpc9SxI0GbHaVDyvJSSWjYqyX
8rXn0KyNmFgB6uS13MM29DvuxjSC8kiLjE6dumm7fGkUdgw6nOxekRQXefwA
vXCvFnWoPHpZc9mwxNMNTh+M+NCmCE0Q6ukQfwUpnlP9YQzuSyMEwUKtRRfJ
ZOR20eUHPvEMVVzCf472UkaoIkYJ78ct0mQjwc+PN+PYWCAQ5W05o9AvzkgV
jMuO4j0Po0Zhqkxrb/85uHOivMy54R8RA+2mZ2vaPa+27FNuwKK4tFagB/pR
A0FxsHY8LtNEURiSYZUj9l9ES1pdlK5PgGyoQ5zfCwsuRssKJEMS1mQjvGjX
0sShoVdv0n66whgETitxyaBQbOC4ga5Qa3H4KwK2YYRO9gvenDc+7Na1yzl5
nJ3gn2T2Dmvt6lrAqNuCjd1FfaPzGeJTwqdX58GeKdi144v+qwmjczgwqa7O
qUjzuqQQ3d3k6CT4d9VEnH3Gsx+70v/V/w+XQp68Na6bgdShZkixcEDtiOkW
r2v4QDelNUy5YKR+MRH1nL0p6wWwughYKPPJnwC7f9J4IqttuHXaK/+NVEyu
zi9DyuImYvSf6tihvo3xvyqzrDqkJD8C1zs7j+UIDumTvjAO05p7U8LruJU1
Dufp6Ic+l3JY4x1/TC3Gdttu3nlWiXiqDyFXTXGPCHqyjbXf3Tqz3q20Z2Z4
HIie7rjpA2LktT/a3wj9pl6Q0EwsQW9wRp8atvGZtSrozVCHAxWO1S5m5V8k
qaoEaVZFjyjZpjarUEC14jh8IEwhdvOXyWfg49/Z9+FOHFKv0kCndFsniQ1W
yre64v9+blAmibs7TDsx8zw26n+1j9D0BINnORURZCG2BE1DqZm+vxLIvyTq
IKVoe2fFFY5rqakXQ8Iq2dAa76L8/RtHa49j/D7npI06f82+3qNofQkPqYOV
eJo05Dyht2Q8dL6bJ34xHnXX41dMqTBeYg3mwP6CkinbXty9rnGgjd+fZV2K
q6xsVbpT6O2CwqQMrd/Uj8RN2+ixCmCvhdhWZStxPyVZDWzzGY931ATVGi6c
74LiRW+ooO8yftgh0e9zjXkS0siNqVgi3pQkT7dLZ+90Ma+5TlQSfprjooIN
l0WtXG7kUGUQe8jDQyB+BSUKh4Me/vIljzPlZWtakH9AhRGcKzjL8jrjApsk
GmJZzg1iMR+UHy3/ggiDG14MD+lmFTK+hff8Pw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mTn9v1Jvs2ikITbXnBUJtlRT7zrrsJOt2xY0WZN+wA5ww7PGm9pxZiIHSQ/CTdgJX9VW1ODTFYZq07khJ238y1iNf9zmW7T51Z93lpM/YfiDiaVnSpqzpRtDlS0WIxLXGF1HPEuydD2wbbKzI4IcwdLg0AlgTnLvcS4zXLGtg4Gkq3TITDwQObMrkjZQBati+0a7eAb3NJ+0aHJ8chrIs7OUfsZigmoyDA290kGgV/W3IOTHB4a+xOXt0+6Wafv8fZ4+7ZyBQP+N2bbWJSZGAtz+SaAS3xfNUtZyX0kZlClPzCH4UPJpFYN2JCpcvmbwtUn5vhqtCEk7UQoiohbDw3eQ6LNtkOY8GqbSzw++RqVHK/cEUZNu5iJbiioJTmZ+/wfNG/tJfgfSLRiJ29Uo1ska1b7KKoH0F0R2z7zlvX2KWDrtc0nqD8dVzzsJ4Ue1o1YxNSe9NED+Xx5nWrEtEwxMKGWrqKpUjORzQk8aAKpzWnc6VwfX1ebYkBkWOSsnumzNijgCxmDhVDZ7s/Sq89lpSYSlHq1z4/iWNk9i0FWx8Qtlj/qHzshtpXJ0o5M49Da9/Lg+s5oS/YhRZhB0z2PuLdh1a/K1qpxTikkJRJCv4jvM+9DEH1C4L36+IUf6sI7Ano9HKCwZHi9GFFezZIHBwZNYBfodY+LCMzpJCrAEiiw+7HyOs2csfHVb0aVzafm8UoBqle8LJZvz5KbSqjQBqUNpFo7LosvhKZvYuRmquRxoooZ6zlKN6MaNOHAyYnelKvYOttjqogfnFMcetl"
`endif