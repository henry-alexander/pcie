// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lXdkMWheTTmdSsaiCG+Go8kIHTQ6ga8wP7oaS/M1ktA+5E2fuqUOdELdF4TC
ivA7D8g58jgl3IPzc2QCRogAHPx8iXiQvMCtBcyKgFN/uU6s1ecsRuPKldjz
ZckTzUh9pR4AsdIlpUluVt/qWWjXs1MTN3GJvFPBas8r1r1dUiuV2JWjOmQO
ozTE6hUqPZIL6BguCMlhLnvMI3w3uy2gqdOEibF0dhbxVwNoxmVpUnmeTjmA
/FRSeRVZSUlxalrqTq5KqvPlhbWzu0jbM1S5uwarqtQXQBpldWS9SqyucDHU
1vcKT8LMG/D/J0pulNNYJHo4n3uxfhuevLgyKRR1Yw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CbsT2t/2tFvvNncaKYFxxIxD8RIK+Gjkw4y8+ZHTNZ+UdAxDhHaeQ93PnykY
mL58HawxcaW4wZH59ByhflUsKwqwvZzU7fY6Vzn6hAMLWGqch6Yy/Y6P221t
U8+ADi4kd4pP4qkaDTsR1peOXJFzq+ztFol3Sh6BqY8RLP2fibkQw5CysNEU
qn1eM5ufiEj2eqE0moxbOuzLJcxJrkLYUE+/Nmyp4l2qkGZ8dNy+bqytIZWg
/D31CfoX0M1IEWaBIIhEsCsx7yOisETwzAq46Gcqy70SnkHCDgSOpjqf7pw3
lJ7RYrz1dvwidtl3spaFFkx9+VW958e7mt6tmB1S0Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qhoxmIpeK3y7uH+8WZmizjFDt7wOTQzcth78Sd6rqs5Ei4oSSs1LYxmtFYUy
QiKH3V1xXhdsxxBKGRx/KGVg0UqInC32NFWQPYqu0B81DeMqmG8CWF9iVF2i
/1q/RWvxDM0KzRK/Tk4lr84iGw1KUHCWrOhv3OdV8Ym4tqKfufETX1ZYvbDm
7Lhs1lsTGUqxlhVTXCxLSU2Xh5hZ1e3uv8kmsId8BoGlQGhlQiqz3zU+XWx7
5akgaxRSyDV5aEMkb/jLpK/ax/9P2WT6SGf4bXF5kZV46FtOQnkAE8slDor0
CUmhYH28qV+CRUcwRxr8CvglwFzRhirM4ufNM9MqsA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BlHwVyPT6KDzCjIGi5P8dAkn3POAVgyu+ux2iZzlUwmdqsyOLIbWdInLwliA
FMYq02nEDuNtMqfO57wdepj16Ruq5CszEZL66LcsXmAMH9h95rOaoWRVfpBe
LpizwlB+AhwcWl8XIKVYIsw9TtTMD8Hmori0jvvmv4gsJmAmNNw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DjuRDRYUVDG0F9psJAWFFvGUCmiIJSth4HGV/Jk7ORigLPv5IQbyfFTjg4fi
u7RL/rYANG1QVMrSfA7wer6hKmy1wBlY3uden/OGzwlmVhen67sOddZCx5pw
aGlROH5Vi7U0y54SPoggb6rBdmZgpDqlCAHYSGS+cerdMSf6rUB/4dCRRIor
7LDHSdZ3acz9y4KX0XjmZsMixhwOdGx7DvgLpYJLaxP2ck9Jiuag4cO40tsn
6VV+RWQCp9nYeL7p+KsmPy9pqt13nc08HPX/f7+AY0lxmYhSntAvuUQZDTZN
EixpYlsqI03sehpGjWYpEDn74l0rmsqwerewhB/FsorNLJ01D6fs2FU//JVz
RH4Y+yN8bpA3Z4y87QjTBb8bcB+sW+0tIA/jDdpnpHe8klVoDGf9lBORhR6A
QRgnRwktcl+15j1ulFQ7I3x1qHkp4auLldE4xHGBwG3h7bWp7TBXQCn0GzZR
1vJNpiRG3iaksR/IvDWLNWhX8Sh53R9A


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NA4Taz5oyrjvTSHJESongzJ9Pmst9SKTudoUx2nzvFO5PpsbcF5sfvSprWWx
00DhYuoQC6L/b5c2dA+KuKpI+xlPO/sbg5lYrClb/9WTaenGsAGq8O3IOCLV
FoOPoIbmWVjp5mCIYOlDo2KN4/2+twN0EPLn9aytVS0sNfQcC3Q=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Q574Oza+y59uLXwHoGxEHFt4FiSKtsd2SAHDH83NIvpDk24ErEKIayPZUfvv
D1ULLDI3ZQCLile+isjyldyVLiwryP2v0aSmy02exdeIX575xAkl5mkA2j5C
kAfrAdKvFeRTQvYDZTnM+0zMRQ1Lm8S7nZ4P/PN0yXDWsrtbxj8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 28672)
`pragma protect data_block
NGun9D5+GahIug4bdYmQkluRWyIjcaz9nl6XRIpZUe9LpKQ1sckPT1cVPcKe
zeSAZQadcgREeUREtxXiCRXUC9+UBMZwC0YFScLpv21ATCQP1FLu/pO70rPD
CAF/WxbzFynjPQ8drtDxG5BZ3msnjJh/D5Dzxt37CEHqQYG4SG6KQFJjY/Dq
cDv89q5ytksrmRxqcZXIzRwbOnLNRnefUpLH9ACK9XWHr4iF9T7j2rUX5i9w
X+uJcUMLtNMR1JxBcDrUbDZk1Ppp205oB46SUV0NVtFE5QHtAMewGVWj2Wdq
Qkl8mOVxW8Ft3OQlDy3iXFzsz2JLEFmR0uGT9pe1Fn8KBuOz6M9nuHZvdG6u
1H0ZbNoYmM2Cfg4DNJCS5WNP/6haVEvgNfxF1beAqj9cbk+E1bZKnXI3JEkD
i2Y14RMvfq4miih8CZDsLoBdunk4sCge9P3/rNC55DuUZ+owB1oqkdYQixt5
LLt6VRBXDS5Aw/iV0mqcEAygjolzrc17BiJH2q6UWDDt7LVVT+MWnejVsywu
b8AsXx3WOA9OWB+ocJhJz/3zs9W6yeY/pHfSbgLj0GLGPclihFI9CF/AHXlz
Dh5MRwwdegwqjvIicd+k5KhI4eFoRxSsnt6jy/nqZ+1xpek43G5sIt1/KayX
QlFRG+UgxeLca2Vf5iMfPEOKfoL3W7zB/BcFoc8AQskutS85MHAtHhlSWFxY
24RfZchzZ8mFk1f/om3Hb/vVWvidvve40zoA2s3XfjF0YwvtbG5ctXOl19CR
s2Ssqc+WtgXnwcvnvlVoFUdMCPbLqa3agw5s0Q3FD+AUuqwjpS7H20zmAjvO
SYb4lwcWsiQgLG1XN7Py2F57KGgObwaloEGaedeewIXmCT9hVFCyE1/DrRal
9qVkebvEO0B73AJfE99gW3KKCtRYWxvB1bg0pVor0xQJRDrdcZL8mo85d7qR
uTgIhqiY9ZlKyHLKgxbFmNcoBmbG+/N1c4BgyqovS82DuaIZ1igxAJYgWRI6
R2na8nVHdaFbW9Www8l07YGwh9FZts/xlsqt+vjFviuM3qFavzphkyTovnbl
y3gOBiHPIkkMJCBI9JxZefrwHGAV51aH8M863gUTYST6uiMVBBy43+4PT1w3
NYFI3bjHmmpa6Gtpga3sKrnX6WMZfwgWP67Hb2JUiMeA1n/PtmZr8aFf172F
gZzjniz3biJvXa2GwYYt3lup7Om86iUfxqhaSHmtKENcsHJWkNhJQnhwC2rB
F5074z2WxSUc+dj4QoeWpQFAoHisHFuljPXcfFvl10p3yWxBbPyq3nfeDJA1
KLz1cmxOiA52hmGjIu6CiT6JmtiDLNQ8c/JrlTnQBZ0GfBaQ6x+985ass0EW
WYj1aO9HoNOojVol/sWEDHFEQl3Bti8xHDCfH0Rsf0hs6843Z25H29f3aXTM
M8PokOYiA0MOyHEeqC865ZQgoGuQHxYrys9NrtO/oNCDOSWr393J6ekO1NLV
bwfBZDj7liq1eMvADgkaYbHZWs/R8A0DrhgoYAe3BY5/0oaqX6yXrpSqi3vz
QqCQp90nou8BTXnYLcqvqKIc24hoaDImiyhJE3ZI0lyFmOwFdBczh6TGg0SR
DdwoS8A8YV72A2m7GHomIirqg6niuYzrOzS3F3qXOkBpwkGwj2BtlzlpU9bY
sL9ggE/9kuoIY0UPbmxoRB16/MoLAPpNfuPuugzDxgG7DkR4wp8fIeFQlZ8f
hEaNVQ0LJl84xPssYXfzcf6afE9sH2XfGp1Wi3nN/CmKrtA22aZgEl0wbSAS
gtLYdORl89knDYbEakrnFQTC7ofEQZQ+8c0zPHeUHh3Ex1oXlHuirwbjTqMz
4UqDa1ja75KKiT3nZddTmCgHJHaIS5SPz1GmzXxGCYXHtsm4nqUANSDBxgAK
fHJjNbexSoNAecYovcXZDtoHUs4wai1qKlthoy+uqIRTv3myH7jzc3aWmMHY
lFMLpYis19FzgbpiCk47B5cjjPsMS5sMuYLGShmfmlLcvDwKtn8u1GvFQXgY
ML1It3tIP11nbPZ2nDXOsba5eBXjgBcXq4ZVgiXSHVgTPe9ZAdsbPxWutxIy
qAsoUpom6bNmaEmpEMkxxTWWqPsBuU6wSPKldUH5MpP+rvkeI0BouJFuHQX9
oYlrR3LcyeaPnQBe9NlDZI9v35X2eMkgRT6YDmTWSeHICPAB/MjKBOFNEy2H
ni6scReTZhVOD69GgZXlUfpKHOXeCgWgIJDvRRdGGkAzn+7oFaE/4YZgx3To
UZ62dMBODDcN8a8I0pPXv4FBfiqixluQEzYChwuXKPUELdzThgHXn+RKwsau
1/YDVD6QEffYPMfSfF1DEzg/KHDHUlh/vY7s4r0skLRl03yz0P75/9WbHd0E
XZcZBzV0LOMkCalcolbHjL7eAw9n86Rs3AW7Kdyf1Sqg+sBluYQwbqUMw8ys
T9xdBaycpHALiH/tsb3ysGGgkdwJP5A9xdvRbEnE/ryd6G81cXMfnlUEQVUO
7XjljrTaR9MOGMu8/eVeuhizs78hWVsfEUXWK8I8fhf0D1K9zJCCgfVKnLja
lx8axmu5kgGvhJ+tCsx4vlZBHpXMId3jb90GpFVQ/pWeq5dWWLkz6U+JH5Qj
nGil/3BbmQEkpopAStuuop3jtFttgmsLQlg3vnq/t3WTzmDg+5q9tLblWCQf
noE3jcqJx8kT4Gx1co3B5+j2U6cUb6llWeLvqujyzzJE4b4tRGpla61G1oPC
Xf4E2PJhQA1Wd9B+Nw2/AqOIgqzTqLTWnwi45XyOJz8WkvyXWx59Vxf0dd7s
KodfilfOPPBV0ME8tN5w1KGz+AWZcP/JHvirAcWvd1mBj1+/ndhDtukhL17O
3yn8EYT3Vlo/AcG1nLQz2WrT0LShv++Y687ZzJZkF8Mbj46gKFniuwDaTZX2
Yqka3lNIGbJw3iyXwu/IuWeZJln226uY7ES3uTDIcXDq4evE1eHT2GzzPrHg
MxnPfTwck+dX97sZ+lBIjN3MULlnOPcutiHZ2nwlvNA6L67o2X+Q3dYcnv8b
FEBsFhXKF6efHBmqJ8ksb/EInmu+HnspupQmlx+Uy4UXExapJl1IfZqhQJ/j
z0Aej9o6BMCRwxaHccNBiM/RSvL2bIFjOzv1vtDHg81HqYl32h/ifvUvLzXy
6VJghfq15DMLEgpGdH+j4w84XnzwS9wLbWZZfT/Wko2A2zzs4nKhScHJGNlL
CFP7BaQWKf0GHuIMizNkm+HNSO1ne5BvmYOiMv/5S2YhEOLeCjO4ui6HwhZM
8PtWTWFXL1SfkhGvGIw6gOeFaR1zOF+midoJqIY7XLXzk6BJI/fQpdIB18Z2
M5Nl2X9dZEen9XBMQbOAtbJZb6hKFQCdHnhav/iTLzSHCvVJFlbY7N/KE4XB
LqAveVPfAUbsAxlQLQ0Z4NJ5bNZg03HH2tY9hLFO+RKgpyxzzvtSbcsz7qwZ
WsXWU/yDawGxKbBl/pkoVmZIHxH/jQwjMDhF/n8Vz1+dosS+WA5Oap7NF3U6
ftcANa+QEWsKcjvmg1/GTXx4y+vUgm1yxaavRjG3KSpdrvlISlEyDqKyOq+I
e2x3SOk0PvOxoram3eTPeETEguyN+u1THnGiZYxteQ5aqq7B4gtKDuKfAEe0
ucUuulD26sWnCT7iynD9ICcyJDX4ymhb815lGBzaCgn6idDgVlgfj68bT6Ey
G12CDhJ2NYPdsJAwswaJqb18fYYqTquBxoZU5h3FVIO5n9bD7REaeqe+mnKy
UFrtyNlbm7bBCcJU/K5RipMWu5KabqJKIoGU6VHIswrq9cE9G6Lknyj6hHx2
WljLrNBBkO97weEwQTNYdAiFbJkQKG5ZUIMUEsit5sC4vUL8+c1XBQy6sIJz
WzrotwC/8jgK0GmYhXAC+jvgoQtPg/AkppBTltLZx0Jm+SRN3YDhJ+4qcB04
MaA4Fq4sNwQcbReLiqUHoFkBiGryGWCKNbRqYAJ84yXB0sNwzGrigNuAos6u
FDPLLag+EojXv45MXIYEhnDGggCJvarAK0dprCuifOd6/NY/r3IpeL4OwKir
sytlHhXH8KVDDZ3j2GAkPPNJEGUw/rfd6tCfyGZEOfhKjNgI2SejkDRUmW5N
EO1qSGtCycm1oIZsWS0ogcrRdGz1xwhNaWlsGnDwh4mAm1bDtoYjr4kiP8xw
KKXD73ZFKsnL3VKbV4NMN3dEuQOZLIP8IM3t+YCfLPxpyw3PyhhfuJSz/z8n
+TgM6pLvQ05lqOXDnqevsO+sgM4qbNEqYhc16BeQDnRZliBvvVhmdFt6n0yM
jYQ2n1GuQMf/+8BB5BYDbXueJS0w6LQCiF2YZYSkYvSsw/jMTct5i08zS2KS
DlTvKAmYFFs/RXxwdAazRD9Qui5xbCS/d9nK8RYNX2ZtjR18yAi7sEnAzLpD
9+ICDCreNDRRYtsaY2GsPurUtVQSEC5G7CadHW847E0qQgmz3LRFd4BJtZ/G
DpmLVPncCFEjr3i/1jgxoda8jFGSfzvZn/I6Ddu+wyxQwn7HI9vML0MoHzXl
f6mWw1ZGZ2p6YY/cSe/txdRnUY0A/H8qrYrM77E4WrU8K4/n9CXHzsoNi2E3
sKIa842Qz79WHn8R0teFK+6OSbprOb7STmEt60VvnZcV+PCTRI3QbMNz0arc
fvWfcBGj+mbxE8ApfxLA+1a6SwZqu3ZzE5vbyLowOvIw7NnTowukzS+TNTRB
m/t1R4VuscRfaEaw3CCD6rE45A5ukEqZ9UB0TufCVPH4V/TCaVUHimqaYHJ/
PuNvqFsIodDD3dNShSmFTB5T+X4iFkzlSRXml1yywvacm6HYdwpdyGUirq0w
jcPR9mcqvN+wCF35J8vLtgDqxXBzML1PS8VtLGXXeWuYCrkN/NySrjS+Te86
oOq2Tnzlglw6nOceCZr0cA0WpE0bRMjGXUTovMT2DhEnR+wxngk0mKLsGZvt
Af/qGXFY3QE2GmM7ZQXDDmsIWKQj3tCxfNNGK59AqmFgWj9RhjTPuREy8QMJ
+Yv8xsiFm+YFcmPQ0etfZBlU/xNIcfqIM4piW99dEPjWsMgl5DBN/vo+KDf5
dhaE4GmH+GbC9gL9tQ5AdPZvJP/5L3dthp9T9krnC7vl8h261TQwLHOhyr95
tFl6VTl+uRE674puBENFYHpCvLeqEplilw+WTMHWpl5J0HBOr+O4jCTM5w/Z
Uj743ebuL5V/UPsRPvYkjAm0WaPiz798+9Czue91B5L/xSyRkMutFvBhw6HK
qBX4YRkC3h3/2GDlZoop3/xeXQHUX66Hv8LFm9XU7Pup871KZy4wXUDM+z/u
Gzq63gOqnjDQp8JyaqxSn9BVkaW67d5O0ISjqH28uWrzP43R+QgU2aieVmzy
NbKYownV3tv5s9nrZOqz7QkiYD0wDFvPYp7+/OTKZqbkw+RS9yEnsXkHmTBk
VkP3p35wZapqzn8U0OfJZFkmi9lPmPfqRw5qiA3hrrmy57NjQg0rdmFp64xO
wAFwWMS3QpW4b/8DQ0g2xRVZhS2WHiBeUTsCIM9R5VyTzNVBqUlP6IjGyUt4
wYW2zPZfkrCfkNFmGrnl/A4088z2Tofh8cp8DTtkVtohySvtw0zulYMJIVLe
qGhEcIn6J2+XohnSi35fQqxOJ15MBorDKsM/lI8izeaC5hRVbYgFNnd1dVtO
ljrwKogILdhaJfI4WXRCejzb0Nys3sh6DTe0M41CHHRgAiLlBD8b/X0w0BSj
4/MAYaLjAToOAfT4xAD2hAX0NBUoeh1UF8mUVtZljOanp8AVWy34xPeRsac7
9Nu2nVfDrZEzn3mMcApnYTkb+6OP74z8ufWCAU0LHhhiOHdFPtVkqH71pXIw
0ZCZQ7rO/G6II18gkii92q0JvnasjqfjU9KA60pAPdrhX15dH6MoVocXoxOg
Ao61NzjjsGlAxgyMLpJnFVotsSL8ebnAyP7gqvYzJ9a7I8fkaSmMw4htBC5I
hAPocw8skZFVN3locE6wwE0sWHksCHpKAFNK9M8gzdC7594TBevxbIVelb7p
xS6kVLhGSK6DHRffTWNpAwfpVFv0aVL1ywFQQU+IhouL76Hvf3BAUINhx5XO
cr6mhUSjxHcAHllkDXSGpidDIfv0+rhkhNyp9FuzzW2whrBP4fCJmnx3y432
Ro5BYjwOkEBiBO0T7bMe0Ufp04JUGrTagIi4IXnd1lk/8MGmAMddR/QnXy8q
sFpwxACxzaaDNUjpdZbC3m4qcB14SHbjilP78+Sx9AbrVy7rj2yBjZw6mMTh
cTrjmU2WQuexudnvFWI7XjYtRPJYqpGegY5vvLTPnc9PR3TRsu/zVSG4BRDT
FvO4Om2oQKOlpiZ8T6NiAzE1Gg9IqloWwLFZ0LegPEf6yEyG67bkyu33C4Ur
dVBos2J7YmbI4hMwDfcErrqcXbIvl8OlNvlyRWEPC7dEJbOUYfN4f0sn4kO7
CfiEZ4lYaiMytZAOD6CbNPYpQjwT4WvNEaNRlfNVs+macY3x6+osSqzd8WH6
INVC4U78EPK6pNgC1fxsT4JjPThKTjJGniRVdhfZq7M/3kkhqOYGeNqWpZOJ
+9OBLmAxxu0OTxr0f8DvTqd2bygT6z3RFIUIszLKpMWGpSuWBklUuTHGeVWj
1XVe3awQjKq7soKYh2FkdsfPAMpogwbDQ15K3dtJulcfoWBUkDTRLVh80jjf
G/qR3+gkQkWi2bpekxDmoV+E0KCaF5HLlAJK/Fc+6F84oCMfKNl/8SUs0ULS
XmZYt6HxYs40MfaKvY/rEz9w5Zwqg0S6mCI9Uq7Z0HYABQA1RoPUz7RdDQH6
XooUjcHGUd9uuWXtqDY8G1R+Xc7Zsog+H717e7c9ZXPromgxHaQLP/s0tdlc
2rmJprLDe2LHJdB8q8u3hvQojXpKcfNboNTm4hSYT9IX/NJUjrvfQUIG/Mwz
YrrVOsBWfWB2HzVT7hnrWmghYd1w5MFWD4LFcxleqjmaAqqzf5UL7SgeEOOp
5MKo6jsHCHDKSRQWDWaAVQrDgkE2zZ4ZsF6TNQ7z4G0HRvM0lQXka6GgwLAJ
9OjLiDSmksQc0sRz2kxOChNPn+I14lmqwtW2694+xru996b+9sPgFm1tpyxa
/E8y5ElfWIj1bwFaRM5VjwthhVE8Zh48gaPsGke1IK1m1a4ccdtaD0kvbVMP
lheLWGTWej61Cho26HT/OMouAllEV6kqpiXscVejlmXOWKhnJNWxPFTQP/Ez
B0LF21JUbzc8UuXa7KVGI9BRq/jBOPU1Vm4VQ0cg/3p/txMcL7/DyZdu+21q
kzS2uWWUttBLiQcR6BaIbwzLpDosnLXwXqMMsNkDU7VI7HrQcvTN4U30L6Wl
QsUmZvzan+lMVahpfpHt7tIMZxMK8xFqzm3iMgpcmjj4glB1kGPvkoDpt2gF
b1d91Cl/67H2qRgQYcX1qkOYBLqi934ol8+JZMUOOzusJJayLn5i5KZnmd9p
4n+iTvz6OHKmBc7axN45gduJxyywygeNuE/VJoj5ksSnTocgb9Zmus/9j+vl
8icXNmh0qjhAILQ6Aab5LN/YWPqLHwCwFVMih0esMTgRyNKOxJ8SvEov49Sb
929KYbNOzZvKSK9pHoE150109Sj6/YmOIYzZ2WS1WuJ6NavCq256PAn8+ATb
O40VMyfAtcLS75tneHsPRFQjbzg/bm5mQl2mZAceN8PDcMsm3a+fHsNy7lJz
V3ve7FsYFiJjg7sx0WQz7FthfVOcNfphE8wiVz3vjEqZJMsnfhv7O8efIteI
xGnsaFeAuayVhj+9C0RgbD1pALbbvrFSx1kCvjZjqpOcgU7g6JlBRZ1wLp/V
Xp3z7zrJtzUj0D2m17t5Z0Pc3t8vrBdOetvRsFO41n9b+RNHVtL++1zrAeLi
blBX3ilGpFt0hQc+UIj5vIJ+MlwSE8nGCJ0RCaaIoHbYZ+ibbZxcmZT+bf7O
R/r1I1vyGqGS/7x490oPk1RNaL9tC64ame3P6sJwbSCqL5aLBzqWt4PI4gNY
VGOgXcPwfNZgjKuOK67zm9vpQT6GFbOvF0iLDimdpWuBDdQpegtWVXPVTyZL
nmJFtMDoG41xY/47f7qy7D+yWr5bT+2PSE0O7a/y9tyLGqJOmTjxxLBo6Yi2
sHA2ljMEoQwSfi3uXOpLV5VPt7Iawprvin8gdquA7IsDMnuKh5Snl6R1uqeX
9Z8PasYCMYEO3CE9dgCiZtMyvtazjQ2heeyFzEKkjeob9eBSHhc+ZyMNsFQ/
ThMUH/NQFVbk88J1mQDrHO622DmM0pICBAp3NYEpDiS55lTmzltHSX4qaL4v
VSNviyw7PVTxygzyxAuVV/prYlcBVqUuJhNyMAYMwpz2TG4gCSIBBuJWydyU
1YH5eGgmdmQZaLhm4QDyVoUD3ggjGZn7rWZkInlySJnqhcgHgvsRqLSiQh+5
P9u0jx5fh7cSxJfgqjVBWUItmEoCJaOO3Cr1oNwTe3jFbbz41Tu6KswYZtem
ArNAI2dl7E7ZJs+BlkvrmrobRqI8Ml+CupzwdMjIZ0Pb6oUPjv+iRdyAsW/3
g/m9BMFKihdXfTS5jTgk3wcxgXlzR88SFTH82O7aML/je6/uj/xx+BkJZyv8
wbdavcEomg5Tm5Nurf88J7FmbZSIkh5hrUnGuF0LAzBJ+0MkobGI1S9sv1gN
4oiA081716arSN+dsSnAZA7OzRL2/HSM7YoO+DBM8fNhqzJT0ff5N4YMh7jd
cccLKnUACBkUM3eY2P2N94V51xdkwt4YWydNVL9V2VxA6I3epcP/YgxpaFud
a9ZP9tcwSASQDLlttuNKYKVJ+vuBcAs7gMYl5EpOg3akIQ5WWySi56eg6K2Q
ClGUAGHtcrg9IJ9KtT1Jf9h6fP2FMd72xZrUA0WnbLhsVLPnvivsBk43zE4T
s/v6N2tV+JHUrrKL0gjOGHsrfvIPNt7UE/jQ1c8UZJl0VSD0XLmmsEdZNiMp
a3mny3cRLSqo6rnAo+VuKa8Daq9D+UYBeWLmFBuc9I8hqxSDZXRJXW8tC4oJ
1eIkOXQ8+8FhZYduZuCHs87oKZuIa85QjS0JVTmsLs3126RzQ2ewEcFN+M2J
0RUfeYj/SfxlU+ywbg5jgnixiei/EPSOHgJexjON8eOAwf2sGuy+Z2/GDSjj
BXAF7ZDkGa3zCj85BjYOFBbb6uWQph6i1zZlC2626MYhLgidzR8iuC5F45qL
n6lWCzK5w6HNY3x36X14SyDvnD+zFwAalxK0kfvID8HA3clZtTv/X+YgNP3w
/VaUrkxE1VF69Q2jCYi7xV8ktT567Gl6QC+hID4JluNtGgCDRTtWAonIC9ju
h76ASBOO/ZGjCRC+lJ5XIqCsuNfh3fCZjFEwKWMeRGFyKkX1V7XuggFNBEna
ZzfoQRMcFRmEFtWWAaRDVVSLvyHPWA/vpugDnadnVb4V8G4rbv1I3GsyDjXL
YBoSF07O6MaHNRJ/b+JGOfgtO4AGkHL4tI29B4mCZBBa4MfJIYQfes/sQ6s+
4dSYnK+e8SHKTEvm0xiKMxMXs8HMqXzwXqA3fh5okPUVTP9T+GrJkcHTeQZa
G9dr8MsmE/I1J2hjQcxSENdukxOKsHgIfc+rPF5sD1Y8Fvq5DwnI/x0Hdrt4
659PrZ+fvEX+VNdLwCv8ItKh2+IMfFDGVIxt3FpR18SoR7se6c04RTiNgrFX
trp+b/TmFKlbHiN6/GjyvrIyN3TnwEXsqIY0hC999cqhNvB5eQP8QiGIUgIB
zXeTxoNPr5g1uLBzeS6Ck1F2AgjRwLDvtuGgiCmwT7ZqSw9fWnGObCBsNiGg
ezN1jlfC4RNRqvnEt7QsqvsvadbfF1nTSXBVnYzFedwhpQZc2aGC4Z0Gk1ai
3eLsNXiUdywcVz7KsBIZ/MPpOu0SMnwsrrxFMyXzjG7qZ7qDL3ehdU88Dqpy
mASpTdmtUj+C4mgKS4K5Ky/d5oYgMpPNrGyzyEsf/HKz6UHmoFQaZLmHHHI6
3xgYadmNQAnBM3KQMOWhr41j0n/x1s6J78glI1rVZSEGwQWuTGlVgR3COjzP
hDYzm+ssbQDiXturHzf1n5qg/on+oDgk7K+cJoUcYdmXpQBC4eyMks7hnGae
J8ewEjaH2K5iKrIcx36Ol4YbFFSdDQ2W/+AlJgVR/fvQrzcx8jbIHqtZQkJG
QlQLMt1DqTHi0ySVSSwNsI6X4i5SqDX6P/0tE2tUVHJOVPO3Fj9IykogVqxc
oGL7h0C+850LCnTzZbyuY6TrvYe1t2ZP3ZYQb6h88sBCgzT1Q2oO5PRewF6z
5vb69Sx+66jxzRSlJHHE4wB7IpntpfJacnJwgfKntuQyxCfP5b6BTA9FMksh
zdlRbX/NbBa/opVEgW6rU7GGvhv5zwl4r1CCIMkX/1lw34K6mZeHFMI9xXH6
ylSdX0q3JgXM15uTaqAurEYp97lg3ZeHhoT1hNtfX24yqbESYheWpvgK8DZw
fcz7ODtQmT2FQl1Ny48UytshjAo9Qf1YNnTI/L3O9JSp4jUo8pygpXSrqTvJ
nibB71vGwoapNnSZM4PMnyKukuRwpWnKwMtMT/PiywFeaOAp21nbe7UbJ+t9
E8djejsTtWzJFMD7ilgF2SgzCfgKOoYlmyWIsiczVAK6QhAR+nv+/HgO3h4N
pS35NP6jW0qPwEDtCds0SS0uMJgqpDAGOL+3OX2fCG+iPfwVRctLnLEBSCxj
VnDGwB6o4yaQNMjkdeupf3cLIGfm86Jh4XJX6lai8eL6QGF7m8pstlzoi+Jf
YPVarCpCejuxD2mF4xN2FQ8kXwaqRI5nhyiq9RlEpvQMdMu/0T458lNT0Yu0
l+sgxDpOmAImCjFkR2Zq2VFajmlx+v8vtd0KASsi2UX5s/02MnsIXvbd9SuL
n6WY6+TWZcHKDVQlYjNUtDj5nW/jxgsSWeR3UpsGEYM1CRV7ILGlehzgpuQe
WLN73UATizGY9kyzhnIZ/LzKIdOXve/OgoPbsUO6ZU7eYstWJBWzGiT/Lx2x
we5FnqrEhsD8FILfgIzm6U8wIV6w/UrtXHa/nAphOUxLFVTbbfXQed9a1LC2
X/SYLWDFlw2GjDUJgXVzeKaRj3kgDpy+4DNSXUT0iDa/gZ/t40bEg6iCgjsY
gwJ4ZCO9H6VOJTnV4Xso3kdEAsPKCQO1t30fhQ9i4sYQwMUxdBQsG8/Sd76I
BImF3jb2HOW2F6HABlLO8xGaX777Wt3sm7+HKBW54/X4bYJeLGd0kWagep+U
fgJZDAyNrCLekjTaulmeGz3YZL+ymJojV94TBHaoOtNjq/dAEK+c1v2UgaB3
BEhdnlSJMvox/TnWI0sXHp/0XQsOsmYXqdjsQV45oUNEIWn5iHClAfrk4Y2/
K+p+WNDYWpV/RrAJsiF3XGjCo+nIFCD10s4QBNvyaAHaIGwoJX3PYgpS1Q/t
R/nNbRFLHgnNmd7S0NRubFFwIG2YeLISyRAD4QZG9p6OozbdrqbBLZ1S2rGh
Y+T++fl3uXf9vjGWf2jl2x84ipdbSq2L1wZQyZVNBmlEbt6LVEi7mOlpMXDV
AKFXoEq3V4rPbzdhXzAYbsvQ0PTgIlR9jMrByLvnN5pSTgLcsskh3c94/fQS
F0gu63Ffg5nus74fy601Hdx8onYKgSX51UScWeH7VIJU40nTlTNK6/azNbsj
Z3jTyVfs1m6vPoVHirSNyjjVALdZtUCHxBnLIvYlP49Oh261gq3abocY7aZ6
4wYT9HQFqJ8dk45AqynJ9XvnxLDyBb96NHjeGV6L/g2qtU+CBJovNr54zGzT
CM2X8C1Q00oCD93qFuo/wh6DShfHuh9/uvG2wJ1USh604A0r7Zopeg3eqh8g
m6n7EPrHBSwZfzID47VpTD8y4PlUO0Gw7a3xZ+94Wxvdj/Ef/SrGST4OWK3G
6j6MbnFa4Z0dmLYs55P1+c/lhjEoEeugFaGDl3wsDK0rZeLnWQ5//gEZR6kM
b8wnkuoLInysNWUchW5+XPHXIHS7vgsoxgDY8MbxbAJrFDRpy7b6HW0wba/6
Hc3Tq8j+eBGvx4OfR0OfzXWpIHPtVIlTu1pvPyyViruzgaDA6hmA4P+UccmS
gVmZfhLCFp1Dn/vw7y50cE+0eYmm6r11l/6aLNl0FKXujw/BzpCYh2wWSdD5
rpzIo1k5V3OgZe4dLUKOyscqs5tHXMGkJHpXIQgO5s/15QUiXsnE4dMsnK49
J7z3Un+ddl4hxFLfp1Qs8Noh6MM7T3xCSoMNTYGlUHWUQxnUidX5gPluQjoV
mpAhOehrE8FxS8h+9eHJUu+kR0fHJKU+87YlQgoN2whVj/CE2lqOWux3qeo5
UjLdbxSVqjAvOVtlrxaHlNDX457TAP9vOB1tAwCkyIe81kaS2uH+D5IpvCij
XNiL8GUf95OaCRR4ehKNYHWErueap7Lqr1lBPGvvrmP4zsm/0o9GmxNxWzFy
uf5pJmYEubXQBOHHv+I+OkLKNdWTURhkciH4ehHl9LKyG+kL4hajGt3VtNYi
9s8Nz3qM1wXCngl87Wf3IMjjOb+IfK3pf3QXvOKLEXQN8e1MtvunoYE3K4tP
0jVS5YGbzNBtrQ1q22k0xw6gR2/ULeUhmOL/ybc6OigE+MOJG6102F2yyYt0
A3uFb7vzPT0uFOmjp/LBlULsIi+ZH8mL0BOTApA6TgJo3/WU4TRXHk8MOzi+
gUPNE8dpsTBk+lF4sYDh+e53UU4Pt+tvGBOI2Ri1Q7pdAp8WVSG17QYXYVm9
UbMhJwwJ1VxuK43ttCk/wkcN09KdLZD8SLlbebrupr0S3sDdKbGqOGCfhX4U
EQ4IHa8gxsGQib2aYTvhD5gmIUoVBWEJOTmoLVi+r5JC0xib4ZpdUPq2Tb8n
sMjf2D1BeL4C9K9eBgNq2DW0nCUzN4Hhph2JT1c//cpItcn7vMfy8TwAJeo7
9BNBnRja5PDLX1qP/cl3+sGCSQ82Ol2rzLQPCKUhjaomtHvGURl02lnv3TQ9
TA5vYa8WiyFu/vEF6xBqo8CAZJrtKi93FrDJoSXZJ89UgcFwuuph61ECZXbi
Eh0K5Fce0Nb5WCBHww/06OrETmBwfpwj4AulQNtQuLLKuS/nzKUrDTL2UADd
8GfY2OlvUpSods4lnkYHU08kmRYZYcOt3b06dtIqhoQlamI4I6Sj0YBTahp/
x6l/XBmuE2CtWWqMKtb9sg+yhcSeniISbINN1QjRD2OdOyiVvcbTPhsXGNB4
gHuhtpc4xgvhkz3zrBWCGzLfi+2NVLZlS8Rn6AjsUPKuuB4vWS0vWdGL8s4N
+RwC8t4WjYV3lM2tqsd5s5QdOSAo8py02ovJtENYOE5jjya40nqbml18xiRr
fIIws4t3fkIHFTGYAChOSE1CchAVcmtjGnmWd2nVJH/5xf76DHZy5WcyVcLb
gw/DHqTw8VxeKXYwwl2AXOsDprfuMOjYwILFUAikzfiLWRk4GoamZnxVlLiO
1BjbKwSZ+31UnApFGwYwi+CBGlkL/RF9h60X+A/H6DQdR2bMNWp7WsR0XxIw
YeL3J71dNFFL2Cx81yqRX8bD/In2Lc1P0AmdU1m5IXmUbPDs/PS4qSCVo8rF
1jlA4hQriOprQIxyBxLOVsHH8NYZFm7qDoumuDZgq/tMKhXnHEV0ZokvjbjC
8YFG4N2b2CEqttOC1/Ybd7yeU4iADmAsDjn0Bnzbhyiz/59o9rYm9cn2joRN
/cRPgqruMl7wEeQgdRt2FPlk0mmZOPLBegiklCLifAwc9jy9dLPzp5Z4e2Tx
zEyZ0bmKoQP4hLYwHy1MPk68BjC+bv9NqBjIUbEgIZNiEx1tWX76mw6XHUuD
L6zQWU2NdgMBZZ8Ix3FbsnHYVixfC3EDwdaEByPVjiSwVX4UrCGAhd2ZUa8W
20JddcrwLWs5LUbirptWfWIuk3h15RTofczfRgUXIxa43OhrTRiLSN/mXFw6
2JcsBgefKTNbNU85F1wTZO9QCEYEo5R4p7ivigHmVx5Rz2XvyfouEnhfzmy8
MjLcd9qvLKDV6bUUmoVplClGQWA883MRLIOjcM78gdgeifLeKPcNyxrDYotA
OrhVlDcYnOgUbj3wIr1RRFrlz9UU96r/7MeY3YLAEa93XOvJmn6wTdP32hEd
ZqO3hI/ZHTK31hhc4I8R2Oc74u3a3H3cnusxCmkej7Cn/yxXmMTXvjxtN+vr
/Rkckz4UX8xS6Z0oOsmS3srgy47iGDqFK4LmPVIr7f565ann5wJ+ZfR5FeI/
BRfB5NC/KLmno6o2jwXJxbF3aVzoxbmUuF4MfLuhrspoWPzPQqmVdhFfojg3
JWmFX0e/zOQk5l8RmygqGarV1ytf38ZMgl+RjE96lfIMQ6MPo6Tr+SMolZ7d
21WTM/fV1Dv7R9vJHncrB3SUI7UR4V6oG7Fd6httLf4K2QdH0qQk95j1LeK4
FK6AeuMt+DqGIJ+gRdWuoTeEWPIUfbzAJpOOszmKkax24UDRjYR33D2FGoHf
d4qhz6pxT5cCYSIDEnjlrC5JS6xShbewWa/6t36mYcMI4a7Oeth9TJwaJZaE
mlxfqTxn7V40HCNULhZhBkXMg1bDaIKo7os2CzzyT6dcukZqTKeX3OjMxhFk
8FdE9oDhCjBenahIkFI4cxZd7py/4jlqEcR53TUslWwADLVi6gTeeLZwp/OA
BSGm5noa7uXKSFxz9gOVvsO8s861uxZvIVEALDcjr65D4cek1v+uju36TLvd
UvXolbk6GC1sTLLD42xOtvSGQHYoe1HCk02sksefd6Uuq/GhF/vKbOvV7K1L
Ofn8Vk3u9X6Iz3ZRLrAommSXHuwxbKyE9z2WREkUk5RduzHU4Y9L57WHdQWO
rXfSIG71CCTiNkL875WoYBR/92KFWu4HRFPr9a13m2rztn/oY8DpaWRZ5Rxj
bVJVTWEQUCsBRsX+4nGofFWsQW1kS7K3MlfSQTWdPTvpjAw4yVtwRPdw44LP
jBjkOU72pefGQ9eL9gUqcJ5hrF6ZCmZWMPgNqcOSxwuSqrLkAun95TQhRda7
GuNVtJohad9sjWxMEoReuJ9RucSo4F6/2ZBFTDZgInm+5zcflO/hfp+WmtvI
AnTWWOvxlMyMBVS0jGpsJYblg21IZVm4ddqshaPCYcm2CMvgn7hVgzfYJyDr
g8NHLk0UF9M+aO5cOVoonizZGZAqgMhI8p3+JqxaZZEYUg/Yo5AnpOSoqcNy
S0ZURgikr8KYI++aRvghw57TWPUDgiBgRU2VObOBzsnjG1x7jN6GmDqUlQHn
bfWYjo7HCZYLLslPIyE/ATr9I+5LquVxUc8Mqc0ojAd4Kj8pEvB0k6c+E+BI
jxfJ1/Q3hPo3qUVH2lxnWxQuzge5b21CPVEc4pEGNNhM3or/gG86v3y2ErQv
pdpg9WmeGoPlsghDKsomgeVRDGgV/wl7xnaLe11qfVapx6Yn0f4mmApKylDX
YGwBuwXGYqTsvu0KzOasYabdqKJbof8EXxwV6g6FIP8tIieeNGqp5fvq7Igs
acS9KvX3w9RmrDyqvu0ReHYP8oq+jQKK8rH1VrbxX6bJOJ5ySJlKZ/YbapwB
SteFKo6zRu9l21qYwLCudEkmmh5jo50UrhW8dfiz0qT3cq0TiephD2Dm7Qm/
dHPNO9M5BxzyXDqyxeEL9cCRQYyTzfhfqeDW6TANkFcLQouBCHNYO6UTcavX
Ba7+Tvv6835qP/xqBWrCE/Ff9CAlgDOiAiKGBDqb5eFRxgraG+d1VdfEQVAJ
2BgP0C3paR/t2UJVWzuVSUCSk9IzFGvOeCVRHOHmcu5hzBEEDWCpCbt8FHMl
Pnw0KcXu/fMe/Wo5JeCQfxZtp1n98gicI5kMXx7sa18L3mfWwuLLWA4oct9n
oegWa66/YdGb9OFNucwvMcMnYCShDiKbeWLUlDtMvdHykUQM3mOZiHsZbmsV
9cpDaCQQJbqQt98mUuc0fBkqnbM2PCghKYxi4MlaqcV7LIHIbIUKgaqSE8H6
YbA0GyumcLxm78YzVj5WNH6mOQl9sDeO7aWHGrxDSOVNcWI0xrbhTDOs57hp
jJHyhI+COzbpb5sPY57NMtcDkkxlzGfBJrDsI2GY2k0Ie8QUwTdfNTVF04KZ
cctKcwpyw6sCCn3mtkX32mQmpvRyc3MzpkiViUzuk1nAv9YNBWZCIyWrfcol
RKBB/NXgDAIKRjKc6ERhZnx1PcXZwKP3v/dEzxPvhJHQXaMf7lk1EvAQHiNW
jgMHe5XR6rI3LyfNOLOOqm+kp8EN1UIUWa60Lk2V34DiHvtmdno9k3siKPuz
AntU3pD3oNHVEXVll3xMRjMd79iVSJW/cfGfmJgF0ysrM9yJvytzKabCmgcZ
SEjMSaap8TEug/LBz/gl/ltLeQHK1lI37lHYpf1nRmfH9auFZEuEjAFWRvY+
KIqL8PISCitKAb4pYd4RsUhKe8z/YLN352tiI3N37atztCaKzgH3xkbrm+Rj
Po1dkjXyTsZUVTA3t4SPpBezYACl4lkAt94RafRGNIElOyePr2PflFvaWvnv
UmkUPW36X1E16S12SRALt/Lv1PXVDFvp79akQ1ORjV4IMZkF0vk0MfSq1j6v
bajBJr4KSACXctqVyZP0wnhRxzqzV9L7GDgi5n6te1XSp49NL8wWcxqPM9Oy
lsd2fDXIcoDA/nUfobCHRz3MWWF5dd3wFayquc8tnI3beReJY1TW5h95WcAy
uTYtn+auxWEL3YxYCrT0gG1Ja/uWgjwMpzEG+dlOF1bQ0GikxPJpNlhS+5Pq
LgL+siSDaLlAZ7o0xhy9qLVCX2lCXlRw6aoesnUQzoBOvcxecNC4FB4w469U
wAAvp276M9h2gUOLTovbWX0RJ+goPY/VYu3sKEfgKPbcaUCsqhbPYesrGtR3
MB7EibkFuF0pt2ZzQPR3mJzBA0IjKCwzMwQdfTUdhcwVoFc9V0ZJqWpLN8NB
JWHtyw62e5UZXshXRmx34DjLgPL4pTjyIs3WsXt3DHtHXEFerxYKDFYgUmm9
kPOBwFq7UiIPSDcBs8b1vxWIx0PxMSp5sbrBWDvBsI+MGOJuUWgCrgwUhrLI
4QCgBt1VPdpnbcPz38g0ySklE3vo2dQQYn3IhJCQKr5h3PEmFv7ar4R13pZV
NSDldJ/Zl1AZPdQwEgf6bSc+W7GH18CI1f4vcPZWzDgIEihYS6j1+5XnN8aw
89Ncwl9fvpbZhnt5EqJSIJnANtrUoUg1osVtAVyH/QkQJli0PeNvXUHwcvt/
h1hJnFkbd1bi28k/SR6qPID4FJYTKU+IF76Ev+lSsNmz0RSDG4alDNqOzNg+
GSWFu0R7ulGgOYYGnk3la55o7ZR+lFqugG6M5dWbVrnt+rRrr8XY28rLY9ih
c3TFOZoD3wKOyH4HjrUIzmWpObu5ZzjNRjBkjirGShnrrmst8OwBJBJf0mrc
4F37EWSVt3YUUxOOnDoXSPVu6n3udY9hg2o3jS3NgHsTNp55VVEYaXAnW81K
kVWuaIgu/yuC8iSaa6MYTLR5qXr6yTmPbDSRf9caojG32gdmOeOWtWltILa6
4G4dqkhk0gGCSbppqK8bttMHwC6nEPP+0HhNUyTOD/lfX/Csd4peKHyHbOkP
wPzjVrf7y3upz4r/ae99GBNkFsA/pAB7p5ivriPga6YDkeUmH8eRBORbCTk4
WaOeO/z2SyrgltlHcKB8HWvRQfg1sTIIevBWDssfqYVcxSnqOVcAu0F3S/7F
y3CAtdHSUQUOjb/q3saY0we9DSmxXLi3+EzDwFVDBgZONvk6TIaTFM+mMkKi
+oHzKx01MYp5A7IgiY2gqqBv796BM0vtzBhT5jO0E/RwxIruMwno0XB2YKIn
pnKO0Hi9wQmnCUYg2egjtu1qECaiZ/y9vOh4lWBOyIDPeCZPid2coNXfSZyf
1NjcRJCcOYxfH1Q+Zg5gQEjbGei/TSvAMQ/8ckmIPfzxzXJXo/DI16FERWIS
iifAvoXqD57tZZGaG2aTI+4w2FgKh9FpOwSUDeqYKfDsfrT+2Pif7eJylPYU
pCsNjj6bl3sYVcdrUIA8L0gEAiPbzy/O/Nva8QimSExMMTa2ekZmZdZSrb5+
j8q8IPspmOrOYXNtRqOrj6Yvq/nYhM9kARMZrXSHA33B25W2TSYTjnUZKF2d
n4dteLzWMGZm5W8gqcDHMRvul6xF8gcDaOniGE6nwL0vGgJ/DzOzQV3biXWY
8cyyk9ZnTEnMUGfRrHIEbLHZDGTL7HWzwyrlfDy++MJXuWQ3YHUCHQCZaFTX
tWiBRQDn4X1qUOOMw5f1onFTkjGuad9U0wZTWFhwLZgNHCyhUmLCx6QfT/tb
aImkAoDq0j8MatlcfQk8kDw8ONp5YkEepAQ0SolQJcmkhFoKfQsaHBUVbzst
oorxifDGL2EnJbqmsTQU8YdxcmmXstbVqNx0OR3eDT3GxrGRiRS0abfTFrNX
O58dRcMIts+L+W4/XGAcwFIooyNllPYllaKdimnG3pQ5GjB/IWBiSOwdk27N
ACfb3RSzrFwAvtKgwPt25gw2a+BrKmRS5Snf4O8yEyU5RlqdrRKFoyeLuvvb
mgTEbmCc5dAzMNnA0hrMgFh1XlniPVKjxraOFmJ2kw3mZSnY0ME2oOWgPiet
/h1BJERxeKPvBroFHKBlYqF5SeCYLDyzdmhVDBxZuAURXo5W+Y8H5p4JHNUs
qwjo6wkzsuVkwf4fII11E4L9v+caPZu6QskzWZ/ADGDSIQvilE4MFhRPNf0O
x2/ODZsAKlhcPiXL54EpbiqRw0AxNLqJXtTRPEOnNwvAxuLtoD+TEMqqJQxT
k2wreh/ntXq92vxTWusTkVBFNavViwB7849cprDYhOyqynYeSN+w3LCKE904
1PG79Lar2Ae7/YCUKFYvGhbQv2w2oLMGoa26VkLh3sEEOgKCFBC/TqDOcC92
4YZhaz8lFb9ep6tOIL5xjSPdHGuPwrE1AnZeJT5BYFSgOLUWAtkciHzD659r
cHYPNyPGgDmeJCXN4NnvK9qK4R5D0qS8CHlwZffEQveJXyJW6LfMGrMeLIFX
KfSTWsHWCfmgOZEdRIF08czAb4oW7AK3brSx7geaAyX47xMjxu0TR7kCeFyX
pSr1+LN7M2qjQPhrDP4HK2rK4rOpeZod6WM+UoTFIKFuiFkU6F4E8HWM1MLy
QUdQN+zJIUGNU1o6rs5V9B6CzRO52iXGvAh5FHQ5nHpE5kIrwV84a2pO2IGv
GC1BKcK+FGNhqRVoTiHpKP2vy/pF/HCyc/I6eR3i2fj8PjLvLKkpUCnTHKJP
pvrDp6uidp4BUA/3df6bthKmH/Xq3Fsdazw+Yv0FVoy5yf1EZpv97tWUupBl
0HaxVS6NGU9YvTyionVsHiFaogti7/+7rnNAbAzMWu0G/ccri7MZ0Qc38+cx
rQT3LbSDATaJu+yKj4gcbLiRr2zIadeJa0/YxTWv/NbbcC/z/RRdWyoqdfu7
cAc+Z7SMAwlHZRlNgLJZtm8fKbbjgSoBITS5LTNPSCQR6sl6meWv02aLtz1S
KtGuY/U0wqTnNRcj8dHlCy7Ph8zjopHMVIobPww2YYk/Ak0tUg6baJ5p1TBA
0AiG4YKkAOBJcYWq5kPoYXNE4paexwf6cTQiZFUhw0nWxMBKGL78cAknNSHl
mOxIxsrMe+GIfXMRgS1oOBoXvfHZfoLXDXLbwWBwP6PzZZpbSLhQ/lI2+2yE
3t4jXIhpn8hJ7T0fz1S2z2c9RrNOLqKzL/Rg7R/bNdAR3fKQk0ro3dtqvEZP
tHepxrU6luu5DfAytMR7+NytOyHrTvMXjrlvZzsIBk568YfApYTtztcCJNtp
PD9u5h5mQJNx0YyE6IPoWDYmWT6/kMT4qJeJmYH/6pqRmHS+bvnwoJlzWdme
hAUcYJhD4rsd6qx8Uja+btA0G9H5jyxYCnno79eAeTjIfuhF8Arze1mdrsh2
XbX5Ck7qOzY3kqhMA/zu2j2DA0mvh6NVnQ96+wkCvKCrfI5dsHatb/nxJZya
nuaTRMymLQSM+xswZgUkt6ox/80xgurxHCOv6/mi5LOjXGv2/mMzsa8FPENH
FH3+MSbqE/gjyE5N3C7sgi65GVX1aVLQlPSRYcGvbOAmYzq2DPT6kg6Anfkf
yo0guei3xco8jKyHZXeY8QpIdW2LCD8pvBua9FslmSpRbgGZILoFhaLui336
v/xmsnnXGNvmBv+I4RDLZLrOJNhBZqiyuTS37Z2zUENYNmCJFNCfLwrDJbuW
e9yvDkSY6vh4Rh9upmYYATlFrM7B5535LIY1CjNQ6FY9e1Ae6PpYTq/WHd7N
RuEa2PsZVjNmMslWTHU/NFbW47TIrrP5sdlDyUlMkUMNdCrEDYZ3KH4hXEz0
Ru3WVKXZm+RdjNEQ+4WVPOlkkisvZ9x05TbZ02GuMep/Aa4g6pYK7WjkTctp
pn+IeKGY5hTlIoK7lIXN6eYY27e+zhZpSUUQqEsOQHcI/L3ZGjBL5zdh2A4b
z0kF6tU4AH8HqvPmOpLlhG85BkRd9BHC4tin2qtR7fTeJ6u7PHcqNC2uk00v
CRosP5dyB05YBwPoXJDBzBxtT3I2eyVUp3yLilu6gnahlhd3ACnk3EAMgVW6
ZS9FXOjhm68/++xB+sjOQORlJ/fvS5cNSoSfB0fWtq4DiIUTBn6syZPC9EaB
5PwAfWh+N3ksYw7mzozpPiBThO4KYxXDgfz1p92nc4354bC47sv4DtRy/rgP
59ZxZT3a2awp9B/dbbl2MPtBJYUgwJq0J4S5vk0+l3k4F9Xaj9YcmLtjbTP6
rqUdNsJTshi6PT+9QZfXBVE5k6zT/GzbRusPqz2qSunq3elFZaTStqq8Vv5k
J3p4hRoRjPTLJjoHDjTGiA5JBpo286YXPPiFr7aaINufuH956AheYa0VUAxS
d4IAYmeSljS7ldBTmCRGOgNxH4HcbDp212W0u8nr8ZL7rgTxWWKWg9YVXNgw
YbmswxeIOm+x2jbTwMSL0pyKz6jJzrWh0/6arFVyOmZe5f7wm7vJ1rV3JJI8
LeJVJFVBu351YnQwE04A4GXZl8XF9T4p7uLM60KedQCTNsGumsn0V2pyhewa
KHI/QdFIPzMXjJKpp/NcmgSIEQE6mvjBrmaynAKjwjdG3FIdaRYf9rbE4L2H
3UlcLNy+72e/xhouw273fSVvBuajxo99gTK3spdm6auxr0zom31MUF6JECf4
RHuhKNUmZyLdJd1miVfsTZpJ3yJ0mazzkMfLtqagebxS37gug0pRaRGgmp+1
q3ObR/3CPMn14tL8VuXPd/8RD4Z5wf1lsAC9R6W9R9P4PS1AtdSvWQtu2yc9
KnbBUBCjYKuNb/CXG1hOLebGApAnKe90gY/kGg2AmZcVJdkNaD8TmJanoyEF
GfzKRV9zLZz9zyuN31F04MP8/D/Q9Ag4GSTTsG8GFAwvSSNKTd64Mb1K0VrK
j4bpy62jXX0ew8p8bJe0BujYDR8KCXjgLYiSiWLoZDRH3UUZsv5IcJx7OIMl
/P+IS3MJ89yXaXx0RX50EegtArS2913pr/ncvt5wj4zxsblA1xs/Sr8HoY/x
EDDhpM3SagfqQyOmzYC9T45KG9wc21idgSTMyzYR435uertYiwos+MZ2elVm
yjEYdImwxwnaOj+B5injUVr6M7TnfXbB2GHqUZmU8kAeisuCm8a6Bt9I6o+j
wJup/DLQAheoLx2l4lsCDLX0PRVc2PV4vlyxtI/p2MMdyTopwfICxaAPg2MC
PNGvopQx02AwAWFDJIH2od37UkFoRfcFZvEVQ2n7BLL4cF9r7cG9pPFop1Ie
rDQZiJwfJLA/z+dpTfayRo6wAhoGEjgsUWSyOOPfNv9VBrbJP3x2Gslg3yot
7d0JMIjFKsiSEvD6PejnX6k08F4u+FikKtEi+8dUebUx2PXJgWDjXD7W8wg8
ch78tDhpfamHjwrqV7anVQAOdPDvUD8C/uZsNyqzI6zh6s3wXmtRxk9wz2F7
UVx9/10Doo6eaCEnF7TEBBvclOP1QAvD49PU/lJpaq/nHz0Qmqv3J178gRDF
nQiRB+NDnrgI8L+kAav+gHJBD1Dp4GOtRhHG4DCFHuJrCLiu8NTUBT9Aq5IN
l9gsm/jKYvNdni0duYA6fXulb1ZDSF9IYvYogmREUYk/XHMKCz7fbI82QtR4
iRZp4ExxcbasiLSVJ4Qwh7L+JIHDuoepkejYeXfAkpBauEEpuSRFlmAoG2SM
3t/38TK3OXWbVCZyII2DCNZvdYAjXt9CYOFc1uiullaVFJRTyxESvr0P/9XZ
OdsKUhj6A2jU/wV3b8Vr8thDl5NsYPEa2wM2caYapoGalkYn/s0vJx4GvtdE
lqJp987WFAZl6eixs1INOmXZSKuEE45K4Jp3dqng2QHCGVEfXq8LJ8yDcc2x
7nVhjqlmXSBvTIYzaJRFPWJj4lMGyC+OXoEncA8P5VjBhs4mz0XiurZntnab
apSbJUfiROzFKoM/oqqV5z5zaVdVaUCYqyTriCQrprr+if6JsNO+hXtgk7yS
xU3GAHQYw3taWqGzFgmRtqJmna05QGKqGWDXkErHUtXgyH9LX9XiSqdiqM+d
yX1nXy70pH+dA0ChU/uE0Q5uzT14dv0Iph5E1GQKxwSTMn2adRgJkq+Mxggd
SSrC7KDL6LYyn8vyC6t+Ctk+/zG2jfuIx4BTofZRGuyhiHxBFz1IlDJ/5ppA
tGlTK4fs7mq3dIq6r4EMPFF4wC0o59p868JRo8tYPEuV+PWq2Be4D6O0YT+G
cjbQxN8bs0MMDO+xIvIL9BKW6XQCL6ScgYmFRPUFUOCs0I0KT3y6dgM/yxya
QiWcdSW6RrJgsNGvj4XVRmbYFGqJHM5xaP5YPihhS9g/dQ0gGRwFKrSRzhTo
Ud64P0PzIgYOAhYEAvq19R8cFzklLSb4tztl6ctJejmvrUHcvBItNN7bN4Vu
Sm5dGNkotq12fb01hUpPNYxAukLH4CBUXElFuf9cHg3+zaUXgfm75vqJYryW
XskPLAk48S1nSBThgRLUNYdATg8cuol87sYbsYY27K1ZBSkh0080V8m4ECl9
cYKOV/w1YcKJYyPBsoAtxH2Eyy3S2xzciP/gLazIiLAdVpa2M9IURofj32oG
GECX+lm/srTMPefIhxXEDcYQQUEiNvKBrdgR4nB4HHzL6ZhJApA2taEpXEsB
fNpID/4AsiBlYsGkkHYHWLQxeX9z9bQxkOAlH5uBBzlZblyLYSCND12uZTDX
Onvy8Y10iCiJe/eNwlUEMU5jZRezHMHguGYrRnkvUSQN2OAwvisutYhmPlOE
fgpJNNp0G88yvNYSrplQMwwrF8CUC41rSRB1gpA+54Wm64ojB8QEcdmJJzYi
2uPfa5Wo0MylrGaivsYB5KXYlgpldkeaQCLaRmHtWKXKmu/rUXc6JAAGWCvG
ughWwIyRocDlATkltecJI/MSbzn8HXHJ1FzFoHVZ5bXbLLOiwnoxd8s2JkUQ
ZpucXAJKFdtZr2wd8Y2rHOlfd90spfCUy/IRiNIH/L3XFRCYzchLq3aPpWhC
NBf52Rw+oBIstbiuh5Y4Fav8yoUy/1DuVCWzZMTVScBhoT9eBKB1MDo0SMRE
V0hsZ9gAre4Sj/fuM/PncuERLicdmT7DV9LqudRO/FTWNpM/UMv1CO9/y3ip
IY7FtK3kK65Zoi2d3mBAk75WTd+2a+H7F01TCJmb2qq4D0fjEp4jap7OOPTg
Pagl8GwcETuaU0T97P72C6K8FVXhbbZmDPrFbDOsLEZ0NLysqbUjOKKwIKZb
hCNXXeQCnEoChMRQgP7TlQ3jVvDIK7/TPkIJYbbK/AFQxB1QLUCzOWffM3h1
tsLQ4a9Ra8gwhhq+k050nCqi/6Fw0gE2+m3Na7b4RERAjrijpa9CvcqXQhDj
RJExpsnac8NlwxAuSEN9FVnkZ4/wS3gVHy7WAeXYGm9mDX5lZhy5E3eQawNQ
XDYAshmEHsNX2bEDR2ROxXyFJROPKVueAKyOFZ2DrxOdPuTLVBog7n5TacJc
XeLtG3+xhUfC1mEpj6C57/9Gll4DZPhCL9I/i8wR8BAoYqibxkSXtUri9TcP
ERMuPPq4To2i+FZ69LeqPKnw+0DJpHHX4bIahWtaNQsBUMDJsTYdy2ZUBeCf
TGXWKDrAOBnuaJgl7x/eUs7beB5ZDi04brJYVUGv9qUuG3L4F4PSHqyZKTLo
nZ29Kx8sxqQYRDueuuRFFdkC61uwdTtXZ+RYpH4oXuOkVbh5jNh4SV9+gU/C
mcUxkooCeQ0lI7+1ybzjj1dAtYklSwZGx6AEC/BtJn1c89QMvJ/0/Vvunsmm
DzaJ2Jzh6imBbSlMnreVW5XgyjpM0VzNcrNC5FTysCR6K+oV/cQGLrrkLs5a
12aYIO0p/BtNe8cfSgWtkEAQW4TIfwcp2t4YsW+0Ro4+xGi0ZvWxcVEuTIwJ
//gSq/cNOz/Vus/QzgEU1+0fU686Ppr+suNCCld/kKGfJEmL2V6/KxXfBL5w
PJKUvAnAzrmAKdLsIsQ3+8t1IkyCC5pnwWDv3+oEOYIuZNyZlgLWHYRDXq+L
wsmoYlwMjG8oV9wQYSb9iKNUrMDablSvHZBHl9uc3gMXf4lmW5wXFVIJf55o
P4bEYNGvkbOAkm27hAlvumvh84zHk9ixRDEuESdGqHF1LjclgVjc4PQhtL0j
e6HqP80JfBnM73oB3sPk5VlvJ9s6F9HV7rPUdV1oFJLnQDQWn+dtxNxbhIPS
L2CGehNn51+Ji4GlCm7H9bM1hWzOJCHxWkifJPtO3IBfF/w5noF7SS1wlxvz
sp2iEk8ESwZ4R75UIaxj4DF6Dr3FCcomJfFGpt9oCVcYIs3WiQ/S5bHjGe0P
8kifCCQ4icq593c+f1Swv6rmni2W24NUUpPjVPRoHF3izYn8yPvbtj3h1UzS
OYNJG1XWjWdPS8ggZGeB6dtwJI+3IE9dvjexI5ns6X+VHN59VZuaNTHkLBer
3dS929BUEZx+iA3sSTPsryBgQR3aeS2e7I609yTeRnndliKkic41j1eHD4Cg
ufvFgf/EkrIFLYkZTbwgq7oFJnUZ8/bPCWTXAnBu7GBd9ndh+JfrjXSyflqt
qi58WKGLuKX3XhciQfwB6qqmVw7EWRAsrbn4ot6XoNbiqbWIiVj3aNRvxi06
TycJJ+HXiT1M46yVAyWddYjcqmTwszD8vkJpyM5HVmvCbued10Ar37iMbiQ5
uOYO7n1nctFZMLdUygge4tUVuRMDdt3O1YwS1GW2rlpdHN+MvWnh8OGFJQdg
ae3lmuDcoqmgN9aBcPxSbi7o6MSDyBbuJJ569Og4a5A/Q0/zqfyhl0zB9N+B
gST4E4CyqyqAWU4s0EX2snBikqT6fN3sEHZgy3VwSAHTuy7cRcS9VAjOrii0
917w//LN9IYupNQ9T6gbjY+IxZwXjVPlDfpHdL5w6uStVua2VlEfCp/YKU24
dJ7LSOZK1f1g1ivOtl9gCPM2be7xzs9dw77R1v/BmXep5zK+mnIO4iVV48yP
KLe5djnMPg8yhBHnwreziLsd4no3yGGIgEh2/1SJJGh3VbnIt36tQAvjnwpL
jHX+ePLRW06j+6PL0sfa7BUzozw+9pidJB45Qpg3eajTnfRXY3PBb9oYJsVY
FYF4ktTOncUseyCOi2UGitfs+Keyq4KewM84s0oDopSKxa9zEWOyaCadR2hi
aJsQ3doQpCMxBujSxBj491cZ0STAr/c/kJjRyvFnEn3pUPqNN/n4kRuQa0Si
MTADNG47lxkbeXNTdyVAy1DmFhxTybTlx9kujT1avRmAwz1pKM8JgFPmnI+2
AtFYHZwprTjrT1WtodTDrjI9x6ElAPIqjr0899l6erfozkAs+P23JG9LRuHh
9aFzyt45uhEqp54JMPIp2ktlPh8nESTL78E9eW5KFVtU7TgJoUJFEbrrquHX
vX5hgJVciokZ4tfwAW5/osnX5VJUN1sprU+bpc4tRWBLEuz19sSCkTy+8qYe
rgJpz/BmXUMkzpk+xCG8Tl7QhYIucAfobvWZ0aX4ia7A1o0xS5gtm57rJQVo
hcqOE54e9+/qWGBP7VgYm2rDZf4M2JkmShRaAhQnhBqcjbFZ7VMJ2B+6dQVd
M8IrWVBaxaWZjqWcOkQUlF3vfvS8fBg63oJvRLjCS+A3P1LZMV0vf/Q8YnyW
CHgdYefcJopIAo3VtMB25zniw9g55a2/CL5UytjVRKgH8PjrFFgG7/TKNRjF
NeDHz/frWLlm23PKojUfxjzBFl1EXwbsU0LYMVIz1gHUPodZpzqOPT1PDB/k
SwrmERgXANy5fD7pZOMebd/aNHcorRiAd083Whp30xCtmY7W78h9A1uv/mSV
qZ7XSULFDE1Bl5cvG8V089opPrUYGo7KqWvd+leHO9b9O3h7M+Jb3FIztfgb
TAn5XNPrgqe5C1O/cp54sEKRr3L2AtBqKZFkeOSGedxem8c92RcY6OdgVxlO
cnqqK//txl75EZukzynAotyYhYWw7AYtaG9hnms1Y3Z29zMDgaTKDTuqb3sf
HKlqbobxrZyR7jZz+ChM2yhh1GGmyHdJaSGklbpmycQmAKYHmPXqbm07Kwxg
vuK71ZNBEp/YPZ8kH58Whl6vXBeY/yWl8l4AEAmB9KK5YQHoVMdgP0SuN7C4
kuzHXe5P8eksixT8jFuYTPjiLHpZ7zSSGqykGso0/xASDx85CJkgznpX4pm4
/Yu+fViYqDQK0sJ4MRamQ1tNLx6/VeDavVazcXEPSTkYxF6xztAKXrtozUPO
soqOUN76MOA0ToZm3GM93gTvtAC83G9Gy2sUxIypa6gQnfUsc7HsN4y3Qo7e
N3kVBhJzq13Gd6axG9sX7+w2Y5A+Vy1nJvfs85jzmXHQrYwngAVF3qrzA6Gb
Hdt4bIqKluUs7g3rWfF5qplr/v+Xw4ZeBQ4dv+Xcq/013iDWo7aeLQo0Bcy4
mfx5tOu9Sv/OSWG+KmKQrgUjtXFfhV1n+l79GUyMoMSPqQ+UsKb5mkhiXe18
3s2dj8ur+9eWPQmsspGUPUeSON96hQ4Y0VvHwtyfD0lVeZWBDyi7ZMwqKMyL
mxZGWoxGpR3mqcpCfNKf6NHUI8jcPfqHiZiwmEkDHWVpA+pLdV5QTd2ssZLW
1V2iFhk59wfyw2A0wfrPEuI6afNvJh5U3EPrI2XB/kRWG9Y+oi8UpuS13u+7
mUP5BsSMAYrb2IrY6p+djLVFmdZIEWAr9jf9BTYZGfJ1aHhygbMejPks+QM0
TfwnqVy+6ov8KqyUyUvPqz/8JI/gTAK+rDT4Em1/3dFePetlCnSKTjj5XXBx
pkU1NZc9/hThoeqZQq1Oz73jH5MOPGu/HfC/UuL4tmIqENjKC4stg8olgJjb
ju6ES6UN5Iqu+hAVgQnQ3HwfMBea1aYgJW46IGLU+Tb84O/HecrVsa51axzF
S65MBfV4u4BqwSG999XCP7qDJoFlMo/lpJdlv02BIp4rizyh9zvC2oT7eOCV
49y/I4A4GF4I7cPGSj9jyDRsRTLT8hhz51JC18Ij1iAQfqU378C9zGrDEr2L
117rDYgB/dE436ObZlnXKQ+qV0LwA8GBkVkI7lnXhhvX8uSEv+WfasQfXztP
ciD9QLXHkAxNTzjJfsPhpeHCSU0SdAoLhliugy4cjNgVGmY9Ztv6Oes98Ya3
Excojcyxugc4CfhCCLsVCPdc9LxWumxFTx1GD7Ju4gv3za+oIMVGTF8u8HNb
bKqfd02VNm6/MwnrrCjqf1h2QsdnztRFaz0RnzjgcyNSNStUpQE78hFmXfbg
VKsFsH+N24A7FjtzptebcXs3PUFJ+Yre1jTVqwdCfn+d1Bk/zWux1FiZSbxZ
BuAFuoadZ2chYNZmFjtfKsUoZlOAbRoI66k6iiezFLcmqLrczK4vAGqQCIxu
OFlUjJ4p0vfGMMtncP8JTmUFcOyTOiZ3DEls7jBV6a1XNYRDqI2/rXM0piUf
FNGI9kW5UDGlUIYqhetzuJuY0m1tRKlGiYsBzRJ56uR0YvUfUwUKMzV4LzA1
GNR524/hJEykIjo2KmYFcz2Lg8UbMZzbcEwML8AmHf8poEn0llChHJiNEhXT
+6kBgLyio0v/hDtXnIgZeqp7ORCwcCeO39W/kxSmG54nMFdxBGDgIiNRiMFa
8cLgfJTjOA3g2yn/09xTIbdXhQ77tUlXVwz4/lvqgiSgN8zBkfReaVdHKcbk
2SLTnVpdEogxDDvkCcvPWKD8yIBRKjHA1Ez5+4GTSmv887tP6t7N+i3RvXLY
imydZ/K1wsqcwG/LajnBT0cBDM2BiEsrr0HxqJVl6OhXQZLaE8fVjLIzF9GE
cCf5o2jAXNV3lOW/5lbU1iRwwXUIi3CZXJjTEw6xS8QZxQNZz1LHAdeSuS48
w2a6zIYwtQrXJFU6El/LfdeibXDYtDpnDqSIV6UbLIih7YoCXoCR7XUbzq0E
Czs7pyU5q2A4CDEdZBsVrxXEZg42LjQgcvSO1AeD9ApPAstczjB611nSjvM7
VHwiA0mz7r4LNkTpGlsQck0rJsmryVcVSbyn/MRpVBsx2tH09sN3Zi+Ec3ak
VN9uvMOPfMHF9okyLVf/s6AmQrVbu5ODxtxRV15xmQVCH8F1y4q3Nze+WL2E
fl+yPpXaN+l+Kg6B6l8PeYpZJquAIVzji8g+WehegcG76ek3c/s7U6GzekGM
L8aG31C5PftlWOV1pbZTYeqoooclXM/SmdLDhgBnYesr8GEnetQjuktubS6P
XY1pXolH6/5xWB0e/yT40VSAK3OhA78vq9OxzpGofEcGtMvZtVX3I2l8lrsY
nXJY8Fu4AUxHh2dyyL6ew3Z8HfpZUaY3zpp/y2PDqxOe8bussX3bTaU4UfCI
lmO+htxuLIzm6G5pwenz0NIV9XMGulov6OpuZqglS+9fq4wNQcNKCMv+XDYz
tv0aJvte12SkYDDYKqj2WQtButefRPuR5cUmiPpbgTaJvvfwmFNeIFREMz3T
S9Hnquvbund2uITExSE7X2y2SLIeTqKqdc51mcNDoSgusfCCOj91cl3/lshq
Sff2OrM8ASbMg0YAs6z/McMOr5wPivblHaDy5HNqUzpFOinijWwAwYeLu8bz
W882yxxwSAnKbqudaiJJbWrHvUiiKiwiyvY2Ovr7VEydlrCitF7fA+LKkCjM
ZRm2shRzUIQmQvwaRYMLWfFBtYl8wjCWa2tMLuHDR3CXOeuYfJABH/zEbBfD
skdE1xRJD8iQnk43tBB6n849/P57WCecS6qM68Gr44DQ8aW7u6ZzsrCWdNK9
TC8EPzuhUAHJIGfp1wKU5732LeINUT2dT6xK+4GKnoUBLCyVc+tkiCHIGW5M
kc7YkW3a17S4D3RzEacZYDM4czc8FEbDA48csq/OT5iiVF1XX8WTyNiwWNT1
q4sj2mj2PS+s0pNxNRgNfAFVG4t/8LQ/B0q86I0uit1A1kWawCTTu0ftkcyt
nKIxSd6WSy4tpTS/uAiv+ymNueezXh+qtmIGgqsTqo8Pm5ICLSckr4J/P1rw
KjDpr99nj9LPseX0PFY+2/WijvZt0LHNM/o9axwMCNwqO9++jT9EpCHeub8o
CUNKuyxppP28ICN9xDOkauFNWtjsLmHRckDMBpQPX6CRc/wFWroWCw11iuIi
ynznKekAUdIWHpc5zOf74k0oK2SpWTB5nScQnI5+Nm3MR1zQC1FrG4YUcQnq
Tn7Z05BlYdL7YYxC158QDBVaqnJuSlgwmx13021bU4e1zMQ1siWrdXDUAAj9
EuhUvSE3uyYi6Pl4pf/6isIn15tVjf8fVAJS4d1DUtUtwA6FCD+sHldI7PLb
mmgDMyN77mHGFw8tSemoxNadwT4IX66pRsDqXzx50ALmNfQ9J0O2L5JN1O5z
zZLxRyEJ2np8jkf46QuShVG7EoGAoq8BiS1pYX4MfCcsovfCXdHtL2i+7jU9
BemWM9BYQCExC4XMenX8NemNB7zkrpYVsMOg5lsMBusy1QJeGQezWEyqT+pO
51z+kxce+wvv8vqgYevQD/VmVAOxrckaN3dAG7FaN6jjI6Cl+e/ktvmtfvpE
g96xJIOeGoBnHJePFBpHK6LMyQncn5Fwy1svUBf2WVwv5GFGLReqnR18sZTC
BPnsktTIOK87gd4l0K3E3JiS+sWO8nSVFEjxBUspwIfoR8AMllAtRD6rMgl9
Ntb6WekBSQ88yYcM5uzAEXjF+o3SDU12Pi+mAMPePFJD0K3O0STOk0jd8Ad5
/tca15NdItgtjU44Gi08Tuun5zZzNbXGH7Q5ES0jsqSIlOUnRgPQDCYGxaHr
iyEDYjXAQ3iFTP04iVUDHpNb2vHFnNA9ZzOt+nRQEunR1fHzks3xyfhDblGo
+lQ7WT6MhjUbwE0iQdW7SHEBO7+4UsLxnZy86minC/CF03KKlt2MFRJTVOd5
0MyWH1m1Myx3f9fXdNwrK3ANRQpX+r3mNNfTMONzcNH/l5F6/O3sFhbOJDcj
BhZk8HzmROAHhCo8VQDlJRyPD5PuIVjSaVdlM/B11KQjWj+8VdSq0aHuDAbZ
ll/qi1JXau1wDffQpSnzSkT3nZM86sudmQi1gQWmyVECMF5QLVfkUvZgkeRX
rk1Y5YmtznbnVN7Zur9YxZMgXpUzatpY/UGsUVBDrf/8sh8VFFjQXZ4aKZ4b
vL2XxPIfJ+kREsT9iJlRYsHzNhCKFPPngJYyeiEdlhOseOxWsElancp9mPLX
XuzVxVBEez/8u65ST+v2yfVXMprzAYObitgF22vb2wXwYalM6t+LS3wG4/ZX
mUa7CRXi1BRgbgi1hLW1HQT0eO+M66febXITUmPZy8jkxxxz3Q4B/hYhEMJm
FJTNX5qAqViLsSKANc+9iJ4Tg/PSwgT6qGhdkS9FL0wi9yUWBAXd6XhuRqNT
n5dqnsLgYiqyppvNazIbjmE+4Fiu2PxfHysB1aKCM3F+y0KuzNqaf4lEvjVU
OWxYdxtlrX218wN792aj3BZmBBxBQZSivyuQuVpFUAKn2OaR2zLeqoGUX1hw
zRKkq///xEjgy9rK3CN700x6gaHRgNQ+81u0CRm7sM0u1qF/JvjZD98j3mXX
HilTI6bHfKMAFxA0jU47vOQsLfrN4eY0E9jubCrrDoflELEhuOs3ZlNDyIKp
wQ3vTBZqbIKcUTLoXmZhydga0yssXU2/W1G6d9PGjfzYRAzNTatFTru1kF2J
vx59vfmF1TnIAy7EjG8y7cYfJ4glNdkmCSGXrSERecuAWFJM+h6HuWGh4aHg
bEHBlCvjRYhNCSwl5J/gRkHpU/QusfMaikCeg14z9atEIURLFOyEhinaqlVS
xDGzZXf7qRImAVHzsaC45tJnOv7gxdpf3+9mkCLaSDp9JDGGEbk1LZUNYYi2
zrskRT6sEQFyyMiEjmbmriKVAFFkOa7fmU/gELGK6sGiGEbaUTzvTZMLwGvo
QNsvIbVqEwCoIQlZG8byi7yqGPY1IrB+eCQW49Fb6loXv0dMz/RZHoL4MtSl
9Ewe9D5A3kQeOSzeEppJywhv5QdHcrO7T3wclGSGt/juF7KfCV7VPJ4Irtaq
UCvUI5MuCjqFlonCRwU9zIfViDxMZY9mZZDtnV/HHwJoiD3k98P9B9acRV8h
dU08lx//HaUEAOy4GYpBK17GmAo/3YEfkUmbFhcFVy+i6/jV55vzifhe8r3X
Wc2zCj87pvCJK9cQp/yraobWgGUNMBaeBYutkIcQZl7bhyIQ1KAIVR+HPaz6
iCcJwYJ+ODGt4O/u6so36n8PiZhsMxRSqW5OYhWuIbL9dqnV5DhfrrjOyVwk
5lqN2wnOYfgeueH0VD4kGpMTL76/0xjMSmzcAo8+4n+Ks/m79uGaAquK+e1k
V4a4ZRzqO6Len7eHHOBFNdx3gZkHii1UiVuy62Lkig5Y4uYNChPtHi03KUAe
kuit4s/giesEKvjQbxhhZ+boYcLb0jvsHEUQiUw2OOqeK432e836dTQrWlgu
LW/Tcc1OtZvZe8eJkOQd1m1FRtTiUMpi+ksrcyw9Guxk6fkqLEsn17txHgXg
Dr9nMXZHv5o2o9MYIM3eSbp6NdnENdNkeeNInYEPD6PQu3XEZq0TCr7b0zN2
/rsrJhusUS9Jgd5d/BuqZ/oCxBQgv2R6Duvm0b2BE1cHDGF/XT06TWKGcrs0
mebGxMc6XwY5awFy0Xl7W9gxCrZWjRZWmgp4/Kok50Ndi5UHFSyWEssxeNk1
mQLqJvKasdebrZmhy/APQDjKN69wN7PvJQ4u9HiW9QKSmkofZDiA0ztrda1V
j7rurcts10Kh1rKaf+h5Pm/JyscHNnjDK9/j2UkNA1Uj9S2idSyPNPYa4yuV
Equby1XeIIGtAk1zgq4mPfYV2PFEHQmrx8oRjHqIckoikCjRNFOQCMcXE1UE
p+KC4KIRu4sKdqqBLFp3RQHVgU24yM7uTD83KSje/ZmW+EuSjNV6wVedhGVS
NXqzbjlcsKy0I8yzanS/pS82Ty3QD865vnI2SBGDfnDTJfqpwNhnOx19Tu2h
y4s5MB86el+8JO8Ye1YjBVJY9ggQm3POLc5Brca0/ERoDEq1DdFS/bXAwn+z
u5OeBx3YJCjBX6iDUzRpvuwaKOAckT8JbZWLzh0lNID/Zw8uA91cbMIyQgg4
ZUPfOpzBvlk5wR9LiVNDjOIc0oletiHKqbLKoP7DDYsK6BDNBWKBsASLQIrF
IGXh5pLIkzp3cNn6JslF9a10cNnhYsoUc6TkFM65fhlZ9ROqiEdQModl061t
VNikYKiL9A8lj3Gz5+r9mnngEK55XRX3T0mUZnKIXD4jBNbWARUmjMeVS9tf
Z/VKVZropZ+hVadz6m6Nrxry54fQ7x1/+KMoo2wC+eQT1BLC75Gs4BoIw4f8
SsRlchufr0zfBgcuMFVwTwzIjFGl5SUKWJTN986tA6syHPQc2kCP1MULAvsx
ev/E0gTGWHIRS4sE+Zx37URQJJcYI6VbJmG7T6KruVRemvlaNj0ZfJ2h3nS5
hMEq1OuilAC3XMSPa48WiT4XcEZxlCJ6adspoMnjeaSYOdLqZiQGt65hjBgE
rcxCZh6M54oRxt6ucF09ciShjqfELwtxb4SEPKV2AxGvlnrtw+4V4FnuynWm
LP5662X+/Xh8rFBCD+SHlEYCB46Sw5p7dWG9bf0GaisqFSIofRTPumRgd1gf
9pJSlopte+/c088hx7zDvKMD8g+m7K3WwkMdrU98yjpFLilBOmAVy07mdfMb
pZWV9kkmzWvqdFq7xjCdhzxuu52xfXeFpKHdH41rZyMRv4zILWPodU1+98kq
UPa2sJIP7sLYqjYu7PYljuq9PCrvniKpwKbPClDFUvF5O7ud2wZ4HsCfzyyB
L99PsuZiy1EJ+/w8jF0HluIRuT1lJNciynrMLroEslwHu839vLia1LTmhkj5
0qjfRWHhwpdolRKKAJKNe4BbZ4OXYY76vpJ8PPC3LiTU3u1WpqI/5QL1VC/s
MS7IalsbpXqaAEeI5AL8m460z5j3w4OWx4yhG/xBkyJqd1Qb1U0AKSxTzcF0
JfBrsbIZ+iQbcn8ZI0aFHXVX6gNTxlIxw5W479z102ichipeTONtrfsxY9UI
jJx4fIfiDA5SFd/GY+TuPJWuDCCuXknim0VYE2qv62pRsCIV/uq/0oXmmZv7
sn9kAj3qmeZWDJcZ1qdIheY+Bjz/7PfSGtDz7vDJrZoLx8JwIbhUyRoRlfWW
sbK01ncIGaaQU+guWwztnS150jXETGudixXGiAixRWL4Rp66eWt4Xsj6hH3B
+6gvAsN54OwQtYxb0g8tBgaE061kA9uJbkr73b7XxnG6BuWct+rDOyanlFU8
ZAtm/8Y7FY8cJp++UjteMyGV71tNAq3Tc7aZ9WueJG2g+6hunyRkgiDwnPUy
e95aN/e2x8oCAvM3O66SGUkI6BDzMvCLfKCYbkJsZotJURPcyw5qh59wR3Sd
U2YFxSHmTTEQMlVGz9V82KAjDfl1Ni2Ei6wf2zJiWDxx1MZPv4hDU+nknp3K
arykctzMVDHL9w6VYQU5PqCEcnWShiR2TDDCwKQ1MHOZU3dhESQojoMPiS7s
a0aTeIiEAdrFJfkM2Z503cHv2ZPuLsBFoFPw/pZySEZMGb0UbYbRBQyObpTz
ehBpYL8roSka+/g2rtNEL22weY3eRsGop5lr6b0rz2r5KvQr4XLe2wS3OJTH
ZW7SXc1r7KfDaqXlhm5q+H0jJ8zJiTkQvwogQIr2jfF4Gqfo0yIZ5pR0kkKC
OAVxUP7c9Gfq0tCwlSIpC0CSvYa6l91ndqzkFkbbDT0XpCoQO5JkPRP3/umZ
0tVOe0kz5Dzp4zBK78E+wzl1QVsGRRojcFTiJ0WrJCAg4Ivd/HGhpikWoTDy
RMbLeavYROsSNUuBOAZ1zIEfdbvxtPfGTSn+0XnpiF3i3jdLGZWtpMausHrI
kPouqmKSlrE5dzEhhqQmbRY5x08fYAA5atmNcqL2torZ7mxuvdVDOoG4JfFz
wLVSRtqCHHON2GMlx7rdmokc9nldaGnE4O1V1iDfVVNxKlEVf1ztk3CN/7RJ
MrhBQd6SBhn/E4FGGOrA/pbu3j/C2gspqfcWcSlYZmmsmrRYoOB94HrgqaiG
h20q6Bhlq0Xq0RSfi/U4eNj7z6BkIw5pMf04mk/YcifRj3WdQEUT5jj/CPnn
GzJ7YcU9ZnwQLilXmoh4lkewfDIJdwYq1BtZ6AiZI/9ycMYLDh+oz4nMEliw
Uz130lYv5fYa3QX1T3ShRa/Q1ZdBAK+rXiEIYYXPjpxGQJ+oNu7wcAJhYdoY
8qpBZ2V1RhFzZG9iyug4fR7YW1IWgeh9sJFmAVcZsPZCXJuOQf9WEi102v8O
INfk2GMwauQTKm4q1pYuVcKalVBQk65FxSdrOJxJfyLyF5H32zgrKYalQxIF
3ZsZ4wI7G7NjD0IJj4BNuebqpzdf00TunjprTT4OY0sFkiyokt+6YvdAisF9
RmeBx8pbSx692iAwIffS+8n/kMu2C+xrDHftv7EQF4yrDBueD5O/kExryBvI
KPAhZKgCKWdBWtk4PaLuypphBDSBbSOpiafn1ItGATfB+KcMCnuAWt/t9lQO
QUw7ZK0QVIJvq70uIfqXRrS3bNp9bUQ5wn9kG9ESIU4l+o4dEcgSei4h78BX
OTihyhB/tGH4EYRJnh9ZZqRVH1yCJWbEulQ+Spg0Dit/i5BN/bsUveAE+SVY
oYRW1x35420WN4KuKnn5cKEEj+FKt6Vhr8NgAE7+5lTRbWSOrey3xJvYZA7n
e4+1G23QmatgGFga/PwRpmRvB3rOaeSjGiZV9qlycX/xRPKv5f9qLdm01xgc
V0KLTMDlflPpDzC0PTYOxNrUCWYsFwj2R9JDvzxW9SHL5wLoItxhd7oU1YMX
vYoPT3Z2vZLyU+F12/gOSGJElN5GoIyeoGLgnQeOuyARrNHo/8Fa6WW2KL0/
m3wftY/ZJ5S21jz0bVdiDCflh4BLtPqdyHw7+b+xm+Yprh2yB+qLAnTtOhBz
CzYI06tNd6KnQAlGMeLYdCTqR/Pfl0Vbn5eEiSa1Ok6/LLFmQTmsCVOftscI
xYkNglr/hHgfn9XRgegWwvy+3yhzRk+KtvhXwTGH14mo3mCWhW2Pp2ImYbRH
Ykcgu0EM13USmM8pzFlaNz83T/W8wKMV66nonvPTL57lBXklXDJp61r92Txu
YhI6hed5v1rcXYVvj2DCKmPhCtKzwRtDhh6DAsbcaELa7OrT0Qjz5eE1bhpE
2nm4uDa3uLloi35fhhUCKRm/MMfgv4veoaYWErQJjNQpuQRwbKy/9U4abEtS
c6uHem/3IXMlH+Tg6EzJqeGtAwhz9/pMHVWJCJDlnXzlKBe/T4vXfDrsWty+
l5tnBsoqpTYs9JP7oRqQoBd1yi4187adjIuxHlsPxTBkOy0OR1E2odw+34ss
1Y5hOeiaKoNmn5ApowB4O3OIK95Ug9m/5BZwBHBwEWYfblwqYumUqKKZyK7M
gw0Legpcg1OPpzSWJiYoLlI72F6ZN34+TK7a5uCzs0vXkNjDL+RnBOYz7sKf
K1g/G48ILsA0a10a7n1We0i0gRBtRHpeqVNMB4yfp04roijuyUC073nDAaMA
zxjBKYieFs33SICsFYc+Zr60fadKPrsjQmCb7cifuyIQ2Zz8aasCs0+Vnf8l
1uPOx9FiBW6NuQpPZwjSw7KgX09ZW5/XLV5jBDyaRvaXWahCXsRfio8QPHCE
rTD+E/Z1FsxaNC12dapQMeO62AYUxVWE/bNkKi0xO3K8viFF3Iw/Jm4gIpsl
neBGOSSw5xklbpHJWqBKNJX9EUbmOCwzmWfRgP6FxOnpXR6uszxk3KvZCG5Z
DDOT3Eu0czvRdoCT80dO0CHSvGMGZLd5/ABRNg7JX48UG5yt/S1UERwq5rlj
x8/OYF/m58+0VVUTvVIGS5UZ4zxsNoedgQldPrS1OZNzv0c279rKeQlT/5I2
z/xFuweROpKWy8QSTSss8A1Q4sUUob7Y1w30ZbVu8I4f3yVKcpxo84LFRzEa
R8akph8Nsa7I2TDZPSKsrtSVoSgj+Nc6i2ZVBLkjVrur/uZkPmatFwb/T+wc
OeZwEXoLKvX5OIBxsQ/gLJyXcwOnwpyD8aVePYGgLFKfE2+YJbTWy0c/6UFe
i94GhEOq3RY8/OdOH4YpObKyu1KZ4I9XXBPx7r4od8kuWoUS31Esl/GCL6I6
UrGgfrZb1nAALoeR6y0sLUZC3KKqgg6nBcuNaa35wbDUEAn8TbucAw3+A0t0
P5NeSrE/9Jk6xg6e2LdppMSODTVZamFsYrzTmdOhNJse5/uuWodTGTsqVKCZ
weR66ZxUvb3RKD9peo+ws+nQC25vwyx7h6bUVMpsuTprCICld9Z1tZeKc7Da
vsyoaOqqfGMxGQs27mTlXX1GLYQEfcJKM/kcHJpG54S3/EKLzn1C6lYjFWNN
ldylruwy01HcwqvGDv2v6Vnc98L3o4RB3IOG7s/W03u+3O1xjWK/z0cix+fR
ib3w8PSlxAHq5nnyRfEMD+AC5Fra1fVSxm0At3ipPc79gddiLSdqJHiedv3p
I3/BW9dOwcfsmxa7PffR9iB0Y176USkJNS4oUryZ6ba5Yk9jR738EbduNibJ
y16bUxfT0Qw8SJpRO404hlnGYlaPsqLG7slmMr0n/bwbAbj+kdgy0FQBvHhz
H1+7V27o228U0VJE+cvb77/t5+/R5MeVtfTcq+uVk1kjpeVZSco+HrDecxQ0
VJ/pbgPz5O9l8hLEe0qeYnCCr7QdHuxw65MTOozBkt2K+jvOpRdH3GTFJV9g
QheMQoy8bHPE2cm9JO27QhowjvrOJSbbNHNEDBRbpQQXgsQIV4zdFp63p+Wc
3qtoVm857ba9QPN1nd3JePajuqSLEae2QtrmxfKIfz1tv07Q6hkzkoMEXdqX
+Ta0djNJVuVtUUnSSwUUAn0+u85PRkJ6R2ci11WX7a0fyhYUXEXDMbE4ghtW
x6X5Cxoj8LvI6hX1Uh6ycmSMiW+884FNeVTNQ8GLwO6yq69RJbBXMIxs/EbB
hXcM5nmOXeIaWXTWJ21M0EVRFOGy/7t2snebbEDXxL7OD+4LGYu7MwcXfCMy
jFCKQLuL8EYYv16KHlslyD/ZOsypi3ShKGK3/qWTeWceooX81cVHQALghcBJ
64gUBsEndJOqziyhygRa3F6opydEj4Dm4JeYAq2Y4BRmOKQu1HMKBU21I+Rs
62UQdMYRQFWQjqiFGGsTN7yztBCEvZsLWlzYqSsUcvyzBk3mvZS749FIrYa2
5PwHiLedRBr5ETQ+yRYLQw8DBh7AZ5b1GwuW7w4gqmUcqpPqFurNeOS72PeQ
EkDOf6SJzv1uI+UeDkZX9Xg0yHP5hJIkH4QKYMDRj04FOHjCzcKpdvq68rYL
drAskQFYqqZMu4/++ECOk/CxmHFA2swZeS4LC83w78qho/liSXiJcjM1XOXZ
xREdlYtFrMpLFDjJqqtWGHFYWDlxKc794cePiAZL8g+TTdwku08hLaop8KNj
fUoPNKHaDTRN0V6xEjWlnjLWa4fPJVXS2o4iV9iXkUNXlgnWFnFkNuZgVEtg
G/58Xu+f6UCTK5JlGkVhUk4A2qnSGVwW1PKuuQzfH8Gtxg8pVPBcez5Uf9Op
Z7OSxokSgQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfS4ymhKSkoV0+dPFpTeGlf3cN8sDAK4aR8ytm02IKHrMzdcl2wUloIoMExb3sw4FXSOOWnBLDI+feZEz/H1n38FAG10HafzrB2S57nQaiWO0RsZ3fpV+ZgVLAvmocutT8wjAeYtyEoPcDdr6NCQ2/rZbjvYAu7cRBCPo4S5RcEdNXkNHqvOaG56Ww0YPZ3AsttvE4IEkoNdVL9ciXsxEEYQ+Tpj1IVT4RdjDZkEGAhJJbdZMM92S6hCxTMF5ttuWEs/1FY4051Q38XZe1GlF3Y9h6eU3irGNu7mcObZdWgqOOGJgSkLIOJVvvdMnmeA/AMDBp5CY3XpVUc2F6/228Jwo8DzmXgtLEsd1TE8/YyAC0aLKqSqIO0MSxIniqzbuItpINgHSd4NM06X/eiDle2SNZmq49TNaZycU/VYO0xFLsD46QprikDx6U0ui45/CErJxFG20inYg3BN2gm2NT0RIgbQSy0Rzz7mHhokFyOHdUi/mARCoZSz43QZ6hNuyljyzZTrrGZFxuxkKHltpKZ+e44yhjOsZWTrHOr/xDjlV3uiKh9soDK1MaKil/frdqMsGkpv1GGQX7atKZD+iVyHCTJsjDAa7ccnC8aXxBIPcvD7b9S8NEi1YJhdZ/MgzHaZTqhXLhh0P33ZIZjI1s44NHuAUW+ykUrLBuT06xVjqtz1y7c7jjP3/Qs/CkJrul70Pjjyi+cr4PuT3jZJO2t6Owz2gTMqAD/L0A1SRm/rpvp7oNocNsHCwN2tRVtCq/Xh4E6cgclWF8vKt2xmye66"
`endif