// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KjOKqEf1H1qcTwiaGDVRGyMrPUzW2RERi9MWZFHM75+wkE1K3Fl49hwITgC5
m0k39v/PktoTH4EYV4lyFXTXU0ujVI0dJpgQdW1CLjG7zz40ui6dDExDkybx
JjE/SOzrUlGe3qjwFyTMn9K9RM6X3/OeP4/0/EFRS+en7ppsJ9SJfLF/Vw8H
q4Z4Xeu+r+cMfY8QoamSAYTx9raYZaP5ONPeJgY1qzWaTX81Z1nAubXSV/gc
frwWR2ffYLGnQ51eiJTr50cj12XM6QVGAIJa4R+t9o92YdF2L6CR0PIgvn44
9XngCzXCTc25R7sSxj9XsaGaeuWWeSwPGdpSM6civA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pmCqZpWwSVlJl8A4m7bjtcKJygVxlD8ea9yU5k2xWSy1Uh0ezj7MSzfAssOm
XZZ18S2iGLcLPWCS49totgxmliCfCe0BU9X6hsb/O1dF5hax3bDsVCYmxBhw
Ol4Y/X8ZwbHHLYSNO6zkNNrWEYDinRVWNHIciiBTazVzhctQz25NJBeAnEom
CJITjdvY2Jee9o4tayd5AURIXpQZkuAFfc9ZfNM1ynhFoCwPe8YeVzSKTPto
qwo/OdL5yrvwF03lbhUB5XrhJ4mqcHyc/jp7XSNb3/NDC73KNWJGRirmJyho
8QWKxW74LGaitMkokufMOWjLN9L/d7qZ/1gJGCmAFg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KjVEvs4bVRfeKz9Z6TXhEYps2JSNcyE1F9/QxBV2VFNob9ZdQBBbuqs0TpEo
AP5NH0OOr/+VWLaRb+l1pme4Y154u6V//nuGfzbAfGw2ezm/I/3D/i0XDXQu
k2rRrY8HLsxRl/1q9K9BahdOqi4CoO6dwoeGWlT91/X2vU0ZxhTDlMp8TFdX
nfL2ibfo3+ecwbOjoxxzUTs1B/J/b2+k3vzG44p9hmta9qXnoAXbOzXGm2lc
g84M6U6MQxseuuQeEdmr5/LlcrUA4jn2GbjrwKvKPghhv3yb5nwNhfcwGv+i
ijAbA/lsEzaqjRs6X0x4F3aB7e/tKoA3H+ZpSJ+LMw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
PG3hRouBEbaxsP1JdhOhKilR/2sLlMRYQhT/f31+ep3Ao4PEHuo2dw9qibI9
KkG6OToCmDnRUtEoH7HsgklUd3eci2tbONSZxVKO4aKBu2cTsiZpltKefBVK
bZTbtMeJsTc1nmsh0dN9fJoMEwWrBJ/FHZvNl+cbmvUcEHBUQig=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VTkhh77uv8OBVKZoztNdunoLY+CZpWOJfl7DYXUV8t5VJpbA5Tt8i2b47LjD
ZisoHbxmMXstfz8gkBgVVKkXhvxTy3u6zn8vHv67AfDdsTI/68g4xLdl+4Rm
rkl6zTUOvM2s/JiyQ+7henQZMiTGs5kP4uxDnx7JMLh3psRTGjF9AsOgTinc
pnLy3O7JASt6DYKORZd7seGRXMyMkNKLwy1UQGbDzS6SNa88bKBPjgPsLsA7
darMgDdPGmpcQtkA+E4LIGFexiQOAIkZQweX1V6QE1ZQTVVRg7xwD8uMKwnh
9yAJZXag8X75ddb86VYDtU5exYCi3ErMfg5n7uM/Bcc0WyqgwvRHLe9V2hqM
6iV4c2nMVrIq15iX3oFs+oIyJaEYTPlTtIekvebJsD9SAQj7f7Ui8Ads9X+h
Jdz0CjhQJZ5S1ofIFP0L9JM41sbkh8xOCPXpagUkHiDjy6e3EkbtvUVXLgEj
wsSxcWZO9qP+3JhVoY+SQYLvqxbS3ax/


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R5tiGf2nAYn4o9gFmd5P4n12jVbUUiaRau8fWCP+6IR8qf7XhsP4JrfGp+56
QiTpK9++uue/3gN5BhIBNMhgRIzL7l70qnWHOQaj6tFqwbKVJFtTR8wvkeq9
dMYNEFNBs4CLuKyops7UsDItMxmtnU1GSVmmPfeqZ5HlhD7Exgo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HIA3QzFG59lTm5uMRdsa/vuLLtvMoDgoUhP1QqakZX6FEvmOOS8NuNY1/7SH
mOo5FzGg6d1sDah00Pp1kjir1oVvxyiApe39ImoQQUlT0hCWFQd0IEWQcNCq
HPscSq2tMMDPZHvN9vH+Bab6aPiApfi1s4rZpyPLW6bHxXX4rOw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4064)
`pragma protect data_block
DAxtt/v+YzxKEWWZ/0/unrQWRJqN+Y70XLs/Yr5pGGO5QHi98XsQMU6uLbch
qe3Jd3NqmAGiZntG076dS1M5c6OwxzDKxqTaR7rVNpWomk4u0300aYwObZ3d
0yOHt8FnMIn8po83TfToUp/tVMvHNQQ2Ol8VI0DjBVPauHiBrxCvQcojJqd5
VSIEPQ6sVus3CCYGxlJR4OnftkHHXv4iXASy6bFT7a7CXuiKDZ7WmA3N7gGZ
BSAAfhHz9pFh6T+zOjtZ3EzimimU63QeFoVbvXJSDAd8UIaJ2IBLi33zbCOP
o0v99qkKmRyZKjsBM6JX9XNXfnjnnA87FqWuTysvOPhbqVAOP4dC5wWQ3KM1
hRcfna6F+0FAahK4Zl8AWaVgZyaMDZr5NYRJam9r9y243HMTeGeSUVVPbeiB
vvg8cHBPxUhCRZM/SDn8v7v+5JAFGSS73+JvmeVxajMELLpZSfNFJOb44NJ7
v5sr8fxWoKYKGZKAsh3raFYBO+OfTmjgcUm8deqwpZ58oEMbVlmSu2j8z9HA
dtgZ78y/IqcB22oXiu8SHr7EVY8A99PS9KA7xY8zYmhDcdU/hRoX/D89G56s
kjowXSJAVcqqjFOpySxiY+kF/Ub8ZqWJrOHMyieHyrgrJ4Qr9elvOp+xveXj
t96YmjZ3zBx2LfSLtBOj9nnb3DRZZwW+QVqrXVh97QzSm+Y9t3bxGNylmwxL
j1S3pvcCMPsKR60ztfvbhau387g/7MY392XSOEgFf+S2SuyuPzsYoZUUoKCT
aR9ukIXEwwBUusJhG+EFGiCQmSRAJ7rWR6a4i++tX7fapvWijxoSAb4dOMnI
+7UuUjISpXyJ4ZrMS+dcxa0oDFaMNEwai4BogVT+CL09rWjHuQSI8/yuCaTa
NpKRw/R8ZbMfqkrb0muGIKQTygl+nZvmqflmSHhSWuiEIGEehRu7zSMDp9os
rNfunLVbDABK5IhgmJofuPoLARz0Ddj75X2Ow8wDQXHnQRyBzaLbxLi0+5GA
GocjkDZC+xwztF92HAqm0Gut5Bk6FMfn6aQ4OutEm3ckoYqBzU4YDiSDJqRx
s46Kyx7a2AtswzqVA4cKEPhiLBL/zxNYtO0W6Bt9kwz+mKQ07QrAvXxh/cfA
63qZozFMHtAR6uwvQhHmKeEZATYD4QRM+h5xDo2OwqFRIvFk5z4RnWSkeZqW
3tpnNqlDik2V8BdLclScCYR22Gqsj6ILZFU7Ww0U6aQTXdYKpSLY6YT54a0D
l5vn5nnvDZs+kZzBmGSXcJQNnjo88+HqOtm5+LHs/YyROu3dszVxiNlgSh6w
xTkXx1V/Zd70w3qe0IBGfimbj1ISZusZ9CKDXDhF+5qjo718q1+0IvavTiwL
dHJmTNAeviaT+ZYPFJrjfvnFZxGHrcnrOOTrJPUnUhPxQkbq1xADmyBYWxfT
0kGoewgSKm0Ft+wFwkeS8fCotQUx9Tcto/kso1nWNayCzDUkg07i6iFkUpBs
N6WYnBXfE7lrlNWU52A7slIY+eQgTyl2FvQqdlwqoIIt/DMQCE5l6B5B1/o3
Is4CHR/1WhIPtqBDsxuDggW9AE+MB8L0rh06DwVwykRHhCraRXtNkFRAOj4Z
yEvFkBir3o2+97wkOkISpogToumi9ZeNs1gJuocEBcG2doqnDuOjvvHJxrVK
36ZH8Ize5LCTzQDafC8J5n+P1bJDM4DUHRAoCp+1+2otDoCH3KU5cEJzgE2J
EQfl64PPC9Kg3zU+5TLtTkFByFIYOvnhK5V2+fahHikp+jSHXTACzhEl5Vv/
Jej+tV7gKxhKYW/JhkXMmFwk7OTk0uTXjcBbKB1OEU6U/B/+HLiqRUMZGhSe
/v46uE/M5QDhxT8uD6UW8LxLSYhVAkTynxb8YiW9UzrHQnBygEBHXV2AqxGp
ixfUjz6zR2F5IR8FSeuYqrpARAYvX7U/dbr40HvmxZ+kvkGEVqrCnjAiMk8l
WTIXitH1+xYbgr8Lh/aY9/Iy1i/ZRCtqfTt9usvfGBms/AuERceqSkX8UtcZ
KgSKfqRv30+b8cEwtXCD+IrKzsT8MQUIYLzhVkTi5SPqTa/bYKCrHP4NN9I8
ikHfAVPYJ5BEQ4e/3neKwXFjTfzb7Pvr7JGn6n5NeyMb0biOiU/Dm0hM5avt
Dpxzo2/Pjaifzfd8Ix4xbvPpjlE4Ab8vbs1f1lSuMtyz5XtBxqJnqQNWSveu
qIDHShJdqaL8BbTCv7emZqF5dXb5F5DOhGhx4cGvkVJZIGCgfc0RWbf0omYK
wfyFelAkrwLB2r7wTj3xNhrd2c2qchzIpGRpHMnmlo2SST+dIjavzeUHogoG
+KPlt5I7xmY337SAExi2EBkF9sJW1jHaud2wmrdDf1sRLPSgLQ8dlvfGmyzx
+snCuJKUiUCTpOohkm6lVAArY/S3b1/1NtwaF/RtKh1sVuqWgjfofabCQV36
Pew5989ixk694ZN7gylCRPDw+ZqJ8ZShHdl5i6xNguqpAgloU6/HDdo6CCJa
0KgMM7xwDZiZQB3IDsn+oRr5I32T/Thpr/H0EVnGDyWsGgnyrwIOYyvV2L8+
oF6AU+tAw5++KSCbGwg7x6Z0w6+rB0S/82jg1IzyX8aC9KHK7A7fq83H5fTP
0FmdGgzK1awxj2rGIVZpvjFh+VXq2PuU3pLqU90ZCjYlOZ6LEiVr5y3MY+R3
kaoh+4GxZxFyVvw5neWRbEMiTXepeftnQJnznybLRnH1GmskkJIpXxP5ezUR
L9n0oNYgNFy8rugOWAXAWrhSWN2ffzrmp5WomubKGeh2WYD9c2BYF2LxjY4x
DVvQANhl9Asjd4l0ODjgRDXiDsCzt1zBkKFnH40jW2/ZkYYffyr7NnLauuwO
e3JN2ojlOCKnDCUGbcq3vrgPcYA2xTEEn9c9i/DTtDRXWc0RESqzABonZKzi
u8QH81IcS7A54a6kFI3lmNh4Yx7oMVilyy15wYat6Vce8rE+EbafgevBQsvM
vD3aBwR7w4wF+dEFjIwsRB7zbV0yf/UGUQFQbFseK7PHFw2/dYgu0iNgS3Fl
IA8ikC+fJJe/2ngiOrAwtGbvDrp0r0F4yPik62ebKOpkfsLrw9tS+Ihc5bZ1
7x08T1OC61ATKet3iB61S+yypoxTeYdbDziiADvx6byVFN0eHJkGTzlHS+gD
ZbxMJvx++8Cqby91inZyL0TwOHU+rIVug8qlaF/uM8nUJCDJf9+WNGpGM73D
SuWG8juayJ2rQj87SSRpjzn31I9cY2OfSS6NvefiNaBrXGh/TNligrfZXcPU
w8QOFOtiehrW27fLV96esHHwbnhf2msgHAVnusPhPHdvv2aDS1JEe4RmIBeV
0LLAtQs9tQL21lDRiye7mTSPaaAYU0pVZrizmZi3gx67y4mtO+vBR/bSKVdd
56vJriBBiOaqe4ek8BK1D17mtdT6SDavHYWnwDtHlruG3fQD+6mdm0l0klnT
n9oEkLoOEaqb3tim49kONN02439vJ9UmyKnFSp7vlfLlS3/7ANLtJvAMTBA9
lGGq9mrmwizQZ5mWVCkBSX/R62/yZ/EGWvvEhOAP4mPUiepcnMHNiyDP5xmN
dGEdaDRuNwgqJRz6zZyWby5SKs7IUD/vZG3t1Z86GK8IOVvTQ64yqpElZSU6
lpsrv4b2W6+oG+weJGlREzH4Hda8Oujh4wUDtcAw+/UiEbaHOUhleC0RmOP1
ffGXpnmSEpLOrDzsY8ytgxHokOMWpI70SMusjQZdIzCzWAN6zBvhIYgUTlu/
8KnbAyRYY228zaxajR/3gtaUut1nAN05Dm5voB1s9Bj7p7bUD9+R/gCkURE7
OIpzyHvIO641cvMVTxovJgK3tPN83C4pN2vCwkux2EPVSA5ExA4Rvo9XwRoT
swbpx/Qi0gzNwx0vEFpm/tXeu7D+DSPE0+iJAH38vDGHo4Y09mczwNxYJVGH
VOMoUmP8fWVhqS7KrakpJxHBe1bfYr7yFl8j32ZzTLFuof/ugKPm7fz834Fe
Fl3oYF5fJwkgBlHpj2ds4YlFS4rRe9Fxt0WjHko8d1BDs7IIKJ65jCnY1Js6
rVMYdSnIPqfn88czQIvl5kri+RH5yo2b8cyF25pjjGXCHbhhsP5piIcm6k0P
tz3YyyHUKkoAbQ+awBurYQZe1ie4U4wZoDB+m8CMuW/aiaTUsS+vPKOgJZoU
e2azbD/VGU2wxyQrWRqYH3+OeKyrPgJr5CFH+7ciyhIQokj3omW4u73b2qKF
8pRhi0m0KnjDe3RgUzNL51CLunGMbv/nxSHfNpPXbcZjl82mE+zG/yGKC6w4
qtTq1jr0A3NoPt1A85xJ6mXYfl9PnO8T7IRaiwUIfkgeithsGpV+OOGEFfcI
pmR964imrqXqceZWoG+/bRgaF6bI1RyeVwWzrqTAZpIQlq84di/ulBZmjGrw
wgepyN5Qw67oPbmQifejTB/XGjqP8XOXRXuD/HLAGUkw94j2Yr8OQwxqJrCT
Uda06HKrJEh9IjlYPHm/wThDwpxWUK+jFKKF9M1x3ZoOe7VErz5VBX+XFntC
kKQoExdcYJBk/S/Xo5yvzZ5osG4Su/8lfVbLE5NOQMLFTk3Y3EUIOYwGEC4r
4QMtjgUBdslTfedPKOKiDFgQ+2f8Mi3MXvfCqeoFRkyx+qq3SehNUCQYohBc
VzrEnactwdO75KLLN8dE9UPyGKhBYlFdTyaNRXkiDrbBzsvqkJ1o3qiVZZlH
tgkBpQaUdwsq2lgo1Hk5AnINC8IdHAFG3dOvDiDbznbXmVxhnHMQ5IA1ORLZ
xN3AQxTCwZ92QpyHirWQ7dT0qFhdVWzkCZwXVkq1gLbiqjpOxmwYck8XigCw
Iek33oKO5Gzd8p8YK5yEHH8ZCNXPomoXhtrRfhMWUP1IWyNrsZQ2E3kMl7MC
v9TY3cD0q6sDPjOtbUB0Z8FA9VjD7AFtfL+pbHXNADYhfVJ1sq2h3dsLLM9F
cEb/hj47Xl5mS8BEiqUWQkKqkKyxW9dzTWIDVc7NpCQNwER+HVHTcoeOHsEe
m+CAzUvF9zw7qHghBeOzLI15y45jhMOFBVS2azIsqw9/5f+y8jUFtRjVaEJg
lbzIvnrZ1c7WwPR+Xo5GrL6LMizb047w/ptOFKg/vnesI9SDILz6zpyeVmsp
6MxEjNeKn2sJbPiQhT4bv6VP2g1RpqtZJ+abBaH1rze3Q3YXcwx0l3agaD65
6BUWdH7FkAyCl9fpgo2qjqYJFpNFj2T2cmcP27TE/LwlsnYL76kgTjxoalMv
/yER3rQlEBcGGv+XoMi6iMOi6dG6SkO695WfG6Oy5tsyNOUiHdBfGp7v4dfI
dayxc/LA4HUQeUlTBuClFlb0rwXI1cOjr8xr8H0F6Yn0zZbXUud3Y59E0HYZ
GRK4Pv0EAZS3JEZ8dFI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "t4xPJbmEH6v4SVL0gN6FMeKrn4IhP8uxgDEXixmWFrfkRmUmHah0woCI0NWn4jNi29PHRr8qC3E+56ObAVSYSIpu2luY1Ux8HxJTmEZp8dfWiQKOAKoquE/rRpOs7kTiASgRERfy/4yFwiIwBiIeSiYycsrshs/YcSPLGlUvkeFONkowA1F3QkwXAeAdMdMqD0IZHCYUiyRDun/uIWwwqKpaY0MedDAF1dXVq3jdOlkqbNSDZeUYAkDYHxjaf4vvQHWRRaHuT/tJVyLQTWTVUKEP08bEwIrtIuIix7uD69I2RiwaJFo7CcyoEN+fAc2F3GZ1JfgNiUciDJfG+stOH+TyVy7CGFF9ow7eX5Tkj2CifXOotCx62q0CVftVa5Ue10aHaXlfYbggOpFgho0MSl9MIbPrKAs7EEk8Ws4Fcw3c+UY5s61H+IZs+qdVa+JfrengmSikoEI5svx26o7sLrnJ+UmJOEsP8W72R4Z6JlTvT8FvfUY7/OJZctMU0o+mwNmwuEs2NnG+1PtMUmBV1NxaZ+/6BbIg8tsbnzTxA/fGOCBAkk87L32SVnsm6eidg6JxpnmVcKk18xanNpodNn+M7AFsqNTmO3o+HlO/zIK5XxHvlyiT0UpNPTkAnAzpY8RjvIKbwm4lkzCOw5gWcUe98Nd2WW3AynNAzg0fNW4SPOR6POlTdIOvW+oCJ80YJG4lJNxYc9vmJDwWRILF9b4T9kqZsoQKhnVUl3XTtywUC8VUZJfPFgPNniOpE2Ry2v7HHonq1JJCT9/13UQ7RAkw09fdsMXSbbL5HWKViGrzGQxiP32yHlJ+37xeT1Uwwe4i0woXUMYcn/FMwm4tQlnhPWrPH5B7bhrkqhY9Azrnl4do+/MycZsONDGVkVbUP+vmE33wNNn36iVSYj8gnPeMVpIGmdZFc7nmwk2kwRSWzWc9DEvoz+17/oQCtydyHdEHJG1LlUeTyhrILKDyxzFW4eGZWW1KOQY++5tj/DLASxNbJFJqGnGdvelc2J63"
`endif