// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AdUiBo70qBDlI8KPixEOzNWqPT3PZiTlS4QucqVnAuoy0Mb8/DGnBpeERjAp
XAYZHgUyGFUD2uFCSOG6oAfNfHBEX0A2eEvdWydhv6t329C9FH0alNtJ4MPT
hFTh6XHLHfWouulo8k2/iC5LVXI0K/DknEggSr3UY8f8e9TJ+QNWBIVh/VSS
pSfhehy8g3RqF4BUVIi9WUvrQsEoNBXvSP5jjI7F+I+kmHj6OR1405mc7rcL
Pn5EWQEZ/Lgo3O54MERJ7zO6s+w2RVt3ee7bWa8bLMGPlC/ejiZq46k7Hm1n
34AVSYch7oWY2k6BLCoFNS3ziHtCtgWWMF4U5fJuCg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X6One659dc/SPW3frxuw2stz/clcGwdVfOftMxVion7jpt97pt/RyaAJKRCu
JuXjpMkPsjAU/V3/MKgGs8rx/+vauVStZCuz24Dj5qRN4bGKhu6LsOwyGi/Z
pU8ZUpy9+wG+oJm2FO1EdOpHNn0M48UAma6a7ZcMxEaxz5FfWMj0dAmZS+qg
sF2jEmREaAXpnKwfwvIEhiVlySlcr2kaLRfOhunBRqHgYIXs/VQUO6pJgG2M
8tCANhwaTFXWLG5Hesi7seKlygGjGqkkEhDECoNtVhKIYZMmx9IRVYtvouDM
Pn/dv6EM5TOv/3S/81o0oVowa24ppDWfqNcedMFvUA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N6gB1Dv1L8jMGKGM6TkJspGOVl1qf+3xxIINBHSa1UbrvGDegMuMvmgQzhCn
boumop/I65PUyQ7OAXFcYQFJXrgMtRwzYmQxmYn5/nOfARu/LFCVvFfE8XPf
VY094uwZ4E3xMpFvm58NW/IwIXupNqC8mCIzrhFiPqcArcTxL9jhzBb34Q0m
GoEW/3q8vvyVqrfT2SsrT8GHW1DxGxlsm+o6krpbF4XsGZx7UDphqtU3qHOP
GRmXZxS6+GifWIBxXM9/970BqxyyGL8eGhjvKGwHyLCPa3wyhMIlJbKiXe/A
UdlXQ1AnJSu1DrhFKdQ4j0vd+JJoRJnXy5b1w3+6nw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ret5xuxXK5hsSixAYPbpwQ92kDMVrHS+XZZw//6V6No8vKMxU1f9up7orzEz
dFOf1yyXuz9WLFw+0IcJgmnyVk7E/imrfu8bYqa+MZwGwYxS/N42OR+PYMNr
1hDj/h+mo3FdYtBg3eN50kdMIi8hpwQyG8aa0iQIeqr5zbZT3vs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
CLes/gXrGu+//dc1MMOeQDpt+7Hhet9Hd7DjQZgsa7f+ZTSIDLoGUzdEOFD9
bIxGP9BmFzoIvjMP+0nQX9kgdLCRM8/R70XGqsgjVjehdveTXZRGMNc2mhhQ
G14Nn0Gd6rvRzblyFkX9XGUJlyKYP8uOlSjDwtQBqLLzkW6DdRpOoanR4X7E
quP1zraTBFwHknM6ckQ5mQky4BIhKTX78ZCP/S3BwJ1fQipu0yX6flyDfIJg
XBr1Zfd2Kc+VBzBrS8/tgUq4RQDmAlm09beCpnBkvDTBGHI9CWN9OLVkF68x
YSGuY0xH54NyLGuf1KcC14iOvvAaptme57EvnSQjVboH2rNeoK7CR0aFXfj8
kDYYVaYo1c842E5ibw7w0G/Q8gQ1kekC9w0uYn0I44rLdt9pF/wxb1blxIAD
KZAMMyfzBs/xf03eLs3XUtpSCRoHqUdR93pTUFC46TDgHAZPhNysf7Tt/E0b
C1cAkffp3LKb5VQIE8WUgzFj4TXbHL7L


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SsQw3/QV7DfvdD16AtcycdFNK+2KMsO+EA3TMT95hgqyjVb5tQNmc5Ue4Leb
2HS47DbPdla5B9fk7zc1O1L2S+CVucWEsyJQjTaZcByuw4cCGB3U2z+dr/yx
qw1+B8swcAA4gjASewEnEyAUXfebjUSw4I0ryiUTaL1BuvjFW6o=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
i52tPpO/kfO3ztDHmDVi9m98XzaKIK7jrFP2IXKEtwXMvPsgfI864d13L5Dw
5q26vyMGhFn0tlc0baGnxPmHq4X5QKZkZn8UV7qm9BYFjSnNB8bKos4FbZxE
ELMn9+UH1eyWXKjW/zUALbEURm8Vbp+y4b9pz7ZCHYkYhdxpIm0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 18192)
`pragma protect data_block
e9IWTjt8I8vYFzBudNG+OCyJe2YpvCReHTweqpWP1OIJ2mtIgHa5nDMuxSV/
mcABsqfy3EyLkaE/gq3s+h5fY77KuAThlK117+aftl520mJ/nw6wPwBC1T5K
9NZq3wANHbTCm5NzMo74CVYg/flE20WHG5NvHlufWFAYkXEstAPMHQNg3SWV
1owVvUXRbrFePDcdbd2ZyzDA1TEz7B8WT+hiDREgVTuJ6YB/T2pok5GXc5+w
gJn1fdYoUE6qbvfNONIt5ks6sX0CYGWi1QOC/B0OlywolS5iqnzag2KKRVau
/+AT7BQ8gj0h/a2RJu/phBqB4VKAI43BWokTCXGGv2UuY6VmXOg2GVyQlhvW
jEL30MuVPA9EoHGcKMA2X67DmN+GxnbQ9ylFMqaAITRVPfviOEOHeKWYFclo
FNlChtfEVHRu8L5xeZ2fFZRGFnIVAILj6z3+t9eHNsjb55XftkHaM1xTwZeN
Yj+07Z03YrJZZ77LM25EwKL2SwRom5Er4IMx/zfzEYrtC478QPRGQxrC+0AS
lea4qnW790B/EkwccxyP1QXuDmRsHA3Q1HdQ33sxQWBhkSfK4+6A8olXnjfl
1EBrAXYM6NgvA7SfRPJuJCDTzcKN0WH2c6k48Lj4vQojMtHwxQYxCyCG2qR5
3Lp4x8IjxsfYhkVrz1Iu9F6gZ+oI7w/Y+QvtB/0fywCsesLLtcSduzz1btaJ
Ehsj3+3MauDYAdGNgO7pDJrvP72TdaWJfQ633Z49Bxn6RAmIP8qW7Mx1u7Yu
Z/fUD7kN9UrlclfzqTfguT+HkdCMySI8MF6mEPbD/+mwz3Xmxf6M3YNSx7QA
i4vK+bKsqFS6uZLAm1pimCFIRG6yAYioZ3PkXmdIjym99lDHBoYfdSdCYp0T
qx8tjtI1MShkS/uLUEYJK4Cerkbbm51SwfTtn+RGKXXViOxFSRXU/B/CBqDt
TgBnezDEW2UdmFSaBNZOBMpAj2dsl/X0wz0YrV7QuR1tlQUv4oMKChRlX2fY
D6XvyJWVxgmDE0LR1sOmhW9Da1JqBp73YUUOlA8Z+XKrM1ArhGh/utcZwwyB
5gxgySWzlk7ec7RZyCnDb8IhKqKELEGo4YHV1YuA436lo/rb+Mqwpf9mz6NV
avxulIyRVDbydx0KWITcxvM7uCoa63MkGIgeK6oNJdnD+CpVmwwKDo1Fyh57
0vKugB0+pzradQmZgeSlVvpbCWc6YPL1jFSpdK0pwoPm7RnAgHwPocp03kyg
4vUR8mFXMl+jC3g0bFitlAfbCOJPbB1mW3GNxhmMrSlP9Zywp0D+esE+ssnA
El2f3IDLeo4SZq9i6pij1QhJqWNC8OOvfX1/EWMzombzsENCLylCA2WEyk9g
0XJsw66krQrWtWsmaf/O4RN74THokrFv15ZmRuLfEkVetjbztuZPXpEu6Fz+
8xPoWa8Vosxx4jsXJcHDDCdvojR5msv4ili0w22Ya8eAFVowMuX+ZdBLkO7k
un9mdAYLyCMPD9nsHVjx7ZnSAjNPoDwo8Kaf17A9xhuht9FSL3CPQp+TYNWl
DLDlkLr5vSdemkjV7+pZnKIZHlxycYOLPzumh1/0D51NGZ9kshPo/7vo7PGy
PfEPCUuYdbLtx+b8BjWGxLN0MnVYu+VAzLKe/mjVv+5Mx8FPZESahNMKC+p/
xhMChJkjC3a2Izoeng66xDEbzIsc1SvrLfYpsKlTkgPaZIa7A/i2mcijs44u
UpDAp7p93QnvfiautH05o5sLEKaAupeKQNYk15sjZFhl6VWnGO0lZ2YmfsC6
HU3CQJVnVr899Q3NCfiJhmyCieITgH3NyhPr73bJ9fq73bivv7i+eWbxwpR4
VoYXYtD7sjwEdjOZK5oF3C1PYyza3N9aZCm0hQ4dTS4ACf5tRR/Eo8kAde7g
yR6CpIcm02ez/vrGQokiH9SdTEDjGpHhpv7FWWjmGh0s6GOuUZNnNbh76oCJ
eOHlsH5BiBXdk0vspevItO6lz3asTp24Fm6Sv6eqlH3HmIEPtLxW4Mkf+kPw
NgNJZL9okLTkA96UimQRZvP5SGu7SLui7c+66v7n0v4U7ki5u3IJxlwjsVCt
MJxq+E5KmhMjS1X/PFpAxO4RzMhsbG7I5aGbydaVPdICEYf6RoFoI0Yps3Mp
3QoFyOxoO2TdiJCxijYsuIVod4VLUmheshU1QYgIW6LqsYWOBlOCVz2SuMry
9ORWd07a3WDJ8cMRbj84yd/sPxhODyF+PQC6iNxRRH3MXGbFPZNI5aicaC5T
y2MQwO/EwE4usuDr8fqjRDU46asi5Xq30kuqDhXoC1QZ7fBZkCn+XIaZ/r78
F2OmoMdfXQ3JNXdf52OmBIqan2stKsSBm6RUXccvJQ2frY+QAkVOFOxJ0aoI
ekt/4C3yQJPlGaiaJmquXi21UVfMSRtfyP0P8tyLFA07XwO6A0dBNVsp7hkv
7h3WjIUdx/adyPKSF2YUbHBX+UarjMfdKABatjQ7+FbGFotFx2nEeIzFhbzA
ETSvlUuWQgsnGcSSmwxtO9BbARZ1Jnuzx2+Yg7yJdv/R98i7F5mX7z5FUQZI
x6/rkVchYiXNN8xuVEQRV2lRvMQtu/ibkQKzyPOlmx/c9fEdXfR5dOdPR9T9
W8ViZ2x2PNgtGcYC7emgzJtppkXgwfdvkpgWu/IAjuuJ2klkl8i7jryqTNrO
SrdXpL/tjuRiy3zQKni0c/XEiQ0SVf65O+xayXQpBf3r/dGEchsDWXCdFwoP
urPgMUY6EsLaSTDprb65zi7bznk12YaZoOiKj4OsZzgiSxEt4IW04xBi2dUB
62Bgd3Al0vNx6WCMgMNAPkYLUEnAK+8Sa8LGntDPeYixJmbi7h8uARislc8x
uAeVZdVZMeu5Fj1M3dM2SJiTEpuiUxDp/OcET9eFzLrNrSxz2JjqYO0/pEM6
T9R1PfZ7L+1PYa1WaqD6k81JL24DD5Q5jN/9gr2sO6tYZVNH4XeGTmLtogAn
yGOmK8TOc3l2RlywXBx9HMppP4T4+Sv9phn3ff0vwd+5UlnjKHBl9n5WDti9
TrHWd5p8NAdZTyR2joj+QmoT+Er4RFSJYlSPShZpQQB8ZGBIWBUMPUPXM0Ic
PmsyoE/4k2W1EBq9DxmfgxGnn++9rdo158UtE5eYjxrLMWAT/B8wWWs6qvCU
CCHkFVe359kP0XL+Tb8BVMdRjM+6TsXjOYnz19mAv9It6e9/yRCnGUfit+fU
PTlAazoR21l4NuMQepXNsWADM91xD57zVoufZGSBcVDRs+PT+8Z0q9mBFZQw
hEY9HnvAf0z+XWxGOt6Mfq3zqcj0jtP4hLRNQPcp5ELJVsH4LG4M44nWCqqT
rLvpQKmjdKFetwjai4yLxb6fsI+UPIma7yYHVskOyQl/qJnqm7gx0nIMVjFl
GvNXWpIJx2lvwB50ZFC0NBjp4/03zv9G2QBwjp/uPjxWa1aRuZ8cj0wUKE4T
QzECP/MUcoLFj/eWbTopgXTWZWonmfXRe7HpogW06h9TClwgUSnkn4tliOrf
w8Kx161ogcVF8F9vBu8HHZYg+YYMUsv7l3R5UEJuhFy907zdSnsk+lj0T8UF
wGfH8W2ObL5eJ8YihqeT6zIPhZlhV1d9z5ONSRz0qvYUE4IYImh9ZFLDTqVg
kDICsK5GrI7H6n0Kfwud2S8Y4kvKzg9xIo4SGmdYBwIAtrf+L+Q74As98NTt
ooXZC2ZtSK5+6q3K5XEGFiB9ULvNMpzJWeopBTszMGyr1c24+HXuKU92BOxK
pntJJSiFnsB2MXdXQn6AABW6luSQ0wIziVRrB5NbGC9U5VrH/me4UFwBVj9h
NL0cCrg8+2+FCCvBLe14lNbDdT8fgcw5+8CQlfGN9wBJce40IDIvf+vMnUDQ
M54Zfqa+8CMLKo7GyQQhjvJovzaM0wD3yNkCYcEhMedUmL6QX3NyPbIPP6yF
G4LBfrZzs0q3MUfbpecuo+S4EGvZSc+sfMj+t3KH90H+fa8223/mLktfJt9d
/BwE2UZkZEWz6aj5/GE6pYPeYoetxNFY6r/0b3Ynl88ZHIG8o/atoydUyt6V
lIm6VoJcDuSbDAP2DhVffgq6QcEWXmCGVPpLa37RLGg0Z6BH2Rc1n3s5+M/1
0KRZYHUbyO+pYAF8ZJBSNLqbZUh5YSSvAy0VQfM+GAfp8ezpGr8MODkd+VBq
4yonwhH2HwDSr77oNiCukLg577ut58Kei0L6d22Lsj8KpE1zRFaO1mcbQ4RY
W0mah7rCNHnjPtOLJRoIQ75G7IpxlaaGdiAFzFxGykzokA87VEn7HxrOP8gl
DFcDy8/xXHgJuaz/eOoDsO1XZ784AVmrKZcQrdxNFYpuT3tyuxA3zQKg8H+v
8RGFSQE6tOCGabmJDEfWOy+e8fyz+HFCpGbOeb+I7sWXwdzTQ58o6B0rOA0v
7MCZjgd/NLJp6xPAqaVHWxylO6HXpyIt0NsUpYVSqLU9P6ShDdErBLDFq4Ds
h59mK4pHZizKrEcSTOjL4XYgDSXggc5ERqG5GvLyXGtegNOmN06BPv8OmsY/
v4EJkeSLId4vVPlc311LN5igbaemDmHpQD8GoCEyiNEfteeBcO7tl0wJYTn0
dx1JT/e5yu6OrG4H55rQ8EW1RQZzJsRE9bgPiS+1AZT/QlamtSBz8PWBkXlE
gIZCqbdFxT5A5MqZ2RHrm+gH0NprcVCn8XpswCjJiTzCzgJ7iyqWzriX/R8z
Tu5TtpiBXN9przk1H4rS6cjRFYrCIAITbDuZFChJFsxwiLpufsg7xeEtPv6H
rq2EKyzhcQTObFh4cnPnj6M+GkMn2voPm7SiYulCHua4zgUxtMit7AdQjYd9
9Gn8A+OK5u57J5Q+SK0UU6xGV4Jy7JchryfJ9Vgf0hnRW57WDtCZR0if7wrV
bIcE/KwIJyhIsR/atIU7ssqv5BcbV3thXz3Nhhqc+6G3EuM0okzP+9jsnJbX
hbUbVBoJevw/TCb9rcvbZ/ki/fTo4og6xsVT8gxrsq0Oo4njq4QJhnLrIXDY
g7XiHvA4DinQ5MqkJnK8wAf50k3u66fOpj6F4RBS7Ly0jlFRQxZK2JLxolMR
bjPgiz/1+wKpQG5XWDbRA0tMpuUDlc2wVdvNyL86/G2tWY+EoTfwk7w1Km+p
HRt7fwysLjmByHTVPJ+UQjCMoHasFyDuwLJ7Mk/1+brCdhMVPaN3fBFGvdlO
fk1xDUn6MZ57qAn3cbixzcvoHdjhRTVy3ANbk1sD7zN1+QjuE8mVvmjxxr65
FyUOKdwWluC1iZhXLs+S7TfHcYxMxtdSHvTpL3HtAVL8Ibz0D+8UB3u0CdBu
Yc4aoiSk013ciEku2bgPLObcWFqVtkvOEF2grCjlaIhUJECuTu27VPszXkG8
CteYUzl7ZPDD8qiiJ1ekGnGrCbUbZHPHOL1FHeXiS+yKHB24DnQXqmVgULDa
NR1+zJcuZIyBhf38QmNltaOf8Lv8O2XBw5aCZ+YzZBiUxUeWTNT+rDC8q8KP
YtSFHVdYV0SwbdP/zUsUdSHSzs4JnAMuo84QfXqSJdhusMUh4sHyaR4MyC9o
Hk6oecR0gLFuKZP592eGORPjQcbBlk6eaP/xYWBqjc013PPFQ2IOwUb9VZ8i
2OR3hKvVsq8HV3RmA4Im79LAPGHnePVELGayy1Igs30bsLlAuFVJLk0IedKD
JTNYFLcY4UzZVCKywnRmYzbXBtFyC/htkhJWi4y0lP1zExTh00R05T7YwAqY
1yKtm2W761ZjaaHUFLh9Zd09jMNPVx8+AaRpVIOvi1JuJ7mFg0dZCZ/mepe4
CNVskO2sk7itSC/MWRvwHbBtvy2JTSuou8qEjROIeOEpX3MzAnzxWmvgheU9
IGEmXJwUIdBN74OB4fEm3e2L7rNcoeiN35/qi9Mfimew0zVrzbtHJsHjlw91
k1pkUoUlkIa8Xlcsg7C5FpxVzfR3f8UGNDdtzUB9wI8gcGUxiIL94pTCyzc7
ZYLpvKk3wSQXQxVKlt+6+0uZp3c81hA/icScASDdFTcPNgIrZIV4XYIZOWvB
oDFkCcagj+HQbnY6yWL+1yT3x3qBVRlBtFFuqYwXP/nkHDNZUx9d7R8r7qcw
RvHf92DM5PrxcD4KB8o/b9JmFVYjH5R0InjWa9bsFpYYniPsRaoyrnmbBhpE
+sbILu/eJd9SOORoL8DKaaejVo6z2sEUjG1/mslMKLdauSAIsKPwZAFu90Q7
ue5UfQvaKw+t2LH2CuT//RgoHQHOL7aITIBUt05sjk/BA+tTjCvzBJUqSU7Y
0dExIUA3fdBfQXMsTUAumPt3Q21JUo5K8wfs+tpfNzbGvCHXVIZfpX/O2ljT
12kwpK63iPUqRm9azmdFYySg2OXxlWS7AXWsj78ydolsI/+M6X18dUOZvPzG
1oqjIE3PcZXZjc3Cxvgmtm1NXdkr8Rca3GTrtFFsEebRnE/+Cwk5jI5Lp1y0
V5YNMlIBneHi8usQqML38G0M6+qriFsIt7lteh2DaZ6gQQwkp8p4jpNFT05f
48iTtfeQLx3n7OT7qTS0VO6CJqp12JTXPHCqlm8L5s9k8mjNmitOgjfG0keG
twRsOC8PTWv8e4qPobs6sE4Cs86fSYQkZ6qEEKrI05GPMAZhhPIebH49uiXN
m6faaGh9CWz8Eo8Y5zyqtq35EkIfxRfd+n0r2evdL7wFLhnyHcZuUVUp6nRh
mi5FomPctdHenctSjt81a8m2hmTNf0DcHurD7irgTETuGcMJjyWiqhaxlt0N
1KtDh1NtZV4HzHxpLlTVxnmuOoSfHLW0/oncX5zO7Mys+dE1h2XM8D9jG1L6
yEb5S51ti9HHz7pyAkddWrpMWqVSYFYJHFRysDuB31sw8PKOCrpAg2bWxbMF
hKZWkkoHJbrU26UO506vAfEEhpxRioGEMBRc1ro0X0/HadN2epvgxvnrJbiG
ygxEgva5zK1IbnGwNNm5OP+yvwOGA3jatK4OZvpgyto358xV2lBTL0nTpIz5
vfwBanBvw5abd7VPIXaSweezLMKCWLxtLioOKdhVSQdEjqdT9VyMezxl8Xim
5dzZoEvcnMba2ikloegarAbUIHYyiOV0AC+kc24oj+daCI0Euh7M0iv+Xced
Ovy8L8KvS6kWZZVYOkiUCZ4wAJcO1pWVC1IfEQShE8jB73Jb90MM5slsqN3F
wUi3bu+km4ZylR86nczDCaGMMSclL2vK39WEVNY/FUBvDb7tedeo+Vp6a+bd
tpCjIFhi/3wlDet0/nMKHRAKF4aKCzOLRrLucbGP3f8M1ceNz38PyU4hkrXL
lFsw01dQMnALuX7ofZy9KdEEUxZVOL9KZjBKV/W6RF+L0RZRDEG4LrPLtIIh
uQ8LqXFoCwEA9f3HtXPaCuPlWZBvUrgO1ehg3F/rVE7CdY8f9DrZOYrTNSYA
HxG/WQpfmlQS/wEYpYsxv2/KrmtaBLLQiwW0ytgSsRbNMR0gT0w5+IXRhOiN
NIRicG3j+cTh3sIjgD2hyfglJcwU+Q25ijJmYnLAzNLt+PZJskSXGKTS6nhu
cOqNk935bid5fVicySUknOTCOghxkZYSihIGiQqqneoyPtMfIwZ2VioGea5R
c0udtall14Tj3I+2C1b7KYBuJn+eXNxc50YGSPP1xAdZJ2V45Aop36UvG2X/
tNQ39z/m4+3MgYYPBA+3rFLBbwLCLCBH/QZvx9MhdZdyIw+VTnkp5cOgWgbW
M3msFK3nBqjacBPA8a99dsINEvegZDZbgpfGgtbE1l3VQ0GhrlpXf/8PelHz
em6t+9/pdwpgkLXfG9PuGl5kdVsXtwDdU9n34RNEDiUsSmIE4l5Mht9IWIpw
guavUesOvIGTJ8+/n0Csiv1rpMbhBdWHXDZ/crs4baMPLM+Gm32oeYXVq9vX
deI8LF0n+FOr/yK+foatN8MtaTemcftFRgQORHJy6SyjSoXLSlDWidKZymEq
ZUp9OdsSGMjLWrL3NO3Wz2BMXj5C0QAQydE2uZD/iuPjBUSrUh4ePX9sNca/
tla08q9qcREf/tjFgNdYOI5QSDKce6QPNgtYtcmfw4coCHPiJXBZYEx7Chf4
y7kKcgkqgyjiMDL3JySuPKJr+p2y0alYHMPQ/0DLTxd2l0XCBJTypv/mdTjZ
3K+P8whpdOw01JlsHZfrLRX5Sl4qfPF5eK7NNICl7zoyGVzrhoQZnFCjlPgs
Gi4hyuZDMMb9Ey4WSwckXTPfzxxENXTRPzJzNcvTAXLLhlv2ussXbKhvrS3d
0Lx3PR9ELNeEOK3rfIuhAOg5c6XTW22wbvQAz05M2dF7DPYPpqTi3gBsWXgk
wok5ErLIUANoBnf/cI0A4K+fJaB3rMfARHO4wy5VpJ/7IjZHDELaOUuMLfES
2KTHnANef+J4XZXi586Q12jt01zfXPwUpdkajlqhVnd0SAPVzEsdqmRAfE5t
Qg4ijchNyz9Syjh+lu+uOBGK50V7KEJ/g/l2VJ485Om7pCRJDMu56cSICaTG
OXreYdvZ1tAeLLHwc/Le3NIq5e5fhRjQbXLMHPeGXr1b2tN1J6mol7/Qeree
Dh5dZj0zuP/fTymyjIIsQjZD8iZ/Gpa7WyNcYiqBVE77iPldgCREqiDVUFnz
OpuQW1OorMYERNQwq3NUR0uhdWiGJoy8/3ql6njNUFM7uAI2ZBKEFRfg56hA
Qxv8Zd55XuXsbj9MVWd4Grd1XIl46Tz1Nacku6FFAJVSrFPCYz+CPIYdU0uz
1aKmno1m3dgj5AgSOfZo/Ne54uvRF2JipPIf9uBO1c9RPUoF/0Ez7NQISi9q
63CS1DAFeVJgkf4avr3MuquZcd1DIAzQ6QqqMOynGyc1UXCwKdhvNMaWnVXs
cslQHzRUlGt8rz/7miTWSnDcXd9EDZ2kq/ms2m3uNa+AOyg7MXMdd0X6TofV
IsixURyK9aINjKrnNz09bIhvI7FSP1bmTkc1BRRBiqRNuSGPZrY6cgGmzZt4
BPH9t2DugGAsSpDyWRFsOdXTLE5p4nOrbeciYWqJ0GYcpKfgnXi0WBlu7Q/z
EruzVwe7sUJq5vi6ke/KwgqqAVzg9EYaRfTFlqU9TBzRIN7Gd5qpBuYC6u8n
cNrYoCFd8fysY8tUXwJwE2CdSNUJxqCFCxB8Armw7Xgm0IZMpG1x4VZ1Kcex
grBesuleg6o9d0I5gDu95dU0/P1TDmGGeK7hM84mQ18LxO70Rcu0LW2Jgysc
t5Uydz/nQJ8N0OnVrWzwHEoW+LtkofwTogYLXpZ+nk3z5Ol5T1A1h9Wd/Jre
NquKFXQNW6OWkmiuzH3R/cw6Ld44UArif7PCPtC+dAIqlYo/UJiIRhOJ5Gy1
E3k9TufeEq91K/KSh1Be2x3X2akL0IN0samOe2a+J/dR3bL6YtTBxOWrjLgr
OryqV9kyd6iH6HYlRxrplXQcdDIomj4/96JzcsBENAWPUY2wvQ9PC4CgB2R0
yOvoIQcNqggIHc5NaKK4s3S4q9WcJtJX/6FED/q+WUJmcHHoP7kmFjdksAix
vYiiNYbGnOFwWXy8fA7psqQtJ8e/4gYfIbJEV9ioZU9pp15VDjxA2mZXEGS+
m6V3B30g5ouPtedaWCBjwvbRtMffT6w6XF9DQWQ+ByyNS9QXDv5Vgp42bS4t
0q5plNPKOtrNk265giD/c9i4g2jBWQ8s71ibmMXBrouZps8jaUo2C10h+WtW
FJdooAi2FGtgqKk8YiyvQJJeTmO97GIFy71ZMyRNNby2fDWh0CdEOveLv0Pl
ueNy5ahB6/4KoPVJipk5ubh6NIvuH6Ys6vHcWFjDY7lxi4LHs/acW8tzJM65
3dbk/4TPCqINLE9hdPC+gQNz65NxopyY5GxGAyDODJy7wzbrfmXM6+9+ldiA
u1DbA5ha6SR9g9Qn11b65KBSs0McVKZBmbeVh1J6khjIutQAsVvyVlGgJ3we
BjqnORYgNTHzY8HFiaHKCsdsX8OOy16OAqs4K0zCRbv1IDe+nRbz4pT08MQg
VDWJ48Zntb69mNHyYtbtDJ8cA8UOUMlFDS1Ip8mOj915+dSYpUqVDpepyIfI
8esJZHnFsangkMYORSc5pxfIzc9Wiu9RTTTmj7rNCSYYPz9ps1fwPWoFndd1
cLR6gy0ekZA5Mm8MwNWtOr2UPB/DM7g2sP3E8XDBZSL1pcpCXt3ibKNut++Z
lpU9SsSYca4xdPHALTkawt6p3/JGjB/ibUr42Q3ZyCX9uHSnQjSCUNtkIso3
WDeueeS/SdoqoY9G56Iu6hyMvrgEeElaGQqWblrIWbU6/ILtEOP59gGWJUA6
7vEYjBXFw1CNwP9Lz2gNYPaVR/DwcvG0b6esLnCNMWukJC2i1zsJv7WLZ0Ay
BGGDKa7IBAqw02r9xZ3QLQn1ymH1OByaMRulJTZmKoK9wFyWK4QuH5RaJm8m
lHZNzS7XvDl8wwuZwrGP/MwpKvM4R9rxGSDMgdXG0lZMBPQj5RPQYNpT8LEU
sUXg0dtfQA2vX+6c4SgTY6zu0L4ZHXT2gtZfDFLCAquSFVKVZW/RCnsQoJ8l
r1kiZtfB3dIHVmNtsBLlWhkqF8algBezcC6x8S3mSatRacbsKAH8i33VxmcK
fpAt7rYBb/R03gsgUZUd3rYprDM/23Ywbx+h8XAUwm3DHMfcsgYmK6dHuCr3
PwHuAK31/qKJEmLQNHXyVciYJFNaYCx9YV0KnoKifEJSf3mu+dN3rzBMu4IF
zCZeyToxeh9M9Z1AOe/nHSRZRYTrQxjWDS0HpEqH256LM90qaNKvzW2i2BJM
HayujCIwIb9tMg8RqCGPk+qSy7woOmYG9wzgv4OusvVcxpGmw2TaeW3TaLYY
rLMdy7G9tsilY8NWlQGxQpGNn3Hyan8g4oii3gyj97eXHG4iwa0Diei40tQ5
7clLjYQrOTiKTji5oHOlEdK8+NVQ1TgNSGjvNAfk00PZOwGstepT/CzuLQC9
H78ymHQLvzhEdsB5N/FNJlFlDKV+Q9G+W3XNsr55zytf2eABkPnc2vRBaTmY
hTDf2S47wzwj5d0y2/yEwzNfRVMQvNzo6OZuSHU5tIKLF9gi0AqR98MPvO5a
xEcawc6Nff08wOGvBvSANznf45d3yhbrtR6CtXSrxTZqEn1va0NFId5p+87z
VGhMBByWlk6KTKNIZJWPcMxJLnHFLYp13Mo2efPAxKce3Z0Er7HTfN/lOfSC
fwlROeY7hnWqwjVm5Xd2g58EEGL1GBuXUL7G2DhLhNSK6oAeRVYpALWcTUY1
cp9ZcyRdTUvSq3n2TSJN9Gj1vpJVaJVdNLJu1Krmetsz9HILQdi1JpwwS24n
fAVomdCOixJA/2bizE4jiOlp12OgTTvbnNfdhKC8tCjA7mb30UhwpzMIoduZ
yyWQn2eQJz62HypYYaHHLsUAGQwaa6aBg4j1cctan+l9ntSYy3x8hAscTTC4
d+D8RC5x7CbQnklQFQzgMswBY8zqY4aGwPeMR0fHoaWHiYq1vSY8OlNhl8ip
dfjIrYoLJKb2nj/zqBGJUxNXtwFrM+EH16lCBlRTtvuD/AUBDRVEdGG4tvop
IluvGi1F89EXV7QPx903Pnm36lNYsRxW4m72t//l5dBJXbuchtpayJm4XFwk
8glk2X6lK5VKDBu41Y45KG2cw2FJy9JwYs5tyHezadxhkbI+zDmxAVlcRMtj
vJMHzdAE0QZZVG2/JY1WX03LTHMXwxeEmeK885NANpJ8eKJDBW7d9e9VjdDZ
6LQzy34h1f/Wbio3KMCGhKqMVoqAQ/vbR/SpKo81cS21AbSUlC3U6nBfPs5r
rrs6JWUjuYLmrYlIkKE90BhHUvgcrzwzHzsQLis4Alzj0VnpUfiqN0zfAagi
3bcP5K7L3NHdSn3iuMu3yvbl2bf7IKocxuQggwjdJjduCUtZKCYbd+3qSdou
XatTuPOS6r1M5aDQJFnk1oxfZZv6KCpINaIykKde7BmkM1ZEoPJjLilDMuVD
mOT4a2IlObUffOogAe0yqBTv8QNquMW60qxI/LOux2heVBHVl7JdBGFmv1VK
J2fttK9HGLjlEaPkJ9S0MGW01KLa558cRwXdTsR3duaX2rE7C61DwPp5jABF
xlPjrZCHBF2iI3w7oHJjLRmS89WD4s0ijQwhSgxFl5Rr5tD267xC4t667sOa
PCFMGcaq1CpFTA9QZvwU2gwO/Ogih1roVy+4ACg1Stm0GiK473Bdiy9/5TlJ
+lPuKGBACOcMa+K/laslWtGprznhcgYWcw3pZqFZX7gbjOF97Dr9LhtKM9Lz
Gh/H3BZU+t+7SVjdx2EljhhIKsjomyMILXPMR148TL+hG1iI97a0U7gBiVGo
sOyt7uMaYx5n962C79Iur3wCQ5ne7s0PKNyF7F2gzDRHvKJxuVkUgurcRu9M
deJpy4GTSAg0BCk8Gt0m4Wmixe+qAFVBFOT7zlkWxvqLnRDDwQWyWeJF5bQh
3OoSy8BQ7ytCBsnDyDWvbgtsRVJsL66my5pLZjBMFFm0oKmJLFUNdMMY0ojI
z4B4OHPZ48Q0wMMN+81celJuQ9DqDpLr1x7HyjtV0Mni+D5GmzAjHxdeO3K9
ws8s8Q4L+m92FSop3PQdOjshMfPccs4NN8lI/+kf0zgtQhgJ6i9Uie8fsQT0
Z3M/dYkMjz8sjXQRrUkgsTKCpNWWK+H7qUOoW6ZY5K3a3pImn5a6BdZI1gAu
IqsC73E6B7XvYPVcVl957W0xOWAaSNKRR09TF+pB+JJLrq6iODrctAwjOkXy
PiB1IcvR59aePjyYxTpj9cwGYUa2SqqjSiCMKOoOPD+/Y53QiCw7jqMvCZcO
xmdqfpLqLR4OihWq3KdhqDGJgWJLQX5XISOmOqi+O56vxWiPzTnGgTYGGGwA
kqnJOsr1kGh2H7mF/xOcYUZeYNdGKFmH6Iqk07/SH4ihdao3HOB3ggz77l0P
53y7RfN5qGIMtRv6pWEMVVxBR1kZcU13rL3r7xyBnXmQ48yFN5AdYYOLm/PH
hO7SMhdamYVyQKj8QBTcYujBlZksFTgiXsEr8rZRsYDd7U7L1XuuxFv5D1XE
xUqAJticoSXHnMOapOE37D/WA9tQ5vsKgmaQOGP5ZDZFFkV+UJ6MiR96aywH
6wdNFjjtcd2KuXA61VDuA2/d8InYyKm1MFWj3a43WT9yBooqBGUunm6kEBOZ
Bn0LeWih+85dy4ohe1PpF+pdMdbciROZykGML2mk6ZYJnFedj8JYgHrTu0Pk
ymCBSu+h4u+aT7hjG9QbCYWCiv8oxPhBnyjrrnnICGjIVwY42y181Lk3RgBY
eo/SWzvxbJQpqCBd6w/hSSLQ3Z92N00qKPWhwNaHWCdN12LrTm4E2zNzXE/0
ry/jJjCnGFPXG2w9rDsG42N9WwR/YgBeR3DwqFxQk4WpveYRPv5wkuPKVQZi
Ay+HpIc0BHriES3A2jFGxQ2wOkwJhL7PCF7ki6iQM+SOg2emcuMg2XNUiX2f
ksT34Hpsjztwm13EGojlyZGhM5qLqxO6eqaivzaX3ZKhLLip1mdJ7zV087ZW
zisVpTMdjQd/qsaoyrdybRb4r7SnoFqaitk8SEyO1wSgaiFaNj30SdLibiXH
7dxtOr3e1pVONUeGnfbO3nJ7w0ufLJ4NI1pEQh1cmNdTJ+x27vissGcM0jEO
zRhVMu0+fNuGiF3INMQJIvZ+VjOGCsBznHT9bQFddeSfU9er+xFSFLUxK+Ag
0tsmBP8UcgJfwu7S/GVLuhr1OV6GDon1NTlTghjPkM3TAZP8cD/9kxVmH7LI
2FdctHL6nnSZwxbYG1Lj1WXJLs9Hh7D0pgjSOt+zA0Y7d09Cl2rzBTyAUu+t
ci8N92W3/BP2OOWWbAdm31RhYGJSgSvZabYcG5yYCCfRDndAf4YS3LwwOB55
9tXQCDYkZvsHAwhDhwLUjA3LmEsxgwnE/NIbInmJH+mBJIPricwaTCKCfz9U
AeojAel5Kxz0HB+4Xm/wYgbk0aZFAdgNgsPSB2rpSWbdI2O2jeHQ1svuEwx0
l4NlVqeuffUoVNzOa1GtrfOdgB0g2QOhuqTGFKiS+j28Oa4kPphFd2B9+yDb
qsfkuFXV+6oD+CFF6ioZB2QE9qgVkDuNTHMAebSwDtdeUs3RZF0aT1kocv7E
NlYbeXVmq3k41FqGg+blUiAlVk9iI77+CZ+nkbvL4C3KWRgtRB1jerW1G48F
9W0Up6dpPGH7+K9e0L1cFxLqD97d473ypZRnVF8yTMEAHbdnqdfqKlvawAcb
qOfz3bpl6rjogqqtdcxj2Bl1UDHxHgJpTJov60KnjyZqf2ozb1GfVljhXnky
z1S7yI3E1znNGFqzju241x/qPC9XFwbMrn3Nj1BRzbwZsA9gcEHJiQd2BbDg
+AA/Vqy7mQFSQ+SihD7kTCg7QkruVHvr3DlFB81Aeg2+2XvEH/hfar5PhcTb
7XJ9WyPm9smvy4mken7/5goZo4ixvWJ0+yXj2f0INjVeKiBseHqWZBipry1+
VWQXTYJ4pAH3ddR/CxaplSeHE3udSp0YAZJEUOxysZGPIXvR07KY0MX4ZJrH
rCvk97aDqRDjr+WdGCmHyiVA0y9HvFFUy+2rI1TSS7skABL0XLQZzNJ3nAXx
4BlnpenVkULLx7fVAnwfeeAPplqgDOoGs58hH96pbpMkHxDZvrNFWfj206E6
Ki+U35O1ilmf5KFdfliv/f9pO10jonUWCfaeDob2twGqj0RLDn6/64ApFf9u
1SLcpRIc1YMgkjbs+GVM/N0MWHg9B6R1rC7MDbaDyofCjOnjYpEoFC+zD0U0
YXwlRWQ3rQgy3ygCw6GHPRiR7Y1lYWz2gTrPj2GmKl9mttT5Y5SB9V38pzlY
6pTSDw/2Ad25/pyF4Cb503oOXcEMJ8Zjcei1VJW94s1gm3CxgtRbX8UKykda
rgWLbw2fdQjw8zbKhNNn0HYW7Iq5VhZxxAxQe1OKf9lotu4rw81XunQzlktM
Lf2pIGBGxvXkKGIEuF9x+Zqy8okdAzfI0KJK9ZHB3MnZTp6+Q3kcS29kd1K6
2HryhebYJOHq4gRG8gHHchT98zukeyb2N1qqedTc25bM4c/QF6CO5ZZPSUX3
1pIkyfFLB1jinlXhDz/BJvLM6U7TAKZfRdg76DqpqdoiTqzEqw4xE7kFHCe1
hSFb6vjD2WVVEsuRrpt25FsMGi1DIA5mrOqZ5Q40O04sUzGDRJ7LXh0obJN8
zZl7UonqZQBmGs2bNQq6Uw5w9AK4j6EJ3RMzb5Wf14LfDSPg8mBxGwUiBo0G
5Var9GVGgu6GsV/2C09i9PS73iOluBN9Zg0OSi6Es0KZHH3qzSWt1yqMIJ3Q
Z5O0ZtLJrDi8nBW5X2HmXbLVsEbj/SgLyNsWm8cnpIrJ3BwJ/gOLbnCPKpul
8GASwQ3pe3mJLCPieX9eENWinmd1zX3C3FCENJ514EWc19Cg6fwhB7/MKG5D
lN3xgYDwdh0WBo8bcvZq0PcXJ9VDfpGHozwq2I+vGEQwZTdJNrzCLxQJ80/P
/tTH0ZtUasFx8X9NSkybfLGoo1P8RW33FmD8gnnj9M4J7a/q/EDUbz/whHqR
rmuHMZdS4K4yuRlGv+T9yM1/aNGyalZHlyrSuYLJfpt1frhbes6rcs1O0ipB
yT7xVxhg+pwa+EmeU6S5dbewFoDIWqwWVlIM2JkVCjOIFZtpD6NKwPh1eBko
GGd47sENpPFV2pjqq0GmnxtyfZvFlHUrNDuX5PiDbYFnpBkaMV734HtdGv+6
i/xi2kXxfN3osUcdY+0VwtrlmlPlimEvHFSg6QcWhlXHBUiHZQH9wBscxYLs
hY14Qo7ckC/LiY2jEum7LFBUUWeHmtceKmLnsMPNr1wtt67X/vZkoTWfd88n
8pmRwai9ccJiEpNany0V10RPfnrpHIffP6L6MRgHFiFSVy9fc0J7dGEGu7La
H31lrR9D59hVICjGyqUDTfiDt8oGxRLWlqKudF7wQWBjDz39EjiW4dDSLjQc
qWr5vVaj0Kj1oHrWAt3endYHUEafREN9rsn4WRFROlv86AT0KWgzUIGUvRmU
lBHty0qaeTo/JLoxd5FRHJ0pi+irHebBz1Pf5LrII5538lTRJ1UQ2KjO3/cj
JR1k+W4dL6VMvoV7+000702zqORXUpOBIne1J1vbZouEUeLstwt1LMXxp6qs
AHUReG5VWF7QhuCcJGlxF6d4CkNhgfYc/E9LTBoVf5ccHUbhr9E0CPZ/SVpA
lt6cW9Pus7WA5uknhbpszLJRheqNjYXSDAWvVQMxTfjeV1GMA6cP7OOqiSA3
pZf8RcftRfGE0cZ/fbJFDHyGNF55SpV4Ju/OAUy2P9G0SzUOztcU4qaK2B7X
wryZj2cZdvb4LbuYFl12xmL/z7myUVkO9I53BDKMD9U/T9BDSxGpbhmFEF2v
Lb1gxtKuphSnft3A3wZ3xNaheJ3rN7ME9mxldCe4aZU+zDRpX7LpeHxhI9U6
m53UYkeKdXufJy8jcpL8WnGW51WYfJoQXGOKoLo/TE8piq1Pb2vCftBFGEvk
gweJuCx8hALtlq9VgGBuDckWEPLyF7xIfdsOjWu6BYFu6SCi3RIP6SkSPEzN
LsEVD9lu1U5epZlcpBbLdJQOemK6TOfHGSqxiLEA5/NZBSBYIcgzd5cT4wdi
RZTSqO7dQ4en0JJOvIKb9fnuICJs4S0MmIURr59MNzxttmwhfY5kMVOwXTDu
wizZM7pQbkIG1+6m1rEKOoa4BjamOyBZN5Vj89g90rgz+MNjxSpQhqghTAzY
YXrHw6nnxNuH1g/E+Z+fM4laeB3OCYrT5yWifuYCzxJeqtg2mqAOJ3By/XUN
88i6ODQAp6aQcTiPfd1mPE7prnNyJpk8XEKQvWlKOhzTLg9gpI/TEhndWEmR
/Djs2qJ20onAdhulwZSko6eE2CRLr/dyR58vpI2qo2tSQYW3WZQtFIrvwG2s
tWZk+ZLI0qhEQd+OOv5ysuCJYF9UL3BIFNdPCiTSBTb7I7pxrjwwcTEgr/Xh
ajEohfURa0B0ReuEl3yIOQfadyBpAfqiS6CGkfHFcihauCk11t6qg56okfXR
6Szjh4XQPk8NENA6VqzwdoRjlKOTISTQVQ05wckejw5jDoamQ14Ucs83Bfyv
/jfuJZ3KTTrtt+Linq/gEVnSAMoUixUWSh2a0i+yFFNyQqjSOSUtwkakw7ZH
GEKrZa5/28RLGqMOKEljxbXcRR96u+HQe8KDvbbRYhWlYM7pGLvjll1NMENx
8wJG+xXnT/V4BqhQEjnyXMw92b5TG6seKqw+dy8rTJF5G8/T8QPj2LhdaoY4
1Jtsqnq72TZq7aayvd5aB1xlDkH2D5gYg0c8D4Xm8tNhPkyXiYyXgtueGmfE
EfJztl4IOwtYd9YJ8ua7sEp06oFdeHjbxRp4XDhkufFHiO+Gtb8md0lef3tl
tiDwTCajN19ivu/6eRKOP+Cylftjc/QvmJI04d/sx7wL6f2DM3VIXBTdB6rf
pqBmXdxAwyJjIgZ+kOaZrmNcfhx/wquCVIEHtntbm2V0U8Tjk+6ENk5N0e8b
IxzOXaYKEF1hso1sRH/mH2iuhDX3Eev4oeMDaQmcJDj19KEZuGgHW8oO3mjB
RZl2jLeCm1+4t2VIPJybIHX8besUA5n82CslVOnbWlCpqiz8qp1xztPXqknt
IhEx/nEJB5mrnuzUL8if9sbu7qxhNkI/zKkTwf2Q1vdYjkIDv8cwusPE0JW6
aCqz35q33Y0GarUEvZX+z1EdIXjGEAKY0zuYlOa4EQRsxQLBLEq8xHYRRMIj
W7DqV47FBGOwGRPhea/sHF+nJQ62mGg7UVfc5AmLzwxuPcM0knmJ2uQZ5faY
minOHI7QA+kA9Q+TPEQ+ylV8j3liF97eZ2AlhqOZerpTZs7CA4+fLhE9A6Gg
kiAczKISgf6q37pKhxh1cHJgVL/qADEB9onWZq9vHwV59uimUryOytVs7a2w
XZJtaYjL50XROmDSucdb3POur3Ab9iWsof+mFiqTxzTZ9PoW+yUy5FUKvvyp
l5oGumsgj2ggamxst1CgL+adTfii45HFe3ub2CcScw6eGF2wUsn26cYdQeBx
nkiDwVNUFcV2EMfHjE8H5CzcRYPYY4RWu7VXMg5o23F9l6kq7BYSiYMJmbin
MaejWjcOH6n40j4iAU6j5YQukw17YkH37hlrw7tmDOJBxwJFHj7Cq/pS5CoX
fXRPXTnp48W+eJ9hwKSV7El4XAZe4N2jSv1joI3JuiSlGB3wNqlmhSOcvhPi
PX2yPSCmr0eI63GAdlOy1uvfKpHVK67oxodLB9EHIN6/Mk/H5QiWuynDIbfj
H8ADhGUXmTXkTgQbv/qP7o3F5Y2PC6YvwBk/jkHMoz7q3ctLgmkuzizZH9ZV
Kn1GERJY09CDP4F733p7nwtvNK58Y1wy0Prv3uoQEQoYaOz9dGj1hpvJ/M5H
I+MUkIHkt/0f7WhAkBRTFiBPVrBojmzShmfe/REkyb5pZPbh8lLuXVqNtpRZ
u5uWgzPGA8KSIfipo+g7BzbRa7f2PoEbBW6uArHFkeq3IFIlu7t7V6joMQWr
N4Wx+rMngkaqfsJbT7JuKjjIAyMX/9YhrOok7cMlmxvAi7geUuoS4EbgNNUJ
STiPzeH70Vpkwgzf9d608HlzG/8VIGxXo4lN9bO3b7nAz49wWo+ykwrVSzrB
N8JU4a85m2KHf6QPiQwi0TlrO0HR6H45XRzc20IofLOO84zmNaeMa+UZA4wr
Pqn3i5oXt7WdyFF7yxEgML3pMXu0IHVOjyKDeUlPpeoYHe4L4rSliKpvxUZQ
PmsTlxz6krmzfEfu00eandtyDRrmQCATCdAjbqE5e1+DpiQeQ76F7p3XgYu+
G5Y2F3whrzCfUrS7NP1RCVCTILBlsUluZk0L/l79iyRvO+NtPyBeN6+olj+m
3DC4LBxDfv0ltMxzlnkTRoTNfmRmQxH56ct33hD/a0f5lrQNpUHyO16lfNdV
7FJ69KQCgLoSvqHsvGIwyUma585Oh2m7XVoZAD1mNpS0oVGYqirHXj1FRsGH
LCMybwYCuzEy/p5VXLGqOrbh/0LLPL1rYw9fGmgMI+hCWc1Jes4ByjI3PDJx
gMO+7QakeLrND34C1EJyPhaai8JHcarURbeb//BB4jPscKR1LBZUWTANgMIM
uOP3m9Ayf+CUYHgWBHk++XDDQH4Kp1t1anmQ4iK/C+JL3U3g8Vs1KLHiPxNH
BW0KAVHs080TDPC0PN+ni7wG5XfRQBLuQX5UUJTV77UmPFET6ZAFoF3drR1H
ObklVSz6+t7K0XNhQguYD/gch3wMFGqsdc6+BGAnA7/BcpR/vsys18KbII4N
xuEoh9M1JnAHOCvctpIMlamuzyXx4v7EQ346MIhqbAiqzFvPpqjIglrPDOtO
K3CWgGRfYxZDeKJOxajYdfXstpqYoUTWh4sVksWbalb/S5xY3dKc/BmmJ3f+
vcKP1dfSXY2oClFzAQp6o68DpW3kg+7xhPf6k7G5qY/UTyWvsDIvECI/7VAH
mPHWCzF7tcoMxdMjDNletFaIc1kKXtPuepZW1R+0BgMaWgvfUKPCXtgsf7JG
pxJDAUjBxEN80vPvNuoaYJP416kprTVRgpc1JM0izLxgeAGg3m48jql6XG7Z
d0cznBHHbG7X/GhPY2HmrlDNmGtWXts5wzBswXMe4makP20pKaScqnaMvCzF
a16jv78pm+HYRYZEz5YDkGTVaV9gnFKV2qTJXGN/bdCF0E0Ztn93WS3mm2w0
Zvidl+GaNY515kAOk9+tFir9q4UgPezyzNnnTZoSRpIG/uUdzynNnCwaagAC
n3HOMY4Ds1OW0gbqhsJUU/C1tl6quB+soxRvNDM7WJ+BLh7bv2mSKHEV7pZo
qGaJJeGhXcW36JvT0yp49trR8IJBzUMpKsP/TLQo4pTP3SO1kODyGMP8KRCl
6EOwIU7UMOtPwyjESCV2xzKYp8FwzyKRmNZvZ3hRMGHEzDMtfLsdnt0sLYGd
QhANhtIL1/sSH/n65DgcTXjOhGJ2wOZKtyQ33qrs2uOXBt3QWvnycogzl4qA
w/5/NQ1y0XNZvHP6P2AssbqGE1zPXJK7ECwdO7l1RrE6NP/MBeEXhv0h1cHR
8zVeb5YhhbJwoG434UfknzB7MiQbSW3ihtgit2DC5iLN2fFFWYuCsE5Rjc/6
zR4twaJBqwnTP6Ak9On71QX++D3tg3Ll9qZhA2365wb0CBCSBl4vwjQbepT+
Y2ZmwrCgTJg6kW94cHkUBJKUaL4B1hb5znvkmYTL12hg+g5uqr6NKV1fUeUU
F7q3BDtdYzYMlg3Nqt75Zcs5Spbo50L9Zp0jWjKDdQM24zYTBJG0KQnB51EV
YRB5U8dSlEiUtMAt2fCYvXi7ruXUNJtMbeVBHzBWfDj7s2qjhqS8Lh0ig+8s
tJRqDebGvAH/TLUsM05dKfr2Tz2Du3Y6unbADDSl0Ev64vi7Xg46cG4kWYl9
YA+VZz8ESKXZcPx0NzceWFLQzlPICSJyQolcVRUhjEoNql5kEidUumGTq6EQ
qOU7quWesfZ90dvdof2tU0vHA9Q4Z++wathXriM/rzj4BLfhWoFR0y5YnfbQ
ZAo3nXT7Cn7nU42XzzNzVc9gFVXzocMJTSlQacrRk4CTu8O5ii/kvPenpo7L
hWGpE/2dkLdS+DqaJg2ByxJz5+wVxxDxVI0kf0dvtqrABERDuiOWLmYPE4rA
bI6GdsJh1awo85/BTK1jt4T75tZNmrZC8F8MMOv+s1DcwcHfpffVlaVoHDT4
EoIEBDjkiqPljnHmxFp0FTzv2fN+SoIplxJqQHI1G2n+u4ApNMHK66b4Aiu1
rQgFgMhYrXTTpA9x21P4FJXfx6cP3nex8utgJdA6X6nt5A5gRlSCleEFmC8t
Qzam3tM1KTJt0+YHdYl2Z7SiLJIO2Sv/G6SasiBAa+HhbSBTuBBH02XRiJ+k
5CPFaq/z0INXqyhzbGGwZ7Z2HOiblaGAAmZ6dphTOHEu6OAmOO5WpkbyxuDR
QhwDHWn2u0dVWVz/63Xs/kjpbeDaKygdZIeChOT4OeaSwRnuKWMuaiiH58r8
swXMsBr9b0JkZHj7QyZN5b67VVUgNYeRlfAGDaq1ITLzGfGfklR/81q+kZ+V
HLHaV7fyVzx2xfvaIV6383BmTHn2jOKubjMfELrr1aJrkpVf6H6Q9yP37c63
ACkvcgaPXXDtgaMyUIn/biorsZv7W0F33XGBz6wYmFFlRAWHMB+aubh50TRb
sdMTa+IV/7AaaTvuywrptn4ml5dzhkpmvuUBA0TzZ3n5bgvrwAOtN/0cKCQB
L7o7kyOJ+Dh7hzuBi+s72/3VAOj5y5Qdpdv60I/kcNFQU42Z0Av87F8g2z1r
u8pnuf0PjZWTV9/awv8rhM0R/CNxU/SVMHyzKO+6HWbSEAHhGrUojvEIJm4I
kJFFZwvEDcPeeUDHo0fgjotK9ZofNrvHdpJu8d4YLOR/5Ldkk+aviWDKzCRM
F3n08MJqSU/+GmzsizF0mih6R8b5JSjn633F3rI4E9zpg2pZLqCyCYlYoHa2
bbuXSj62+oD8SXqNT5y1NgfefIijQHU3Y49orfPNGfrWh2naZ5aEl7NgwBiG
lgQFPssqzK0Gpc5FAIOfFuQZpLtVaEJrfdtfF8BEBotvBNX+raZh37eV3izK
BcD9sHGXNTbPdGDisyy/A3KCzqaeldIuN4ZRYtEMkfacuqdaF1C0MwfGQWR+
YNQprOPo/xggucNquQPDnfBg1pGIF5MVz0L0Dm+ZEp+nEhPUw1RmkyAs8gsY
h9c1nEKPwN+2QGswAw456JV66eU5QGlwFEAjak2wuAyCdRuT0Elp9R/P3lvg
ZSHuMR6KtKv/b1umKwwBjPldu5T1bcVQDubn3oqb0zH9dji7DNH4b8HsNJ5D
SiONLbzPFXUgvNQIOAdSDkDt61iM0XViBOruATJZ7UjzM1q5tJaqxTC9IH14
qN1ILqVDNq1cdoEDo2i2dTFD0Fc1xrYVKoxaobSaJsmlnSS0bi8abcgIHhn1
xtHzXWU5vuqtumqGJzuc4iW1W5lG2YF7IcDwWT2VrOrHPgu//kSIR/IN3Ue6
+a3Wt5w+TDKHmFXcnMMbKDkVCbaf4mhEsXPfEPmv1uCxrmsq8Z1olEQxvBrD
LpgNXRITgFLS6F01dnmX5jKCSUuU6sXSkPtKBDPpYLaHMTRVHW/hyaXmAjIl
elAK5hGs83xG90VxWIUnD3W2lEX8Dg368VGKSyQEC3C0F0q/2BxOrIlpYbbb
Hjet9sf0aMxzqpMtEGj74RrDKmihuablnq3ae3zphmdQoglKiPSlpU1VM/zJ
Oktp1dPony7fOQVufnKs8DPSb34FQt1uwdvLzdgEEX1yA1dn2XFyDlCj6wez
jONYJaUgKVh2GeitetMqdIDr5wWJKTibHwSw+ptSRQEi+2t2n7hybYEpb26Z
cX3/yBZmHbGXKPNfcPA8Gtera5yPkgujt0cQ54NPSu37M1OMewldJ67lXSZj
2zmw9sBiJvrDH6GtBHgcEPpvCViucI0W+57wj1rTeMNwkzrsi22LuaCtuKmt
iT2NduDA2LIioNtglZ3A2CYU5EVUwrxiOreY083lJ+4fOO616oeq9J0NJFvz
y3kWy793VLvdJ2K/wvYF098L1Kn96NcUALGC+QL4oHIes67BS9VwX0dOsRHR
ridpFlEQmuWMyV5ongw0JEPQfY9Ve1xeX8w2NlCkBzRyvaPa88kJTC3YVbhI
++Gt02NaXqNZxPUNmm8dcNizhgxgumpoFSO722rRLy2/dpXkjyjyzbHhkNFa
+h0k8gFUvFNwIkSQH7Z47Zm/Xn6uQojBELm8x09CGYY/IJ1frOIi7XDATbZW
Jp7b51HZVJS0IpBvRD9YQrfrnhp+29OlLCmvNmbjuCKDit1jQFFfthE5gqOI
nKyh9SztXqUx8K+yK1n6G1c9GjFAFuDfrnuaSW1wVZTHwnqSqKEn7b5AQhhX
w80qlCGo7RY/VhCsq3aDDB9k0g6+A9cu65LClBfTj7n7Z0iiV0vHSHmGOSDD
cqZr3F3dcRXj0rtbjblznupwSeEg7NLxAavT4bGdnmRGrNzAMkFVzhied8AU
2eueltgIyBYeWiRBACNMYVNwYFXRDTDYDM2rVLOTVmsnlbEFEvgTQZbKcnHy
PxFYg5HKY6xZFsoqJkiEd2IgN++pZBLB/7nZWmNQrR89LOp8kaWGmMzPQMGI
0Xpqo2egCq1uiz3KqYkMLrBR2uAbwNHW60Knp2b400tbsLoJQwNJ0r0RDT5a
nO94FLw8iaU2nz/RxJ/xjjpU5m/BtWknLynHZA32KiAuxzQ2w07mBO8uqHpW
ye9TIWBOhB6ZF70Ff29grytSEzTJDCSwhFxQOWAucTfvPl9HSZsnZ4M+4MXw
iRjPAXn4Payk4RUHGnppmbTHOATEva3QOr4oDkhZKAzhJlxsnLBlfc/tUE4M
4KdH/idxEwSHwrIdr6m3bbZjv1AJlDYTHschOhz+8optgLKDXUv9BXeHRb3W
rxWUgqqBMw7b9gE66Yp4IryiB3uhyKnykvqz1J8c8TuBHPEYZfHZdtMoV8Zx
uU8gNNbDLLMcjZMtSwf8snXXem1l36ZR0U3bdc+sTIaFrDhifrvTcmNnXi1Y
h0PQde92dyGM1N7DtcyIuZEWgQ1MvQ1wukl9bxypbTjRwdgz07JLdLFijKA8
MJ8vKYcc5XL/fnDsXRKDa7oVLbhN3L+iPUvIeEMyeFwMm4q7EvSkQLnCEXy7
/GuyFrzPhxUNbAw0D68HFhGqhVHobV5h0YkO8S4ntLfgYttBs/WSQ5iGg8Ob
/rs0av4Un0BqjJl2Z8zesg2dypq/Dt0mnF2oAo+Ly4scZihp0OdG6G2sgbRb
j/ghZd+eXbr9jqSLWz69P7jq4CMPD52iZhRCtKqjT7r73CQ/7xnbkSpauHcZ
7qMJE8L7QC0qXkFfj0foAKLbLrysu9HCw+xfu8xfOok7bUpMwtcSfLcyu9b0
dsz+aV2abW8jTLy2hxV5d4yiB9v0XCkAiagaXQJIfYdYRYgaYl3dDq4WiHwf
ds63BEpEKU7MxS1Nw0hzfqG076ZHWNiCGEL1aeVODAAvpYkBNSyrPHuXf5BR
V6rxMO3+tAmfIftyZyhB7A9KMM30QTEKU1etG3c1BSayb+ZZB4UJ/3XrTko6
tyUKcC4tFkKEEa2r

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3FANQ23RCmB3SnOBuBKiakIDd3gamK0JBHXkoeUHvnNhCaGEGstdUd9sWtOW8pBYKOsXWB09rNhcwnzqUWDkX3df6zyhbOmzh9NYqyAQuFEkYtpMT3IOSsGrkwr3/69EBxdo+W8ZRrmig1uvseQk6tQEgWrtJNdpevRNLj314dAm0U2Rhm5y7qXpI0ADDl4gBInAqmdytpMKfobfcFbmt3HkIsuBIO+WPaQOtqcyNDzNzGLLK142optftrds/Q7Th3dSe3lvlX45W4zGqe+inoI8+RGUlnMrRQmWRn5d6huNeQRCb88wP5EVXpCnytm9pE06qL8U/bxWqfnAdGDUOopCALxQxmKR1D1TNE6H1mUcWaPHksBYlpgasNWSRAeHpWjTnfgwyAoepwj+V5YjN+jkxt5Vk8VO5D3zf7P08BmQ8qsiXNC/fi+FQfSZxxq/efZnn48BMrW4OH9wxZjMFqf7Q0FRWGZPpfDQD9+yG4gMgdM6zfpzdC3sSnE1rRv/gU32WsUDUBmhfWlmRGFKhJOdlcx5GfsVhQZuzHvEixqOfVx/tsjUT8da5hrc+aSBx+qBSQPZjYC9Ttf8bO5CJiUB13pygqzN/LLiyu0HPhtr++SAEHuSL/ds/c2g4TUOrcHBS6bE2PoSsOLDGTAsdSt/FQJCuQUV4swbboyWJvrLjWqYAyynjJPlN9Im6Un6tTK+SRCOE4+3LVOkB4NBMa1PhrC5/AQ2NvD/Af7qqQD3o4RzJpn6HY7q9MW6OOu30ZainnW3jh+FQe7rAnC5Om/"
`endif