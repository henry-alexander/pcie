//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lKKfGgY4yOXYOtftOJpYi/15RRo9smpkLUXG2AyXzlRvzHKSlXGri7OGXH8J
E9AIHEtWyQ0FCBxUf9SfvWLVaoFhmkoyMIbjwrB/L8B0QNc9uSUnxGcOpSRH
JNHbNX5uq2cTSu8B0cW5+DjNjJSgBwk7ZqJ21ZRY+lZf9Y8HWu8Qj9pH02Yi
cXIDvFvcVqe4cDrOaZWwgyZLx4+OxD7VF1CV873enSMpPiw7nCTsUfQ1sW6m
0CXO9zYHB/7sOhR5Pb/Fb82Td0o4dN7PfoAzqDTKRybzfQGicyb6okLML+eU
a5U3l+FaP/5EkJhKffQHf0JKhCQz9V4oCCQVSmo6rQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L4IEVJLv75t3i6aK/wrdVjsnlDi8+pvhDVJZaiMRBELv/pnMZMTTuVxKmEm2
pNvZLqg7JBtAYqExTdz28L7soLpMwmI4Wcj+1K8B2uny/OFPxaQBopF/cHaY
5pJ4Kqo3MLIZFquzZjAFY4zLVVpaBnJgSToXtv7Kk8YanH/RlxZaryEx+IQk
ha1m+Mqgyfitri3OoP2Sd5kQjeSiua13yQ5ox73FmDlouhS5Vwvt7ucGM9e/
AWiSomJBHGq1hISQstc7HtA5MIY1GdctiOvowUqSyqesOGl3xCWsZj5H1mxN
g92Udy4BAAUE3JXHxWvMOvfEZpICQCWJPNWX4Rt7Ag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VKrpnAoYXmWWA++PvrcuW7C3CobluLCDZLXWOOOzpoYp87rZWJ1Hszks7DJy
aGMwD6WaKDOmvR+F958d30Qqdi6stWgYfddx6Z/sLaIGO+RjAnwLyFNSdGY4
2kKeuP/reMB4iBM6gXvaww5SSQLunjGangooQVpjDCbyKWor8ZsVv+Dbl/EI
yn5bPBvbVNyn5SL5scJ5fZR+elBGUR3RhCHFYnjz1MrlE4mbxQ6SbNe2EXFN
4ZBGpnFgyNHOybkF67koTuFYX8DqxNJQ6SUxwpepCNGA+4/MVKrYo9u80T/E
7/mSRO/NWNl2F9WHz1XjMVniNWJCzQzHzGc1becYmQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iN0UzQ9hgJ4ugeO8Tq6PNcs0H0hBFV7EiaJJwPaKpCLyJDZraYLlhAxpxn3/
vFIh80o6GcV1dbiEcVwcNE98rN3xt8hxPb5G/mBklc4B2723Z5Zjy4f3B8ST
VoClxdl3JtouON41AcD843olRPPGQLQwe7Ap4bayrPA1ssKFmN8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
FL3XOYmJFhsj8vZky0Xsj0RGpHLuLnzIGAzJaB8lTY9ZJRKmeHqYfVOFtltW
UsylcMEAbT9MsLCAK8r7y6CbjLtJSx6jHABX4eYIOAKdvJUZOowvJqXYemlL
hpsrEayY2cF1WiIo7aRyL2KNIhFdROUvOiRkPUN79O+z3TmCYtW8wkLLXUYz
WeoMS9R37ychOXoNnnP7bQXrJV8sZ0TykC++cqLz9jnAUkGKh6PzHtm2F0uS
0/wLoce3dqIBdp/D1Y+Kwo6f5TpLJe0AYPnLnWjwoIQ4uq1gKqhJaUrbVM3q
EIkHDnAcUN9QznYmdoJ5QCK6DJ9M5cjut5FDvSMDCJEcEB0hE0MKCoVn1FUI
sduCmVVrrg/nfZxEUHgpVFMp3A9sY2HxArHZ+jF5/WxB9E8/PNhS3BwVew9x
VAUsFF5GyTNel7AKb8XL4He/Ad4hTobZgMAZpLzqZeX3WogaFAdDKhkXlgz8
TTjtn/wAIc79rOnNOH/tsClHEhVTiLfp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
izgO+wGpO5KmZRBfsEVjladyYUfMFsQWswsXK63yqm+SCEoW6yZtK+JHpEC0
k0d1Z0Khzg5D/FpIcbC44RyukQOTYhJEOUGGOMZG3c8jQrZzyf4373iUH25c
hMFnEJZNP8VnWvv8FiTAvhGrhn2OtdyNzpKhoVjEltzWkcomlvw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aRg65U6Nj2DmcgWK3mebBm1PNjpR6cK7sOfHftTzx5baOWGhgyUCm64rb2Su
nUkqM6O9NLQzJKxxHT78sL31HAb3lIYX1T+8zCptafLSiW8UwzivuldZ6Pa5
XSNdkKXZHVQ9zpYOg3An87+NszEtDtC71gqY+N7jeNKlW+YIMcs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4912)
`pragma protect data_block
nuecANJ3pqu9dxyHDuzkIhFQcZg3MwumlsHkaCxyFI32gfwvEe8s0h8IrClR
cs+ctH+7TWJqAhFGaEuSixYZhcdaUlXcgHV8eT3ICGYt411VgHE4ghT7GeHd
EuWoy9Z7okElBYghdSL4tfzhMBfrCxMs4ugf8+RiSJ9Vll1cF89MjLoKnULV
0vvP5oHnXMXzwb7pFVdEe4Tv4qhUqXTGCqpGxQi5MA7k69K71MJ/xxuybYAD
1eFDsUA4XXD9iRH2kiSYISZuBGV+gT5ZYywjCwO9SKplDDYlK8ODts3RCENu
nJtTTQyLyvD8Rj6loqaIEx7v1BSyNw9jAXeYHLJNmKmrRuVWUHMMgmUzz5mg
f6mn4bhnkOwy+YOlxzwbdWCc7u61tmdWPIftaMKkFLk4pcp7mxyhqz9+z/fg
tBKdXEHr9GCy06BNr83/kM9MZEWIoLunLwZWKwrKNKbg/HC6ajRjMpa6GLwQ
wvB01+2RJNzyjvhQQ+rIjQUOnZslX2zyDkOedBi035hxWo7lfFmf8Aq1s61w
MIemTCdtyTIpH99hWpe0gLt+rYEp0WfF4FS321zi9Tvb3KqXZ+cdV96IdY8e
1V5z0XQQoyFYw2ibO+4w/lf+8PPtEyvINPLGeibehDfk/7iSOE+Cqjdp34O1
kYUl8l7/LE13Rq2SrK9qa1FCSk3JSIU40dYs4I8bI54Albp5j+vXVOIL1ZMZ
2go410QL+EAU/4rWnKiA4ZpHGKKOpCeR2SdOCNHkqjwD03DZNc4dLV/TTomd
eRoBvlMU8f1oW4CvgPsgFrvXJrI4DUNjX4QKgDCMUjt5YqgQ4Tssry/j/iF9
+P7vvkoh1IGJv1Z/HNvpZf3MMo4wiJ1ExT6PRDUuY5oRN3YMwD5Um15UiLsQ
RfVH/K8RWLe6xrb3a8/0z2Erq3Gz0/HhfFP/ZEwjvWtSeh3PVZ3btXtT13vM
0qkSwI/AeWtB2EisyTBBS0D4+JZT+g8T4eNUZ3q7/73em4VCXAP2Ibn2K6m5
2vuRo72Vh2Sn337V0tTgwE1GOLLVbhPxPxdnUb7jXrLyCs+XEIbD0T1Qc4wI
mM3VQFP4wHXiA2W7K6k+3midEJ5HuRAbPa+GgUkp5EBuQRcIYhqeZGlH3H1j
bCMYNFXYd2bnYzvFhiCLXRIi2J6d6PI2ZkpmWvAbeC1XHFHca3CDWE5dehQi
Ln1aWFUuRkYyEuCrTXnrS8jE7q01IR43IMzMMWchySQN8Xri9J+X6IenBaZ0
dGn1w4gjgtqF277COJaaoN9GDFK3PtsgMZZdFt987beNa2XALWu0UiSKOTwc
COuh1FEP1fO53SuGoyoEHEwwPTRlW3J46AhT2OZkTF/9F0TauOjnCpaSy3VE
oKTTeIXAKkCKJgJV54oTLBN2ry9/vfhdYRjjIRDDbvIwkfK8dVwdAM6NqPjM
zEQVF36xL+sHa8T5KEYiRCuLbek+vzz0qtPDzkqW+7cB/6M0hyO7vNh1+boI
hnb+woTloT4XKNPWfF8qGn483VvPikWSIVc2AmgkVQPjfEKw96MdnG9sLMKr
F0wG7PT0LQcVVZF3d//1ZG3se9NDUxr7WdFNXQh2qXZC9Rndc32K+wg2y5mi
GVYMGjEZ4yM3rds5Ih5fiUSDdHCpzTXRR9RiErk3Hihs6Ktr1QngZ31eWHP9
qPnYJc+4YT8MLJsN8q0dtt5TNZwwtS3fmLTZNUfrqEb4DaWlhfHlJ+npJ78I
xIyMShI/VwsuKDLrR4tVkSPVKF7M0wSz5K90ZFnMqAKHNsz0BC1mqXQSb/2x
16LQxyCMPDPMCI9e3EZay6LnYhsLWNTpeMyI81L9GdLfvP3+eujf8v30E4is
JUQf/ERiHq4/ZsamTsASHciylRWQPePVrJTCHvAVkGqMRcsTLHoGMjyZvkXj
5XS8oqOazz+ixmnNHApnlgy+BYHQD24KIbExmQVFP4Nj1viVIGmd6hJ7CsE2
c8uVhDJ17mhOhxKqov//zWqVkpSvuZLZpcmUQLs2AXd1N0O4DEIV5mpH8oKk
fsAAniJ8K8JZJHDhNkZtoTAYYH5YkN4Ypnh2RlGu269hmujP6CeiiR84zrM4
K996lrByOfCPZoNR0o0qgZOIoGza9lvCLN6K1XevaCi+23MXhj76TAMHpicE
uiRtbwMFY6fRYGyWNTfersfFQEF3mfguCbAKQoVq2oUkn2UWLZD/bvxIF9rh
PuT2qDs2uuZRTRq2XszJxEFQEpVQ2WU7/KqA+O4LlQiCzSnL4LAk5jtaVaB8
uzduQ6h2+1/XkWkHKUjv1Ce9Lg9VNnCe6hOUWvGHzvNth66XA4mRIYNx3Scd
E28IoPFpVA2w7taha5S2rOcxfPEvIcw0Uzfxlhw+uuHquMDjH864gOv+46gf
+tkRqTH9ETOCoGdhI02pJp44Zs6sIBRQlfzsFOoRjPKE/OhdEbOsFd8KNpEG
V6yxcoa/jUJjDGIZOpHJhMkV6+uTkzhnlb827Soz7pVfrIhAbDliaGjl0Pqt
A8PiNVKAzL6O8fENcJXK87CWpQadqRcRI4MuBcwhrzspiYkWo1CAwrUibXJw
a58LoBCJt3HwfIsym6k/9rgZgrA7idWqsZ75wqdtY7H/8n1IpHanY8DLNIPp
ijFq1OBCPykQ4f3u1hq/MSWrcFxVOjhb3hEkX5kcFrirHeIpiw0J/NlUR+y2
+VCFVVMdGZaWAgcZQSWcZRNLGuf4qDby0gyCajj1Uorzg34azoogcBCOzI84
i/5Sgs+Tq7qRHJu9INkvMGk4hetL7ORO/kdDEmRufuLx0VMK0mJa88Fg/iNF
KSCucP9SgSjLAnC4ChH9+0MGVCGIl050Z2bOCoCRH21SBeleV8/173khQ+uT
WZbXZHpbNP+0+aVOXwTk7mQic0enbG//0AroyNvG7szjcjVL1nYabmtap6eD
IeOakQeH4EyzFHadHNLeBI+l/PpdNevz2tsbo/Rkb8h2cAMVIVNCpoh4CIgE
XSGJRtTNxX4JOoNMHug4d3JAtzdDxaz5FvONyusP6uQrhCkr/72TCntHq/XE
h0GvlCR9FrFgteUnYMxIzuHnqC/gMo/pTYORmbHY45l8mjdjp01BWgRZMdDn
M5kXskJkGN2MV4+zsFwtQCO5P/no23L7MuKbGYSRwdq+wXbq+Wi/t7T3O08U
R7yn9mCNkQoEKK05L/KwKOXbrmT6xp76kvR/vb1UleuWyZFMqxKydDpI3vt/
qGzjN0qeQctsIa4awZ4cgdE0I+5ivJWTIeefTl4eF+9IN4YjippuDohqdGgm
tuiI31EjJUQ0bBN3wnpNprD0IpJNN4o6uMLcgth4weIpv2vCruoVBdlHQOfZ
+rrpN8Ds5X8gTbbqS+1tsArstgG6x9mf7avEle4JQ7lNuKGlBW27Us1zLymD
2yVABX+nWu6ttV3oxMgFir9ltu0Qao4+jT/4nwAnCvYRciPcay92hrTD1xFG
fHGdrUbbkiXiZCpgTuNrINFMLE493q/FfbWm39c3B5UuW2vJaoBBmje5ZO7a
3k3TXan79Exw3hUh/2mScw0cTi2kYM09pWXoQb1cT635b+J3QKX1fIiVMyKQ
eNf4L3NKv3Mk2C1n4FdX+LavWF+iZCVZ1Gr2PlooFn+c4kBiZeymIa/IFj/G
SOobwN+lmStKiiRL+h1f+r31mt64Fx71hkV+j9QqLPOsgPsM2fJBgtuTxq/6
f1mqkOzH6hbTVm54TPzWpPnzVr7FfJS0c8c0OLha4UvI+VqhIsXEIN+VBcvC
2shtrc/wzeviAKgVaNMURMNMsz7vKpqqANm3q+AwPaafeeJcx7xzca8/07eK
FaZxM/J08MHnBpDyAwWcLLd7rEwyZKWj9BDyGALEUo5p0Kq8LPhCMDatbNLP
MjK/eRrhCdW60pmINUJgpGx1k9cVV4cY+7af3jzjafyP45vIhMyJoo/+J4wn
o38Wb8P5I8GNiSEmkcrf2VbFYFtN5Whn844KheYg8RGRf9yLwPnBpbACngpT
zDyh7fRsqp1IwvVGOpF2WrQpn3GUV4liQmk9img9UVwaa3fxWBJe4yr1KFTs
HgDVYQEvbuV/fKTe3q6tSNWa7bULkTr9fm06VY0Oe/Z7qs7slv/rBm0rqrzM
70dH2qtb3P4voi5XD4zNPINjYOFvziDM5QijOopvAOyz/vqpXjSxUE5FcPwr
+/HghY2fCJg9Ub0t3hfNFYAlPXT5AJLCCVUt1cqpNz2lqy+RyEBouT3dG0Mx
5qYtz+ZUx+mT321TQ498cdg1ExVoWcmfsQNupzp4wjXzMSczbXTI48iZYezi
k4Ruc2sU7Zj0T0/1gWhozM9GIrACauSCgkRJ8Dxh7kCdIVSa7L1b/P+0ZWAb
KSkhqUo6njhHn4wGRaXPHyWFIOdhz8h0GTcb1ojxWhd5pGILmpU3dwOwIvlc
CPl1/AO9RII7WEq9g/y+yAk2S4FVvMla++kUE5jTj6F6JTheI6KTyf4vqidO
53oFILIFMWFOXbuwchoShVop+CICO+ep1RsaLorsbhR7wogmsCHNnweSnln8
3LZnqDDu4C1SriE5c55VOILnX17qILua/RFEpN/ZvYPUybomPYCk7x3JHW5P
XNGElLkjA03gSfAHo+FwX6X21PvzuGkyCiio1/juTbUFsI8IaUEUJMOlLme0
FPeLNPouUIOUpypnZ2u/wec6QqriyeBZcBxeOvY4Y78bVj2L1k3ZFCxD2Np4
AKcOqfyYj5D6y1NomwV3D284GwSZjetUxCfTpSE2Bf6hoNtsoYjgYn1gF+Ww
y0Mud0wQw+eHV5I5xHB8saLwIqlFSlXRyjvkXLpTsa9cQ3KVVZeJT5PPDHnH
SIZDbtG1ymp1pO0HdzApE7OnoZICU3t2ZnYAt7BY6sBPw2ZHl0jSr4EHkBUP
FiNVpph1e2M942zrleoClie0VMsUPaaf3PhjUKHTorwsP523rxDmJJ8tcuPF
ivLt6mnUxSzjefN+zuoZ79fS9Nud0y1sKtz1g1SISHPQ/gJ3MFZ7zIEXO7gS
7hDri1NvLWwqLgqmjSHLkzl/aFBCskOmWK3ZZhpqs04sHhNHSDeZYU4LgKz2
3UKVlgQb3eoQ8nqRTV+hTikmPDT63oJ8jmqBwFwpx0RrgNf9tx0LSLESAZbU
pdzeWGstkO6awIhZOL/ibBNTyFQCZQJQBxqmsgSzbVqki2E7JOZUHeVsqSze
Ppoh/qWOICMN7aeP99DncxWGl8tiYw7AG/0BLYBz3rL90DWxvb0/AgXPTqD5
tpNAAL4FS9QXNClDwvBnbVvB+nZkxJUmQD0aPZ7NIZnzwuP74yV4+UxyoZjp
WGdOTTIWFuwyTldgyWKuRrpRpWHvnqegTf5OwhEl7HtLc/9CYt5NWJ9V8NsX
6Aai6D0Dge+6FnsZ1iv+sZWUrTUSOFdfAv11SykoSTLtBqy412g3j69cbJfp
AfPc7/S70ZgHropGbf6j1GIPiCYrFIp122XOZMJhEBS3AnVQ7Qeat6YI5h14
EXLfBKtFqMqP4FVeUEygjABJsOynLrsfS5QzQzWgMTzPPK+Coe46SE8F1NjT
PGiStuLug6BVF3iOwSbTNH4t2nvU0RE22wQHhGIRHJ8pGT3dKQP+vNYgdxLG
0XH/7fWuA50WZnA6JCzbike5vHdT8vQvoVLPow4MUIUS9kLyMpGkBmXh7xHa
ieyo233B0W1JG8V9ulpx4CVp7wMr5BzB3eAh/6LFx7vEt0vFafTUF254xl0R
Ymn6NZhLxv6jgPPkudHvvjoOb5DBV63hxTKPhpcDEvJBDbWYCu5S8F+3+7dQ
+ZKPfjG37hc7DvF0iARnfK7mm+c8BDtKB7UskAy26cZOVGB5An4DaY2ZvR8r
tk1K6f4keV+doOeGY4c3w98YAEgmfqcyNwPxbS3gNfBa3kHFaZ2lbu9EsNtD
znX9fixqWdtIMf8YQOsAT7k++cnLw/jIEK4YbW6/NZ5QfvDbxGaUboB//5Q7
8rxvzldfuLEV8KxZlNd6a9qEERXsPrde6C8gPKIdiZEDi4oGn5Wi/v5ZDnk3
8XgaLzCmgw38J7yyYUIQPPnweFNyuD6QU2Bb2K6GFFWwLN5sg8rjHPw6zaY2
mh7b296YIswMPizIqcJM3QpyvInWjWbJ8OzyjjueJF6qz9Dh7aFGmIOXjsrP
b7XR0xSG5OMoJbCvgGPA2p5z0asu55n7nHCSaY7qBuHgzMMASviDuuGPxHNa
1NilSg6YyoYkiGysx8+Wrmey75vb+bpOcRMNbDFOI5qmV/RyY+LFkiIaty3m
DdoXvVcmWveoZtnENzAjn8YuQcm0nkRYhmT0kHaZTrPYR/w5J0o+dh425DQB
l2oTi2g93Wo+gcwtAD2rTuyjZg1QfOeGbMVHg9fq0NmspJ4HpqgxhqUIcHkA
gz940QDccBl1XsSTK1yBfCjYeaUFU9J87d0DJsF4zRL9KO6gZt9mpoL0ZTy8
43EJonWUZDZkz28MiqW5IPwhGUD80YPSmo8ddf6YgxgNTmJJVV251vM/ZcZB
nJimu0hQFQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mD/0oBULxCWhX25ufwJSbFDmqrStAdsTL4UIdE33Nes+2I7rOUb7Yoi4XXT1VhwTgheFBI6zaifd42X2FqppSonILu6EpAdhVaEYVDeZLbFVT1FRtxorGvcdDMB8l3uNFGUmr7QTALDTdOPG6yYrckZzPY5lpeKtGHDzjAx2hUS4ikrubsf3P4rKKk4URMGqa/lMwt3RqgACTMrUU9+SOtDGvZ55Vbyc8vxU2+6Ha7KRVQZH/XCaJ1VF1/t4a3uTa19RGHiVXS1JhXVeA5B47FGEbtGpSjELwXnfWKVS0nukh3qOdiiw4bz1zYOusr9oIt0OgRF8PdHtwgH6L6uXCbxcMWoGjLMFIRuT2e4PhAALN+hwu5OyBBZdsHVnszR4+rpbiE+k9Xe3U0JmcMkLrE0V/Ff45pjfbX2vT4vTHHGzNWpKDLiGeWNlXr2BURAD51shbU8G0RnJW2BVBXm1NBKRit86UtNZm7dNrglZOcNj4SN36e03qO8JUELfrzzUv2Ja6fui+TLT8K9bOKVnV+6HKXhh+ofvRMdGUWTu8A0f+mikXUk0S+qoJLrF9GbQuNjeztz/uztf9OTIAiKfo1q4zC0+bvfreCD4rkSrHhFZdq53bpePvtsVKk0Gzgqrz1LxZoK7hBytrLEMcFzOXsndyB/SWj5jF2RekhVfjN4C+w9ynTF8DDyhmlD2tRaXPwUPLR8fXfPQD9xH0sN8Bl/ttu04aD13R2zbnDi3qhw8JWkT5YJ2oa8yjkJ81gx+7rEmylbW50J/I7TW/hmKth"
`endif