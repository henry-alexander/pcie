// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lwKqbEOevppelEIgqB5byZvn+uPRl3B7zsYUI816p7500j54d9OQu9Z/XjL3
u1BkdVxtUoQZJbHmmO4PbJu0vVol65SPocFTH/LFz9l4KFhdWToYee15wAOc
6marnF38iLx2YsbGTyx+bliCIdAr1SWsLXWYwQxFwQ0vLL/E4Lh/6FrZxzGL
iP0OAMsNtK/4zLTq1UoCson0mNVbyq3BPDI8m/LmFodrF23Bms11SrMik99m
shwC+Y+4jwW51aIzpYZzMPuYc5w2HA2KsPAtzfgeSJKkFNequqI0U9z7KGAc
ZsZx8J94s6J3twugY+ZeirA7S40gGmHfxFr8csoL2A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
jA4BiRSjO0W9CSZSAzjNN9MIoJSlEZJHB2SB4D531HkAlyM5tWMcThUpYkJS
7UGVLvGY6zXvJP+0GD0Q9O1a/HjwxvBNdr1XsoGfUrkV7OIx1Ad6nwMkRsDt
EkHlIQBz/95iuUOwMSJVP3Vtk2KOi42hKPKQ3Q6S+O/JSMX6lNYR7Q9jTPTW
j3/0TOud5tJ8scrZaEIThnObTsAxyYXAG/XsbWDGiRHlMzwqBA1Kv9GHoEjy
uoEB6qfR206IYfj4ExKS3iDV3zkVt6iBb6mRhlcnR7Szq4T+mxIUTfd8m6nQ
wUbZBAXBqYAyHU1oqeJn7cbXeDLPIruzkMdEQD3Mkg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k9M5U8vibadQJ4HrnNnEeiF+lsh6GPAp9A2ICXzKIi0sPbZ7H0U5KHhd2AzO
HaC+bLHbSVpup3cd1CV+JlJy8rVi10Hz4X9/HM55m2sCXGgYzmCyfyo7Wq4+
TmDKTp7eW2qmmDDYUahzkJi4kK2sXQjs7Ys6vdttEqYhBMScnjHDqfCz0TSV
Do8dl2lCkUIOzegUw6RMgAMhOK73xQSOoR9xbKanWcHvc9vfFa6oaJs7gvMx
j2Xe87gTuBeDs+UzEBdgd2C4qP+69NEia/rqh2Z1zKAKYg+z/uiiIqgmxpP9
9a5GpMltjdWQ/hQOytO+PVcPFw7EieXq9Sif2DApmw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KYqiPIa5tSceed7fyl0MMtQp2qcQkuSvRs4PZqfdOtSSqzRzlE0ms0x0qnuj
QZzLd4N0IirCrnyTytiOsTHvBBoosGHJ2gS3zqDDmdJSU9hqZzgm60SzZkh6
Fxk4E9tr31xDo+w8ZI4Lz2hvGNfl22iCRwhlukscG0PkrVpdc5Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XD7JgF/ybHFARxRVJfkRrGumzV3xP94rwLV6mPvvOak7CqqdNSEnBHFr54yV
OMlWCE/exlfD/Rh0UOsDkgd4+H9yvCaSQl2U4HhGxgpoAWkDfnqbUzWlGLJN
qXfgj6Y4xL6UuijSgaTTdoMTZ6IgEFvgJi+VetZRPWdiaTr4/N0qxa+MrRBj
CxVaRcMWqJqhWGtn5gTouK7ZJWW/rHox60NjYcblmPYTHOiif56jaRlt4r77
JzdSRXnIBQnHYB8PGaSfYHGNiEIdOHHC5RyYaoSWS7FLxvWt0OkSycQ4mEKv
6Lmuv8kyPpQXrO8dF8HBvjf/BFZ1mL0Ytzia7C4aLLXkVoVUEDG9b7uy+67c
1J30Y69/uKxuZe11fZv0YwvL5qlMs0FR/GfoEaNPjjFe0Ism5jAlbvxM4Tuc
pcjEKgQLE/gkRMnW2b8MHw3LncgWknG2naKValFj1zgK2mYHQKgo+UgFX4hg
SWyUgErfg8NnF3iNhJRDBtUfvTakNhnm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UDWCKdJnZlFmmfrxH6KjowT2OU/8ASqxTgLCWVrp73DcJNvKDhdXGdK4QtgB
D8uuvfJYP+/7V3ISX/IQLkCigLEMb1Yi99CfwFQEvLOz16tnafSxBDH+D8Bu
V1SynKiKjXP7kFGiEzneOnhbpftVBqGQv/cpv38Yd3BNZx/EJ3A=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fP8WIPM3wScuFKHQcNF38FRhAJSEo2Jo/tpFOi5iPwdos7ZS6JjxMLUlhpWE
I50aDvsosz/obFxFLxTnfwcOY3girwkhdKnl5CcracMyYW63cvI9jAZx5CTA
PdiE2nYno/z6seV1w7WRnK+PB/rm6aFf7VitmcgL5qC63PsWpwM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2432)
`pragma protect data_block
N89qNqp7HCVf1Qp2TdS7Tqt4UeoPlA9/gfgFUvqx4nFb+WjTkjUf/Cedrx4F
xTWwaARBZsPW/cq6AAQ5hdUttwvxRnzKutDCj3+04ajYEXPaYM77FwX5FR7a
W7/KNVmc6m1PwKvHAhvewPnPtXyfID5VcJZ1u4Oz6Dyk5ike966UJQl9Mf0c
q5LBFDPjOg1CxhYkU7NKpKQYq/rrQnpRWUxliiSyKKBlEP6IOuaBuZknDJq8
v1RvQ4025W86nWvTzgrFxz/RNsrXg3SNSs8G9aDiW3fBfKKr7770uJdsnLzl
WsdMpr06N9buPxYIjaOQ/44CbuR7t57yQBl1Sg66ttEfmfZLjYP52hXzfBnz
9jvRMjwv9ZXVTpWANnD72Wlm5Vranxni7KK7g7l1wBcz3u92EQ+twfZ+wsTP
5KK1E7ord5rQmokfED/+wBemTSsOAHwmiIR3R/H/eUvYHekC3WsH+us+331t
Opr+gV0eyxyw5A+OcXUmh5zjjenT/KczWtkihM5uJWgdvNtQ0aHjCcnAnzYH
XvMRCeDjyRKHmpKKRI1OBBIN1/Fw7OHLLeIhRleoK47CPT181q6VQTtjidXt
1BaoxZqe1q1mL0cnEXv14Jnaqoay9VeQtZzVrk/YPRcdRtTDC472l546lFkH
AnbpIlGvzzRBKeCVfrFDclB8af7+p8dZPPooi9qg2zmqvJnyOWH/HRNQJ4Wc
iyjO78hDbgWeG8jVn5jAwZW0XE6SzYaEI34ef7oDhMd5z9XwDKsRy0Mglagf
haScRBqZtcY9jCL7PNspK1mKjnKacZFOeMRHu8RlUDTckD51bX+2tQaxzHrl
bCpgGVBPHCp6O5NNaaKw6Xvintz4BJ7xUHh5w/vi88FvQ8ekMGc2tHwGrURL
ufJ9M3j46oGMZ7s/YGXOUoneRkUJgASF0LmipXRYYTugEw3uuLPUFJG1sRd7
f7gQp1LTYuxLG8tjsMe/oFlbp37y5DCGc82DVkUARYG3tqU08Ppd7D6k1UJi
QfCYZzDoZGgnWiWHlUT5pd6YPVMv/m5it/Rj/3Acx9KrsjqoOUzqgnWuQmu5
/fX1RXWYJHwRAiEa5SlRl84/qzNpQorArClvsVZ3eQ2wn52Not8e2+ECKSp0
pSdJhWL62k1Jrw+tiZhaDZDNpg72M3jEKrFdjnzhpdJo8DhIzmidMmPbK61N
FdQN/uILa8vM/2RnXF4lsag+6aZ2vfPVheqM4a2asu442ilb4Osg22fzyBbI
VkP8mXa//vw51IEfiSeT6yXeZz+15LVfF3OfrLz3jsjmFwCqj98EBh8RPs71
yrU7EAkXDyMdDH6LVGdSweybBKc56CRnOul75iqKyJKu9P6w30HQ+e9+5357
RO6fgo3HoJwIQcu4HZMpL0ovN/inSS2vQE0cQHsuWwRGq0iDZmfjuhoMbNNK
V4UPZXi8ICUHunW9ARwynlIM+0+N5qSDYgE+0oJMtKIu7TJfw9+b9/L3PvDQ
rsCp9EsF3xTytO4kYNHcZ4StG09aQwDYb7oy4xdGmjQ+Bxe6tntYSk3KcxTT
SnE/QCiAG4NvAoDLho9DT0LDur+Em08/vGbLuQEcoNQHhmo1Gvn0ak8yOUr2
wuYwXhvPQfr5w3lgFR7rmtJerR4TkMsexs9ij4s/4AA5alSUemskbVkHKqtm
jTZFEEeDZn7dRWhYVYbcsN2kwR4A3WEFPAHTxv0AHXxIkitKyN04NE7J6Akz
pN0NVzDbKU9NOKv+dKgQgQqAvYaVKZfMoJ2vv1m/sjCfqYQAv1MYXR//p4wz
gX03vnBvyuYFqSD+udXF9uKTlWgQdvEiYGv7+B1Q5EmmHdMj8GJpn2BsFO6B
4BAHtTgyRrU3KNWeTZeKFiqjWTZvo2+zoyfsFpOy3jw5Nfa8T4B/EDq572c2
UjnqLfY6pUEPTarylERlaJ6rUxnuVwVQ1812uJCCdWM9iZrHzo/Ya+rt20vI
BBGbQcOEm64RxzdFeLyScwh3X/ldw4Ipjnxo7wVFNITyPdjY+3lVUqUJE2dt
ndMPi2RFgOGAHbdgYfCnzL6FIWXp04mmpliOuoD0JU9JOScFkQkxdeGTeFWY
RJTLWCesYpBbLq13UOuMqY/y0wVueZyTV4NPhW5Dd24sgED05SAwUR6eNFgM
OILKOCHb2BuU17s0dhFtshzZJ3Ht61kx6wCQX58Fn5l50HUVcTiralE15U1m
TVRvXkXta78XFQbttTetIbA80IfzlRAzp3OoTkDsbLAC7JDKYXHkGAoJuQ2I
arKZDCyV5qCVWV7o6k12ngJsWkEa+4yCIzhY9XBBtndUnjAtHcsnmeRPsL59
4n4xLsXwrOmk3FOpzx0IV036hdzPA2IPBk4UvY0wRakKeVLJkLeTjoHUfYp1
hK9JGm6X0I2LVxkrA3huTDFXkd7ARObBSXwKIPy7NfW2ZLkI0S1jW9qjeKuD
UDURuFas3CpKW2gg8fmiDOx50Uw5g5Kyhzf7qkrqmW0PSqHIwvcMe/U+aAwO
wZOe5ypvuPIA+k7SXV37l5VbNX+oWrbgO/TtkfBehLLH5rE5euUF6NWyT6as
9gAzxvRnjSIA0swkWkutBUD1vnaCjJ7TFWeMiXlV1V9aSfjzyQ0wjpCoMsg3
j1OhXP3WGCEJ/FiEavLVQv+M+/cL2g9a1pvNxAF5uWvtV1fMMrMLDIBX4D5t
CxSbwBAsXdr2MKJvkGwuvpq9JuLQ/jT4j1N/Ffpe0cghW2nOqOiZnmtjSl81
Jd6n57T8+waDLf9nuA28D0V0LDuNXRl6dSt6xpkul4kTmRxTE9pPao/AGEBe
q/ydXcROE7laAcy9vhazloIcLe5km1GMmY/6VkkAmCptjf/evwYR68pLHH/Q
L18IiNkRuu4ArQrIUWiI0zzIeUd5Pbqt7AvzA6RqjiqRcPrwlQFMVnnPMXY0
ua5AdfQt9mkP0gDbfBo/GZWq0XuTdEBmdcnNWGZMYvPg9hiyN47BMQnAXwZI
TucSBnHPOCPNt+kPLA81g0zF8MlFHgBwxbeOVqDxGc2456wB4uhYzY3DaR1k
YNIPPFif5y4e6m8ajMUBN1ihmDGKBANHx/uFMQmJNxb1VzwNT1osZo+Bkv6g
1fn1+5cn5l2kRm1go6g1Js2Qv3pTKTHKhYWrigLjO3b1v4f3jxnqaQSpjNaD
byYvoSJh/Ao/SKhjLHr0Jju2k+ftWIL+G8Ym24XJNLbI0UyIphWKDBNniRTc
Y7g=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q6yHuWkcVSxXILMxT03xxn4PZPg/QDPOnwuvv4Ls9+f7mbwHUHmgth4nXVYWZfrzflD/isMpTPpGmfifI0y25fGYx225HLtVdQvR57LoIvMRNyz9szYivVuRRVLOqEhgpofnoUgw6BfZUoxI0ZhrcOQbL3kMLx1fRBVV6mAe06QN0dZlQlxSgZFlX7prx0FDOSvlmROwGOgJi6FbpFyEqcWp7lEvf2WKY5ZnW3R0tqGuH1akUG+mjO6nkWt91PRXJlLyicURHiatz2oaHqH2S+x2tSMxmWvsXtnlOuVFa6Zaj30PgcZGBenPPCGNsI25QnbR6FJHJGGPK+A6gWL5HdqxbBPFiHH0e6LVs6TNEJ6KcMJURQBI5Gi1SlWP9k4K2IgmrxLUhV53N1d6eOTdXUlJq09a78gFShje7qFzP1QuQZJuf8hoOhQvXfb1eJuCS90zu4jvToh83FtwxrfSvAA1WFDfQRtUhKcpJ3b2krN6KE5yvgqNOoHWO76F58apcgYSZTFK8SLA2wdHd2PGTqcNTj7wIRW0mju9Yn7wOkG/LFAGJVKJmKyFp2+3+CAGcPfarUfedI5U5H+Eypg9OQ4cfTf46NIOpHBv61STtADlUvQhsjYx9CA8ZSTUMezo9dBTeiv6mJt+HLPsPyNL5Tv6rV10tR0mVFvKlB0CrScJzqQRcajCGBzxw50k+n+4I38YFsMxiyOOtLBXrdiwPL2sphw/lxvRpazVTSwVCEFdaIWvpAbi2s8Jtwj4CgGS5lWRjqi/C/MABgvNE7MyiQE"
`endif