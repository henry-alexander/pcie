// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PqIwJXYfLZLhJ/rkT5uaaYv8i11mPyHcvRWO/DDBOJyefXynA/zedY3MarGz
PKNVdwWdYPwWixs34pADOmHEfsoN/4UuNZ0AD1JK9ZPTK9A2g6n7PZoBtjnd
+Tt7vc4ZLUgYU7+WmoDrNo1tDb1b5JSGBllfLxKlacYpB2gYe4piWg5sDbPO
N1M9Vndl6dzoRin6S6ESbOJ3H9Wit3OehMWEJI6VnHDkDiJy84M9g6rIl5Dk
eWUsrUY3yXTFwFhc5PVKszkOm86k005NzVjKm727Gkdi7lzGgMx6t+tQyZdk
+jN2HWa3rdwQTneAmEmAOzhJ8XuuDyHqvVkNskYrGA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fI1WV6elvyj9W5uBbzPkpUjaX+8cieB5YbeeTFFKrJ6vhR05TSRHTtkfrJk1
1H8ZaWMqc3tG/kPuiR80xfZvzTUOpUuj8ugO2Sb9z+wt8GkT8IyKjnS4CavK
7c4Y8WhOZOqTciRh/07Odivj7mfD670C5aoYGF4oE3w0uAE8Vl8y3keBvWVI
XjePoGOZt+0rky0Fxi22sNDGrHVvjrJL6zFeVREutID/R8bQKhBRknyzRiF9
kUwzbQOMt+uqM9G/poB7xBkU3sO+lRxsvdsl+kQaTnQN2seNacgSE249K1Ir
xKyoAOy9rD8vjXWkQkHzLtBHW7GpPWwxtNrK/YeXZA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
n0ADF7REOhbVvotAYA7dCmBl9wCYpxPSrb6lg9xhmgQn03VAOGGPlOwkQqFt
M8aDDuWiKLMQVAbYjEFWVcDcztp+2V6G9DVH5LtWfwzLWrf053ldgdK4XsZa
GvPIUDYqGhgkKubxljzkvg3/RxxNrE/o0uywduziv+uSCpJw/deEN3Oh22oa
14+ss9pj9zwIi5VyuS2lDLMwJlgSOJu1UauLhEdBGBJNoG/sh5rCBbKh+4EO
idFcDigf8L1ofTLLXv8aD4mN2LT3+jh5CJQ32CdL0CIDclFMI+08FmYIS+Fi
p+XX5L4JPtIFd3gPMOMQcuNupFgDcZdDa0+uc/GmDg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
W0bsrqePxRmuh1MWXrkRLrrSNyqWYlQLsrrk3pQsHmmK9XVCZwgmyNHUTWSR
5gWtPvBNzGXtpEwJGM5HndW8IhOn1t6R1fyu+pDI9p+sE6ODvhl7zG+Eo2z+
ZsDSwxX/XW88oroQ6XZco1TqdvROrWKnnGeUcA3TsDg7U6reA4o=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yKbZ1pACAHxcCmy99lPwzGgMnAHawCU+DrP6W6RDqd+7GvOekDz1OMKWa8yd
JyWsXb9qoTy2pGEXLyaM8IGJj/3WCNcFhNZseJtjvSLTZ6Mo6iVZYNJ6I148
Ukt23ehPr7N/Y6r75SfbrJ+yH2uoTMUwHxf4bpxZmal6DLQU2WIs8LA7Zogu
Mhi9lcISRI7zm8t/a8rKZJex6hpfZcmxIeHccDWpwiCsXZ+Z/PSMPtL6o9bY
Jdp6WabOn/zki3E78zQJz85YWQ+W1BLWVsF6AZs63ukVtZMLhVPJiH5/aPAt
fm+Ie/jJp9koG7G19LqAXe1zo75BiA58XuYbG/LP5Dm+J3QT7PY8tq8+N1pb
DDCTJf/U5HgyM8wTPQXXDw/Qkr6QKN8q1LC7FZnxxj1DRc+fPeVE5SUh3NLj
KrlhWSq1R+3SaQBk2Ajovr5Jb2vy17uvSPFWayW+amIMQTHv7HRYYgYIPazZ
Fft7Pb48TPTuJHePLzhxoP0nsuFuZZs+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
o8APin002u/1/PbvzSJ5prZk3aFkLj9EOuK44SRd3WOw+G3s0qYnzwYGvZ51
8peJf+jfaL3XOBJhD7/zJpKpDLIrZet07C62bVOF8WtYk3p/JAQTLhYSeVXh
PJ5Hq/ruflWKfeqsobBg7kO+9oy46LweqpqrPVxLEaINvclqt5k=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uJd1mnzgtprpsXKBqr/p6ffD8g5tBkYqMapNz5tfCK3bBTJEDevvSpUI2mYE
2jVqH4XL1PSCWXqxaXTbCZ45r9InTwQ4BnNblaz331D22GkGGXKGdogY71Ly
xJufXBgXqGx8ELpEkSRcFIXXvNrfKV5KU6S+kQgLsa/A5BYhccE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17632)
`pragma protect data_block
SlRY3XOIIiCcggabWV4Nqc32zaK2Wqb2dtabvzE/apCZ1Y71mKIdRFNXbnJK
ne2IfyjhLEA/9fqpl5tRKCq7NdocOO3Bb/ERUTyBv62W/vcWGwFNbj0zxs7Z
H07/jTkxMSoduPz6qPgHwSxh9anACyM61FOrFIu1wactkqrTPmi0vR8kvprw
3HZHjk5ohbgrr47SB/8WfD9BCmWHKN4blMsaYQ8tU5vScmo2pU3ei1oIxl+H
lQnWID+ZeMfCOoNPhnCW467mElODj6knKZAJY6TPY7kuQ0LIuopMqkl3pHWA
5H7qb5h/CibYa7//Z2wtDJk4L58Y+CBiLtS9esSuZJrZ0AqbNXVZ/Ip3V2Q/
J+S1rlzjfDX7aBlljgfZCLZDbxBRfF5h4m4lc0LfuSYT9tfVBIE3g9zJF6a5
G090IGSbaaveJTc5qUsLt0Ngp3TC+6u3uRy/5SQqn70XD3y9w24km/XdKB2V
W8HeYS54HmI3FHACHio7s6Go5shfmfVmi4pFB0qjvzi4zgL/7JrGf8MSWXz/
KTAAazkSwwRTRdqHsoaJEbQkXh0BraICc098bVduyWYu9o3DpvlgIirBm1U5
UBgIXsTpL7EbNr1i/rrLhqbw0j11Ljj1vohFKcndP2YhEFnW68pKW99qZbPN
MA99z7s0jpS2DaJjAs+1JCkfBzG+pls/IVbchDZwwVEf/dK8ST2swBjTAaWc
dEkrfY6sM1lAKSSnNLMcINUpejBhew2UCszgwEIb9X/5UwD4vMe4hlPdH18D
RlNjbpg/nDCvEJuYJ9d8D3sgguWa0bGQA9v3fkAER2L/roWkKcyFih283XdI
NCk/VddpaRBUURNukqWNmMNJWTgFusmVgJO43RwWjqtPvOs9gC6ItCtbqnk3
H1iieKmh+yYgKs76co4ZYC+JH7rzABBqnI57+uTJY1wvWWwh0RuS+8qXATJW
VJTBjPoHlhZxecmuUIgdv1nio7kI6V1hQS+XrOtEKV1Fb2EPPNehGX36TlVv
rEE9xaqIdgrkAay3t8ym8HjNG0Grdw63ecNgE03+fkl9I89zaIkTo0nJI40o
t4tnDaaO4BPVwgBMtUnW1wcH67mOA+N396HJ1+22TjDfbAjj/Qjl5h3k4vSG
e2SNNudelUAtWXAmfO0mk1q5uPwCXb0Hf0aGrVH/AyEJyJcbufCnINUiL/TG
L+H61aF3UQH6B/KYgofTJNQt3PNNERpGRvIXpoSskdLPsUYztPV9sBkRbiX+
VGTl1Qm9nCXdaMwhpWZk2vGg6BV4Rg5mgZKBP1YrtkwlGeC5ryHnHDa5NYHH
q3j2STRjvDlq0cde46KFhqfSdZLNRvqOmuEgYNhn7V0E6UQV2Wzx3fKNVtJM
Q1B2WUKYrO7/tnkq+qf3WrfZ9Ez8iLnA+md50HXESSe479V0jft1cH7EfX1o
by33Xfh4HMsWnRcoI9m4mSDXRXdXmazdEUCiEAi4yeNq00JYIaV9q8e4A9Ac
0HtOjSeKs70qSTm/ZO0E4Pxmh/aMRo3k4lYFpqBgCin0YrveiICg0WErL2ne
9rQcGo2Ts9JdFvoDGlQPAglpQyBPbQ4L1lhZcc7RThQ3up7k7WHWlprHQ/R9
5gHaEJznRLtjWw6Alrgb9UWa2Xa/38czAJE0U17B38HKh8Lwze9JOJ6jL4xE
nPFEBHZ9Bfx0276OUNofYcx5NiZVmeBJIwmQqqFW1RdmTHsa8nJl6B/pC1Zv
wvgBhwu/zV+l46P2T66lUuLROb/jUB74fGSxnGRq3MsxdzgqMTT9V7fzqwLz
HHkdaWzkW+HO9OuIsqG/0y7D//je48m75y/yDzJdmh4FhE/0a9dC4bget7zw
5pwCeSr/JDXjkhWrHqu8pRY7R3I0YPFJALE/JaIehd1sVPOJq/4Gf0HBuiZI
5tOeUcO/V2+HP6CpxwCPU/u6GqSayXK7iWYmVu1T5RiVAmFmeVsjD6BnVbep
Q2EWwaxUh1t5jwKrCCZyHSuSMRmlQU0gpB3PZrkTFyFr2TPhl1qpOAUG+9wo
FW7A3gjb/S3AuXnEAuK73VWnRjEWpPj7IGTNP+Jv86ef15eM5Q5FJ8M8GKck
uX4GAAtZWjPwBc0Kl8e1SlffM2f9e8f7MFU5PYdeAQqH7DumR0v9w3mujQeD
vzysrm8+oHJPtcrvgkI3LCUEKgGLTBMs9gcuBKsF4+CRMr17Ev8qvTfRxP9+
AM2PzLhRS6SfBmW1TBnutgf4UzhX9w6eRowTqR1YBoBxhZFkezMqYnR4fSfE
cCPBsQDzhfyvOd5IsW1qFSLQuDGMiIxVNS2kXVytn4DNMUj+QZqZdPUcw2Jh
dr88AVlwUqgidZO9X3nAcbEpG6MQ/xRipPUnuvcGAmxduTcQhOIkax7ADC4/
Wxj6S9TWye5qEKLl7Pn7uj4nzRhrrwqDdajZXf6J7V7s3cIOtL8GDywnoy7H
mJL+b5hNXTw8MFrrUnfRXQ21aR1qj4kCtOxKjNldjT0oIk30CXmQoUijESnd
ro7xLjTtCm/C0SaReXye1qSTYWf6njtEood5H/+Hp235C/mNKUU63X5p52Nu
58hNaIDNQlYieNvKDmhQfea9tQyuShfH4+9D0kPKyjAlmbylWSQnfnEI8ais
i54agnDQ9wTvNywlIERibSNOBNif/U5L8dq/bNEPJybndt6r/QOTfBehPZZJ
zHS2h4eXcIFF3hTbYXLd9gqpDK2pxS54t3uYFl1kXCnjeszwnUt/41YInl6+
rVwB2WIUjyLd309XC7nKzkjo4QaB4HuAHqGotHUpaT1xnu2jd5SxqeXz5hRZ
nCzaY5vRYyQQ217fL7t9vuOFWghcUwlHCrvCBanEHRlb8e3Czq4n4oOmAB1F
th7UA3KtltPIGUtujkD3YrJ4GwGAw3BPpQTkarXbNPPp4V+0M5r/LaUs8PZX
i57Drm7MA1tHjYXQk+mRG+cbm2OhLNT/lqpQVc93mvIDvpjYjtwmjn3qk2NV
gF0w+8CCCxwBBbCIhlC6HVwRQ5R7hVu310taOjwFgBNslXm2lVBqUGZZ4gc9
FXjFK0r9L+cp5CKc6UqWBDq1abVVcdRrFLl9dur+x9/9UjBvLoYs7gC/hOjz
N41MvsAfxYlSvT+cFp/qIBu+OtgUUpLjRv7k87hlXrbeGJgSo43CHWgvvd9P
wDVYogEFknbq3qXSW2pF9An5APgKR6TycuSvr4SbRKv2jlXgJds+ROW77n6D
2Wb6MfeI8oJ7BEhKa8fFNPEn+rGSI4Ty93Nkjr0XZ1fUkzoHUamxPePqbXAz
SHDvwylkrnRXtFLTUeTQ3I4yIY+bONDD9X4nn9NMjiSzJZqpGxdNGT/evvCB
9Vd7NlK6Bqwi2mlolPaEoR35wdEKYpSkLixiO7BG9Q2LZrD8fydq5dTDHL6f
F7BUUI8opG5bjTTppDxIRUFmlDF13R4AvWv4Mlkyp40YdJMEf9Q1yVfhPpfx
wOIOIkUJNEGKsBoO56igSKXQ4/aVr+axTnIO0bIg9sBDbHtftNdxp8hc1HP3
V3lffXP4wzj4lJC9BdEwviNw4kQvz+njjPwwUUJ83Z9zAqqATfE0O7q5Yxjj
sDUJTXlq8iLsepdG8taJNE7GdYauw8bFeEbZmoWAWKpxk5xJ6V+o9f08Rm+w
S5k7T9Elxb9KkaWX44QboxTS9hQ2pRjXP7zkVPhDG7ndoNgn/cN9w3E14orh
BofPc1zGFZUlyOKgqmfpSyRZADKX7oiNjYINqSPrdIK4C9FqzK4oektQtFfQ
f4atdkaXf1VfEF+lAnB2I5qMYjKJ/kGBSsuZhOmLkSLqITu0uDHBkSPhcVwI
23OwOck1LM5Jojna69v5BHcNVzdkfWL3qML+/82j1+Fy+mnJj+EZghT0ttAJ
+wayw1IbvRKVy48goAwros21CYuOPbuWcQIegTNjoypPOItjx2ExHrsbd+jc
Cn4uAjCHOQihy2ruf9YN5emQ/vLIKRGRukwJfKQ/zY7cW7xgyvFNg8c5cbRA
SIdbs/Vc4i6z78m9or/Qm0gFs+CjcLv1ZcHhwujFK4U9kKQPA0DvOxkPtpQH
xJuWVtr6oW82TdbmXIMgXbEJ7kFBWYvUiH30n+VZJW8WnfB2sooYQ6oNmKml
O6ySfw1vLF0PUMk88GHz8YisOV5GqKaBHYFscxr8zufkJDI3McvMFLw7fc8L
2U0x1WN5/Dd+uKR5zxDezb4upGNHzretG03B+FCZ/mSPJOWxacWWtNzoiJ66
tyJWNwPuxCA0HGSyS4v0LD+nhoNAgEbZWHOKvHN/j/25KYbXqmBcqf1u0qZ4
dvPcNopMU0yf5kSroFNMgzcuNqg0sjUjvIkFRHgbkUuc14+J++6d1cZznihW
CemLOA+iCn3DlNdP+Ee9FlQzkSDRzOBnqvGxN27mnrMWiuSK3pqdSaivC7AW
cGlE3b/JZJYc2rrCA5wImHTzrK1AVAHcVOk8e8KfjyN14zwMZ3UAWEE6mrSd
4lRfYyZqE0eDb5d7zXe4o+MuhtpraBGpr5VWIz7vBXcMaUsr3Lrf7W6KIx11
DjANdbiwkoc7dzO3JATZUxKC6kU+uKSR17UmflgkPuwCWSr3AJZZ6pG9tCg2
ollP/M4Z49vVBzKD6MTP79VsH3jLFfEAVkW5XQUBrX+9dhn1pu/Hx7J8BVFk
2i4A9VZgdXtXdMbih+BNF/ct+IPLvoVq+7792lWFvUFVd1eutBe+oTeVYfhW
xTlMqz6PFNmPmFgz+nHavSIv+W8IgghFnAaI8Mcc/MpWcqBc/UAVGt0+qbH/
49BZVQ/x13+ifYoYlB1GcKxejajzz9Xx1uSzV+BKmgKC63G8YVDQn8vB4BhZ
E76/yR02IrPsRezhmACPcfxyNWK7At00v6HMaJV19q1vhCIFg+oRjCKFxXK5
ws5c+6qkqk3H4JircWX7J/VyNMknSo0KmPH8qvzh8bckkUuLENmfrvSu7jNZ
MCQEp6X+oqypxHkaVZr0sO3i+3rn3jyT9eaixV5JFppnpX5EeIGwrYA8NXpI
6EQEHc0Vw4AMRtaTaRqRcIIRZGK4aaHkvlo3kVWMTHLxMfMtZDarysAyxNXX
OggsMN8SKjk0RlH+ydqHcmQSrIZYoJ4Mo04AjdxZAaBtK/TrBqbBet/zy+um
jLSfiiCDflAINUrIg2V6hVdO1PR30MRAwLQPwRqZL/I8+F1vxrPyLZF3b6ud
BjTUS8c3aZy2uX3dkVYT+EOvsUoFI4o36o9eGnRxpfj04sqLlUOmjMe34eEQ
vURDm7w5MQuC0sDFYNE4HE2BWSUc4VIkoFSnmJG2TKJ9T/ms8QPggdPphzO+
2rIf9YGJGI4MKjDQuzTJoG3HekwPOEQUW9QrvzR1DeGhbJ/rCIqMuBXrV0WP
FYeFzkk34ZJSnJ5UXKAj+ooh4gO0LBcp5lk1WqDG9RtAr9wbnbpJcJOTwguK
S3PAe+lZG5n4VruJaqUngbMeFIGkBfhCE6TJMldfAFA9qZ85i5XrmJB2F2xB
DRa56uvJSvZv5wVC0s8UeAfAawwYhB8pbLZhlpkz1dcE0qdG8lWbiA8zPiGd
7DOE8rTIOZpW+tnaGxWBHp+eceIl6SPSFLge4aPNErBpl1mnGFbIj1klnFxI
KHAOKF3FSaUnwR9l4TYhXlV6uXqHWXITgiLRLgyOLLDHHD65yO6DPpmt6lQ6
mBTfF29I/GF+SETpETwpUjbElU4pzRXQEiOSfZ96FbP7NchucK/7w4sGz85W
idl7TFc7qHHG6lt/96+4DdCu/4atIu7kjFhosUXpVJ/2DCjF5TbjqktXJod1
bvtKaIAK42q8thWQbV2ySZuQeCC77X2TJoZLJds0XasIB58I9o+DKVRPalZW
6sPjfiJlOkD0s8jG4kJX8sL+Eor2rinZ2bJGDfmssDvs3l5R+f4wyDMm2ZEF
NzmVJ3a98ILPy9Lo5qnsWxhbJIGKsY+z3R1H7EUGgYsgkFg9Pm2GKAxPXlhI
wy6+UcqkiZHsj1NLsR+TIKQJb+w42btIRq58IOvSOetO29PHeY8gMSPc0g9I
COBYHGxRGz0Ld0B5+k285DcDE1IpG0cDUovPSFLF60lIEr6UtTad5h/xNifB
Ar/g9jB00vzCzYQHcnS9SlfFWWF6z2VkCOPdWfy/PSMC02PzizkLPSij53ZH
nSPuTpw/mc8dm1C/flqSACfFetRU3uRaE86hZ958M5yULeVMyDsTEE2OXYjE
44b5yVpu2WYfc1gDvLvplBkNUbiAfhTRAU9VtlJBMbdN+XbSwn34mUmzw8sf
YEG9nAxGGrhl6JjVcYGuFb1lZINj+UG7v9hIai+3rmMzmtDuB3IlxYwWUT9h
pc2y/0BB2GoA0NXQAPbfpgZ8Nv+JiEeD5LrYRFEXf81eer/hvOAVgeJfQdu1
RS6KThPxWTVJ4uq9tX7C/5mDxGHvjXVpn6iX9nY8YifyccWK51y7S7F6pvQy
HjvrF3Eos6P4cTOf50H4tdTrcSBMth2ZkOekym1A9sSxOIECPEJ8+xtkMj4B
TWhYSGFamVZz5Ye045eyvaYPeV2PphSiOg8ntiQjA9d/wUcnqdvwIaKPSt8F
f4FOB/3JnpLhHC6nsbSdrz8Rf6wt+6ipxLvtcSgmbMjdzTIy21tXSvzrnrnb
2qx6txrSaRuPJjW7LlfTa76bNcJiKd7aiQhObv1qob3XBBqP/1UfoL82zlTd
UVu/7j0+btGWZSL0BV1fKIFZ5Dbcs5Y8QfNc4tfnpJKwR8nFk8UzQ9jpmXFo
2RR3/0bl+jvBNEn9XPJdimsPOTBVYOqyJdV1aBEmJH14A04D0eWhZasJ11XG
H3QHrHUfdwp5tj8riucZldhPZ4d+WDUeTvZzW/8SLbqgKz3bUNsF+lHbkj50
CDM71kKLg9hHQ6F9iwXsVP8ME3tCl+KAKwFMnBpf34mBh7a6Rn4witMjcroP
1cZvdwNuYWk8QXhYs2/uJ+k9XilKJra39L/3PJldxSw27jdF7erAFHBo3zZ2
Vf9tvm/M1AF+oNKPJGdAqSclA/ze+HpLOP31Loi+huTOA4P73iBAkSQfXqOu
WxQhBAV3OPdDSd1/eVA08X4ltAiCnhVATcKJP7CFlIY82DlX2Kc2KbViWtWq
dH4j5+zEtTtzW8bjYPGB+T2bNuQ9fSrZ9zzvxD5g+rgF8NqComy2DKXYjq4s
gbwk8oRzjRwG7jPggXTb0GjqOhmGQCuk7JgIn3LpMjIKrJTDNH6V/Wrp6aPw
7C0OfXkB8yAoCru/lUjkwGvqNZGjOVNpbejWd6FvySpBrfoU1kfeWJubZiB2
2euJrrE8X1WcjGbMX9688VuZaMbp33D0HvuqqiTAqnNTGaiwB7Ar28FHjwAK
CgKST/X4yoMHzbBBr6a/Na5Whgx9dag68/Vd0Hw7QKQ3+C5BS1c+gG+faia7
98k0zKIoNuUkwzephpOCKYVIVWygX36yk57CTVTowoWOTlQmG4uTRin74m20
SE+jcybEzgJfGJw0zFyBXJvO8Nw8ld7ambll0NiiO93Zltbz7Pm0cCEZpyZO
VSDoeHtusZVMtgVsy/n614ZRqFbLeS8Vafmlf6LOBk8elkQo8V84AqBQt6k+
WUIS336nF2+57RspLBBapiCOm15W3/7GezwfN5NQ1Z7Gm1II5t3Exif8WRcE
YpmN6hhld3lES2KEzRUqszmebXHG7VHEjnP0vFbeIOLAg8bd8rOHuoQvUkLW
uv7RLOLCk0ercMRnpEigqPkvvXDbZ7jX7MgXlU4xBtEf9jZwMWWxSgCcIGDl
ALjOJxH3e5IL/puoCHlIRlRwoj+kejGS+vL/xNwQgndH09G0kd05+Ff5HIe9
+bvTALO4X7lxhkIfdKpyEN24SbiF+CPt5S4tuCCrV7Ux2K9VK7xeftF6aqB1
iYDLmX7fTOhPQiCdUmFN7sXJDBbZI8QfafbbXfCDOcu0J15yCYgHW6DRGQgx
saUpZr972GDZwh74Q3LNu+8u9iIMkE5Si7cNJk4lEUcpJSMYIv+YQ8RUdhSq
pN7Qa0Mwf3ABAv7EaKlEQJ930B9QDf/lPgksWjgGTpWPYnRRKXS3vG9r6ANm
BbcnYCoX9riNdwiINz5V2FYUrDviu1iCBkJ4jDzt1SloIYZrVmyBl0zMd3qn
b6Kr0PeqUEi16Xtbtq3uSYHP/Ogh5FmsnovfCsjsQNP7bffhb5Pxyb0XVNqZ
w9GvGBt89M2E6RBboCNQPeMOAQmqXKzPr72v7IliGsZeUcLbWtM4FGTIsxhZ
fv3pgHMBOCNxqRqABboHI5TfNMEVCXTjpUSU0QNidBj+jUcXws6QHy0x2S3t
+hxloOan8i2HeQ1LBnUyFsD2L6Qulmz7ZC8a4yFACIs/SVnvFTrSTKc9LDCB
FWcAlUtqEOGdZeUD6OuK6eiLWJEBJfPWvnLfxp5AWWPxTSE3kgzjq6GP4Z4r
B+h4ADgYJpvmtudf64laN/Mds8Axb2pWzex7DWsHb2pO2710lk04J6U6AODD
dGQuhpE9nLBisZx0eK6z+D5oThB8oYGie4KeQ7HcHHfLUu/7Ncw9VAPJV5jo
pydABIoB8L3Nif190hi60HaVP0+2BN5Qqh4k57cKTlQKtNK2UgkwvSY9zJSk
eAPl4m7yph5EJtpruJPTEStbX0+4Ej8yG0UI2Rh7VadLF+7/j4+vEZWPRSX2
q+rVeojmn3iXsgKSoSNIP9mMxqk/pLmIHW1/fXU8pK1hskyP/ZAiJIDg7/gy
6Bbm9G0wtyTpDOh7XCMGMwNzQFpyuB5sbOsZGj/U+CT0XnWmgHnTo+8a6NHw
P7vVg0xRuX42R9MMVPFR/XSxywxyau99rvRbTyg+tbSMF66f/XnUp9OGRNg6
Fbo34THioxbE8iHMQMHH5h3C63fUXJIIU4ftYEsepdarXk1PizQJSUwjJLSs
Jtg+RZ8lNGSLbMrfVtQyRVnU5AupYhmFq79h0d95gx8PLxLA4MxGxss6Niyt
NamAh6fL3/+AKR6/huSWZr4IE6d4rwArhZoQa+HFkj9vKCPvG07uGMJzZ9Cw
0xAyJcYA+yMxeOK4CZKALh9WafI4rr3nfTHfqBVtS1YhWwYYLcFXRsOrYite
p3dzUMw3yN+cFsdVFLoHa+W/bnqVuNqsTrlgq80JOo/kn1sBJ28ippsMvQr3
MPcaqNGvknW9k+vKOkPXAjLRjWVW2cih1l1FV603Vfi/4UyqIgToOlYXeUt2
+M0y/cmgpemWFu4xq4zxJA8FZ4d6eq6cAqLPXTh7SxBaa3SMzmz2LVr7a39G
vCW7NZFfwaIeRZ+UwsWavjWej4WviKbz3J3DC3xIvdOmxZrpKeIHqotvi8oT
K3A7S7LNkZT+E6G0iVSovu1YmxizlqSNvQuCX3x2LlH70Uv3AgjJmYXw8Qdw
umtEbyJ6L8Nca2h/Es5n4qSVzMm0kDcGoFxH/wWhxaX4O4rIgmuYSyQzyH8n
ue/Ge8bFKbevBVSbyx0xHZt97t5JVo7gAMKFxbaG0gL0dprqarhJHxMJR9jo
C4kDQfIuKYUCTrdUlA42zD/Iik0yPFnG774baM7z4hEiW7k/RVnkyIKoI7PT
KeskRTzfacJZuN/gt+qoWkjSCIpIsW8pqX00smXiI6kbB6i70orUxoWM5KJt
kGFBBbKGadqEECWYz725qvpkgkak5zuwytP3bvVCWTyMuRfcF5iJDUDBkVx1
mdjq+VlKXKj2yadBX29H1zqYAq+/lyqTN+Op1XKhBHvr0gYm2vBbCay6+HLa
mPoIjB4PR/Xb9+D04Kj3ls5qKda5scnnlHKBe6ujQrTJZq4gKDDO9iogLbjL
rqEmEpapUqJ5K51L7DD1eLPHaC6Zd3IEyMcPcIvgzRGEoUCbq/Mk4WxGpRQy
nT+bRWtGTGM039CAkE0N9DxFpv9w+kAMnEaVr+5uIvZ8wzRLji0fdeaLHK8V
0ubhnWN8MdedBY0xJ35m0xVhD5SBnnpMph9qqhonLMiPQEz//n2tDS4a8zFi
gyhYUNhv6wM01lMVS0g4jIFyt+V3kXABUlOz9rg9aqyKrsQlNxxrW8ivgYd0
30yXekYjX5bTUFlLVqCHDoVEvJkOsCJOmIXKmSRtv+RBIy2rSVMaqwA5i6vc
5rgOb8TkxGjW12ovao88ZAUvIUDAm2QFQ0iGsaB4HuoEmzjIB/rZG/Fb0Sqz
TgNTbMMBdKfNSLF7jdqn1ILXxwT5sBPzuksDd914/y8e3rTyS/HHl3FkP9wl
QYXTlc7h0GHsIiogjWlGr07X/OKQ9wSq69OjwQ7daJpKnN1F/jOggvT1pl2R
l1SogLDL/B/nyRZ5PQjsUvZ1xmNSaSepM3/wUd7YagTQKsfOvE5Et/QBvjTw
/LpWvNYUWyJG0tiudyvYm/EB1/3UiiAUSo7jE1In59sub3e2pOIIq9tvGOCD
4pbQx1w0HOHbXfxzwfLWkfRaGVAa3Oof1CkizPR3kqz38x3IPnHnBUEAXIqV
tb1bnkw6aCGfRumepxIKy+1OhfrEh6qAllbIX+F1jnnULd/wZ8KuCppk4LXn
yhNFhd3sgvORETargevTo1cBSH64r3NNfakzXcY7rc7T+7D5tpyJexSWx1GH
4vovBX/kolrtUWAKXChWyMNvJB0lHaQZCXIOLcdgc+chaXW3pNVA/I+XPHpR
9zEao74Q3ziXf5kWqkFriO3DfWQH0dVfO/0b3sQTfTNUSwYiO0GS38l9JF5i
pqbFoRWVkLM7cn4i1TKFig8s7jNYwjz5R/kiOW5XM3e6PRpmS/pnO9RAA+Vh
bB5QkQWuWmIdVq9I5p/1TIRLtYw/q0n8GRWKzAIdP3x9rT9cvMovSsVFiGee
TR7kZHc05SJIZ6YSNYQ56iHuXFZwQaLzEB4Rp84rckrcIodrImn4MA8DQnC6
p+1Vu8QV40dPVz0BAspwPANcCD1Ch0EqPH+EgbRaNdAR7dGJe2+Nm0ED98Qd
r4GoWU3rMKwLAZHGh1NpBY68jztFZYRHgJDNt+/gciSPWjcOPG8zg04kmYCB
hSE63mLLUikG2AwOsylmkPdarHLpiRQYhRAY32MVn3tFx/+uS3aiJhAgk/IY
9BLuccX1xEwYAf2Qln5aF6vmU4Nt5kr6tuGexfe9LsPIB5T3HSsRtClAEwon
aekxo40a7UMDQl85gEvA5wlY/EfPcDsku7pPQk8KWc7MAkrAS1WXHvStCxis
semfv3vid1pvq4ffXUzY1ajhUob4w0ODoSSxHYflVKp5qTieTT7XORsF6dRr
/FAxT/cwicCoTmisq8i8Jk+o/wHzbrhDZJyiOnPSeJt5npc4zIwbxjWgrPsV
dhAPAF03ewH4w//3IxcaEo0gFbgdpGm2zVGoLfHRtUR9zmFhQQ1g6jgpOr4K
eG1qYsOb6F2wgk3N+lVeVFPAGDtw2RuK8uMPK5D80UTUEK/+IWaY0IxKyAs7
2Pqm9XD+7ANXvtosS+ulfeQmuU6+0LuptTlaeO1wXNYrpXB0mUeGYg0IFdrV
HdAJjY/g6gfWrmv8jK31MeIAqoukAY86j7IPITaGqD6GqnOkVyFbXs7kZiRZ
IOImwPnKBiVBhqQJgc8jPfYrOYHqci2CXyku22SbsPnauqp9y6vAF+EAFDT4
eaApJ+HRvRd2qzaRrICaoXOF9f9rQ9TNuxc//MzMS3/Gmcm397mOJFoEk+8G
8oRZ3ih8V5pd+ZYS+hcC01lE+810p6TpYxYo8NTzmZOEE7ubM4Pw9sy96Bvh
W6OcnCR0R0ec0kEE+8gcDAqdpjPiDvmkw1z/GWCMOC1oiId48U9AI1N8huxa
xIweSlSdH87iF4AxI/6gcbwxS4VWk8VNyUxhpP8u+Ay2cmnXBsksrwCLmWq3
UYFL8jXygKS2AxieNNrpsYyab7m00wRnrsiPpSYG+9L7YkqzIRvT2+hqFMgE
M+G55lptdoYhoV+EqnGOshqqCjAdrta3nM4QXQWpU+WcAecIjGLGZDB2NCXM
SGUZ6u12cp7qysHguG00cNix1BzEdjP4A6vnOnk11O6NK8xGfqT+MwsSTf8M
A8ljwYBrEpomYJoCpLjAB/xvzjPX/shwWZjbMKT2j3t3N1dyj5A6UGAfP+Kt
icS+qRWRTLfXvatBKYBpQhxXHMr9KGI6/HlnBhGcwpU/CPn6bVrxlS9V0EmW
VruY1eZWjOPCcr/AvYbpRHQzYNWdoPMjqLiSU+kk/ytiXnF0KULYF8VCtcvh
ccC0S34WhgoaBbueuGsDdoBvE+bhnKrDhVJWhweYPsCoDcUcLzFYHDcz0b87
UG2uOIZaKTFwuBnvxGTnBl+LbwszvjvTF2LmO5EvFzm/jj+BQDWgUYGK99r1
kVw4YoDk4/lMDWT5xg9o0lIuYRY23pNCr1C1NR6SMwCOLnnV+i5PLNysfpnA
2mjNO6/YFdOywv2kcOuFPXNHgXFA+zesX+T38g1qdBfMAnt23IbIrgqOUKRJ
j/wlmstWq4Qb5mSmS9ROTz+aQ5UgliOOwB2fQM+yGVcEEkCC2Tl1vfbJv8Uy
9eNglqDTHFWuEatyq7Y+zJjBJjKCIYZk0FX3TjuUpAFuifd7Pf68bFjE4eLc
a6r6MlmOdydMbP6fL07JnRpG1W+eStOesXvZU3OKEmPAk48eLK7YfB5RRYYU
rTtRnSSNeGsYNF64EPnartVbW421XAdYj3Gx+sm7f5xVUhZOpHtfe6z70IqQ
XtFgEYAm7MCTHBlMQDHqi1j/8+9vvuGRVMUkzUUBkaRrwMWLLo7xJ5Xqi8sf
szc2mUMJ7Gz+rqSsTvBdaItd/8ldkOq/RaehWBFBTbV4G9x5VK1tLk12pu7l
9ZWWA/EJhWPSu3upma07rmpLpUeYSgke3iB1qcoX8Wlv6Xbv8ibBBmHTaJia
GBsd6kEZ26HJ+lpU2T8swdljD9hF/6+3pq3CGLEKHWNknAcMhhK/34ADWgfu
f+F1pUZEuQjmmk43NoktvcVCfRaE4vgNqSu/RgqvEFJIHkJOWiQDEm9sEstV
ju8Qf9peCzayhutdVLsq4YMQ9dbQrbvvd10+frQwoTdk8ZnTR7FHixmE5FiM
rYHersMN9eUq16AdlOPNZeK46zqcs3q7ZItsoMNh6rjoVWKQ/wP7gX+rzbNt
l8Q6yZp89uEL2eaDahTYa0Ko1ZO6dI9Aine1pXasvw1eYkc0rBidvHItLS21
u5i7aP7Q831tCCUAn60TJlHL2pNXNOOt3neY0PGPdnF2qwfZOhrqDTcMfK+N
uUIKEcu8MUgOW0zSiuwYcAtptYB+3EWsee0EFHpVhqR12uMsBGghg53XZe34
NaAQK7PR3gzZtBZtyvoG95W2ttvplwBhgYHSJFWzSEfVEJZZj02yURfuZOcR
oKVcf8Ih+aFc/QKNGe2ylh4NVgBpy7hosoV3LpCilrpoyQ47QRAl2aCk60Wc
GudDxYfLQUSBFiyoOT11mnY+/g2jEPcJn8BW7vcVj+qRpD6fwip+h9aG4NWo
fAlfel+QqKGOLZAuVsU0LRl/V45fJotZxOq2gUI0XilJIdyFuSaDTqvzpN8g
hwPH8qWSNHwW5Er7C7umejOD6t6v8rwMNEmPPsioOR8YGivODVL4mfnvahlN
/mwPeA+VdVlMhyNW/MXlsVuakeClDGRsr2GUxIXXSK6pBhIOpQnseZ7looC4
AojoY5wCLZPYTGPrNPZQLBN2wDMJ0id7PyDYZoEITG2ugN/qIuQQHuQUHjs0
aItshFHCsXDgnP8kLLa/CmB+7nj7T7J3X3gLqtGrXqaRAXkiUBBCE6PKFl2V
7OX8MOIuFM1O1J8gLUb6Wb7wZ78zJVsqPeBAO0rRYKzCIZcec0y77uF+x9Qi
JnFGt21XbixfiHUdnR3h0yybosLXgkJXAY+Ti7ZQuYcLwdy0G5qkiZccwA9S
fP+39FjXidgg0FVCuDfzyW/nRD/yejaDH92GRdmtGY3tnESXX3FpFMEmrqqk
nfc+k3YSTIh2ZgGGlIG1O6tcegErOUeHuC93JWduIzkOlCF07dASH1fEduin
eGUZcX/RY3hA0UdTzNl+/hvRZssGHVh60k0v+I2K86EzfuFvu1+orNJdw6eg
LTpsdI1QeVkq5qsqFhQHX/p7XHKRjU6YI75prnkNwL/tnhevhQjXCSYpNw2O
y91pM80AkHd6lwfEyeb6mKIkZa2G4JfZGUcPuLv5RlRGGL4y/1PTmQ83csPu
qSYzNTN+B9XaVeqttDDq0nUSCwTMn5jXbPsRkl6XFoX1YPpnoG7X36DXir6L
GCovcWSIAL/5bO5iesqyYRWmajJJtQTTeKrGQ5m0gYKNAwDUWVU6fFB/6/gT
vxWu7PIodoMsIFCl6x97EZjFAC+PtObkN2DWfJTgxN4RRq5s+zINH/OdqUVX
8LgJ6wEMH0pKDy5zNe28ytSqBmQKX4W4dExLicsLdTMvzQpp3BbvC7jGkR1+
bbju3MxAx7dKjkXSDeEqAECl2F+TQDn42EALMfjRvDUguLUIdDAQNuL5ItRU
M/4DZ07dICO7jL7w4kFxp34MmVODfJ4CyNDNQeIDZAqVXasNuqT+YQGJA5jW
eoGMBvSZ7jbpNScPOaW9NFAySk4DKjgsUI5MlDWDU+cpiPJKmi4tS/XYSGyE
P85VnIfyfVL3Y9SIEb9J0LM8fFSFRQJWPw/LK04Y/XmW01y0T1W+zbylwn9o
ytOU6L7dx2fNkzRl5YEmguhK64uNjV2tH3VJc3JBFsmRZ7tL9fs/4ZwnQL7r
tfYsqZMN5tbBnBbcWuAvEIeNCos5PupQVdfENWrjYEWZAxD+BMiJ3EgDsWid
sgPGgzIo4TaIBr6goKz4+KjMRUTOAQq2HLaURzsTu8CuMBVQL1JPt2Vhqr2D
wTmWUqrPhc825TX0A55CZT+wolH2XpwOQHHnZHS80LobvvZpckBdU85Kot0b
MTx0qyVtjBfalVDpwRsl1cv2cOafHlzGJNeWb58hYnWa6EQvlX4E5nvOHkGs
Dia886cACyk9eAzLSd1C2iV4felyDAAOlgpkQDMNOVaa9cjKF58Cr6xACbAi
Y4GCGZKSh+3yfVIobWdO0Pr+AZhL7a3JUwk8xL6Pqt1qbls/1ZWhuiogMRGu
3v5iHHKNmAxyfhGDXmcLp7RGhjIkfNbP8V1ZuRZMed38L50cpYcFob/rXl65
mhu0etklEe+DpOzVDQpnfiuwP/q7q+EYbiXHpLfSgpBdKAIht48/IAnJbrPJ
CJ9xaX5uMUpHKiUqPLOnVxRhsB4Tvo55/mLCcG2kwu7RQybEMGiggEWYM0NW
kzmrID0rCpMFi7VOKZgsPDFTX269Xyc2RLxtgnKvevRB34sZyPx5CB6Pq3ke
pdPUpQN97LvmV1gWILTQBjPmRUUKbE/w5ISMLiGkmweewJ3ukd3gT5gIYPyU
akTLnE5/4KhBT5/vsI2nvH72ddHf33v2iAOSz4EsRQsd0EuFEP+jnTK+KKIC
WUbUhHi4FmHl2HWOMURxu7uzGOHguOvgVCZSqJKb8GA85/zTFEUoYqDLZ6MC
Mr/p9nCePYH9r+Mj3yepdkMuF8lh+/9e6+1dONn8d6X5HqNeB/tGDS0WQFIC
9slnkcJuA0Wa78pUb2xrESWaHtZYJPixrOIT0c2s38H2GBTcg17i5tl5BiVS
4PA5kSuUN+J0HpvfKwdIlcZekte0BY+8T+gkrSm7zsoAH7pVsFG8bzz0wVPs
h4lRS7KbON5DjfnY2Qfvu6g8OibltNQ86XVpJ2REu3QG+256S2MRu02wFi0a
8ypipi5U3IBCvixMJVEY1AexqJB0/PpRZgtRA2LhNTC4TnE8J9RMk8BB4z/8
8dR7VqJRTzcCJMv2xTwUqHBpwgsmo4AyuUOaLw64rkJ9QBiMoS0kN179w9U4
ndg6xi+VHiS1QzCTPk3ZPhPiylVY3Hl1lvN5zJ+VxyBlEDnq9am39UEdNFZl
uK5epMVCK+yMFxA2qZeueJcuhETPkQscpl1DnZ2Byjx87T/7w/GpfR8S9UPz
01Za+2QMJOpYdBvStuLsGSru6hj7IbssgiQPRKXzPTexpKaPoOPh8jKs/EHL
qdB4vqhlHa8XKy4/vJ5y9fu+a+qZ7hvpFV6HXnCFPvXpUeA8qqLjZOa7AmNH
0TSMblm3lil/z9WbkkX+2/CsFfOzUTcLUJpuxd6NBYSiEe5XxFHjjitPq5Dh
nhmsZyQd+BC87/y4kMw1KorDy2T4OIo6+/RrYoS7FHtplo3lmKI/h94sctF9
MY1N3t9Hi5Tar3dNaJtEj6UT7obtuMlxzG1qd2ennGUdZGWMR3G3Nl7JQHd+
KnQrzj0yZ72fLyMtJ0XEosZ/HwhLu0X0H0CJmgkQUofEck3Pe7ytpqom666a
CP4D4BgphSLX+mw+EU8QBhOHNoMbSkVvJYo0Xu51Et7LGTWH3xnJKLyjbxpw
Daj7R9GBfYZIXB83QbwvanknZclM3n1mFefD+WgSwTXSRJ61kgFtwY8qTqO9
FW+anXW42wulzHBemxDaxLZFbe6O2lw8P6PkWgLPZ/rQcypgavvyuMvt/st9
CDV4IwJRlMAJ8UMgTJ+FxZ8B5rma0X4NrmAun04OLexNFAafyzBMVbNbVKty
3OGeRIoLVrF0ZcpEZGHPH9Je+ZAB7E570VFwe/STogBKILgdsG2UYwqkOJBf
CjB5XBMgKin+IhoZ0hGrvYPTCxcuD9uqR/fVxwdCp67Mn58pD81YBQT9disF
6WQIuf8COsj1xeJ6VpUzbXkAwhHW+198oM0tEZ4ZJ1f8hgBlV4zrLSDAehme
o2m0JIFWXwu1H4BOsCnkkR/HTBWjvJdtfxXyRXk1w6+UwWt3zaNxCoBwJe8n
rwbL+rEZMUYXEakZ8n7q00K6m8opxoe1vQyd/HyaHvsQFQD7lDegMSWc8PSq
52UPISCkQiz3EZL+K+wQcR5GHZ/MkRPhFmwMt3dm9UrwuMNF91ToicEL83ym
pBKFD6p7JIIixMU20YlTZo/j/NoGWkhmk//nfCxA1H4O3TE8u2BF9pDc3pJV
8iGxm98BvAnp1MEifk+WqrQbfr/z8NFamxVvOHA77jYKbVfYPXQ7dDCt/sJW
nzJP8/m9C/WGl1aUKMpwxjud6tyKSff7SLIMEcza17YQv2+sWVzYjIVep5kH
TFnsDdGt2Hwdd7wzWY9cQrGwMTAqtIHGIi2g0Ezj45ReCqoJAlHKDUPpYmF6
iyXfUSR/zU5Xf+40aum6vhz/VzVIMAlBWrtFOwH7tQEgNAysy96usYqRlj7/
e23fU+MKQPyooVWkX0xNtDt5CompEjfsDXOhIdl8i+AuTDK1uvQo7Voo8QBv
DG95Y/jyt6I8oKsBR/aDVlWXZZlQHyf/zz42FEb6KH1kYWFYY5dA14+GwDJ1
xTCunPSpfQbIkZuBFgnyITUaYnJZUKZl8lc/qYyIzid0Qs+9mDIUQelOSRZT
4AvrlC61LCWyK76O4C8jJ5sdZZA/Wfx9n5YpmochfGO/09SQ/hokTdZg5dnQ
AKD59aPpSFHiBvQCYIm1pAriFAmM9JeTKno85ZSPe/1F2aTZ7ZAgF7N0lYHU
mhuI02jM0ymLJOJRg01Q0ZB7fKCF8x9XOKRE3TnGf6DxdB/Ha7cpRJj3ZYY5
Ug2UJimS58ESOB1Rb3ENxvzkBDog0bHw29sgxgQguX5gr35RUb0u44HCi3Wo
8YM4vaz3zX0//X/BoGv389pjxyOKsIkDsCPV6/S4ASibc5cjIYsHWfcc7U/z
GbMVR/G4NBHTpHpAVJFK7OSdfDDNfcXzlMw4iPDk/XH4Gfvkxr36Ixbivtg0
p3vPLOCbK9OhgJA7kmjQTT5vGoaSnRJfynjPUXNOC015fHACOk8fJExxZvcR
HeQ31NkZD2IolWGja+vAnnGzjUtwgnPPT7/Dz9t29MlSiBvd5B94R10QEozI
ImfxxU0KC41C901Vh/35GXd4Ml2tDO593gGESGYcPSI5pEuLXx8PextCFyyY
uV9LcaT/p4OkNaMgZV+MYKceNSLmEvWL29bNc3neSeg3MFlrf9hZuh9w82mu
p4YnpNsKBPNwvQyPM4G3tWkBt8PIQHwNwMz6pxc+JUGE8U3BwFynddEgbSIi
vrZSjVALLVPZguQY5EOTdhWg+eC18BXm0HD9OHdBtD5nvdb2bgcGMU8xD8DE
P9UQ+hYAyRhmNh9XadTe87xuuBnXDakpAkWrXQ+AWEbDgrfW6eh3GznOf/57
BAmiSFxRYOdENBjRALlj4TjPo5AWSLKDEykpDxcb2dmFPAln0sluduIBkqi/
ao8kIFFHMiqiGkofPXqRLvLD+72OBJeKNcnM0Gq5EujewAwWnTOQfJI9/oCj
74x4uoLMzzPUrnN+JeDKtx6+NgLoDfmIp3xNvJRuq8/sg+qObK7USZ2RR9II
fDsGBmqIUkpCFR2s1S0hpMnPFa5y+mG5xcUDWm8qzkuiACVlBZtc8oirNOIw
G5FMMicHnNBFL0Ilfw6U7vAGESG2vXiPAYgzJrOu/MG/no1OihIU01TWKrtL
YiWwh/s5PcOU+DNRjC6QjRo/Gm7TEnKDXdaxeh7NQp4gvMx9fryp8ijfjBMt
XQDhA0qp87czRzYtBQKvowx+aZUmCNGDfsoIy61QEd5XeUWaFeI+5EbJ52IP
5i5brkGysC94j+QH94oh3AN3DL3RMG7ABg9rVKFq/79lQL371DLLCWtLgTC3
PDTOy08/wvWkweF8dVq2De+TJLM19L3J4KpuvijoMoWdmsAoU73Wl186flA1
fnQ/X25fwXboP0DVByNpxy9IfADGKIYYLLMcar1O03FCaKY/off75KNMY5NF
m/NuyoC6zvAwfFRQzTcEQYOGDnUXHJeGoAJ4iGZEfOTiu64Jzl0mdGKeFNm2
sbb43O+hK4ZK9hJ6aHyFe2vdvfy8rLYLgSqd2V7GfR5RIrfH1F6A4HRBDCmE
9JZ0J30tTuJ7lLkfyVxsEm5elBXlEkNkl8pcaTgfbQavTG+pIyKBFZoYdqqU
qW9347SHy1DT2e5ohdoQ7x0dyafbqdWIcidT3BD1ohm8Cgc5ERPVY5nb/Cpb
VT6pE50+rWhHD/Cs0UC+PSgSOpcYrPWKBKf10kVvFzYAKqnU8ZkVS0rNdDOK
LaV+AdEw02479V6knW4/l7ZEtVT5PcASmyDRQSkNPvMvtzr2pqRVShPHl+yH
B8dU3z49RmtZld4mW/XzPZkYEN0r6Ah9QNlHPFJDfxnO5HeAnwRroZXn9asZ
z180qFLo/MtEXqzLz3md2+g+jTmuTvNfBV7U7BOM9+BNLCpBnsXe7qONNLMp
/i8Dgj8rzudtug2yXvuEcsx5ynKrSwZSu6ISfSByaC6iDH7l9dA7wQBotXDJ
CI+rKBxvCT4ZfmvfhInIBv3HRUe4SJmtuL4jGb6eq+2pJMZjJiCiDK3h/jWR
/v8BQOpSO7foFMoluuG09oh8X/5PV4UjZwIE8NL/CCacqRCXpF27C/8pWIxg
s0UhajXCilFGvfcneLtwfCbj6zWPa9+BxTzZvXfaHzP1rwq/jxHR6xiTrZPe
669dol2rJAH76pcPZldvUqVLZDEqdX6fqEjn9AfTwO3uMSLxZJvm0zRufgnr
bD/LGsLV1YdRTvsEPo5Y9UOz+6SEOZmUZozBQSircdQb8Mx+x+5yXs/DV5t0
8FgXzB3R2MWIMJS0B8qFnfMEHiUBxYd2XVIWycuVdZFzfow1H7d9T+qKezzr
oTB3T4JQPuYmP1C59SZ6ky5RIHMmIAg7JieHDjxB//VqCp4hApCTaeOoHCiI
6Zakih/wyCCUAg/LVY85FeG1T9klR0aUKubCa2/0ZUnDxBW8XL9WZ3RMQkv0
1kXNkNG0UbByGqxYQDHQ+mxocJhDhckuvPhPL1xyqftWJSadDZe6cX9Wp7gl
xL+/HcD8ofTz01RdavUdx+ACEQn6AZ9TwYK0GIL3UYvObGiGPnLz9vvQVM9B
CtDd7FNH+t1EZKMAL/uyxXtuZ360bigNdplCbiG0THEgV35b5FTZDbF6Mqa+
pp05x3Ts23vks7oYMZRQ54r5NNc9SbOlfOaUl6FoA5/3EfOeKMypLqjkpIwc
s0qjBwwr3GLm21Ekl0mmCapSfoEiWdXGGwvg9fx7rP8TBDMSjPbXzqX95Kq2
jskc0kANfrweetmSWoOwJ6xkNq6Q06nBNZSX3facpfA2f7dDJ/q7Su7bqAOt
+leIGh+sdAyR1qGHTRBO5wTmfSE+lxZTvgW/LcoxateMaZwTqOsmuzldfzlL
g9CAJJzBTkCq8PSZiQBgzsU46aEgIleGFYg+FFoxmWhaVshTQ9YmVlB920cE
T3GJiJcmWETHc6Yow2KLfBEvvxQ3Zvdgf1kfblGI+EtChJRHy84OOjrebY+E
19tsDituz3qgnA2VTzERlRGWNPBIukM0UY9r3vkgawQCgy7V26Jf+WrqYthJ
kO7/i4JnZKqqDW7NR21xjxXaatAwEVFgBd/vnAE4vDt37qJubSz0kmXQIjxB
7REqHvYsxTReb/flH651odXcpG7E0ZdnD8AWyfh/Um5QV3+S/WXELZRzl+ge
oANSFqLlrFoFQnv9GS8CwpIzuSY91p6fJI/e6hAAQMSSJIS97jZiQfF9vCWE
qT/fGij7MCB2+GFWY5MTlL+2JEV3fkvQby5L1l5mLbuuazG2+8z7O8BS20Ch
cj4LaB7SHC36eJArPEbHPlBBk0E78X/zqtj8f79A9vIbVfgfxBt95c2V44wv
HgCkwW1y+RowljDnTJ5uDjevJKq35gfpmrnvE2sqPUrN4Ff0PpbViJSqPd5V
ASqiC8bLSD4D99a2D66lZJJbt9Fb+zYIA5AA7bxPKIuy7dVyTq38zpKwEIdF
IFtW36on4warjjoKVzfh7ChW94o3geKToZMOD5wxJwV018KY1D3n/jIuRjp4
B12lj02HDIVP8rBJMBvFbyfTmG/eENOfEBhM6P7VckkyapPpE8mtoXLcNDr3
6rhab4tjmtBKav1c3gDZQ/fhZRDt3bAHojVHDhTjbuT0UoKF0dEtbzMAMmL+
ZvaV5JXxXcHe9pOtcP7DYyFvtc4/QxSb7OFitLjYNQindvzhAPyuabSkg7dc
f6VJxp6NoRpIbHHZG/LgpirK0cESZJgY2XA+gcYhkhi5XCxrksL+cj7mJAf8
LRrVFqqV+dcYhqBQTamFEQDJIOpp9zuMMTDq07e8fzGOHyaKI6G2GeRvSDXa
aFypBuuaYsgA7FES5c7wVeEa61DIexLxOje56tznjumDcFGrEMeX3GMa+IdL
TXiDRrVzCeT3R4D5EC501P2E9PzyVsTnUVFfoyIV0Gd30UsG0zlLnxqivqU7
9CMVnvYicG8khuNK7pgx1IxOl2JXfl1yCV2ifLeVsQNOPFcHmMZ04MZnQ+3T
s9cwWMupK9eGMEAwivB477tYNcUnHDjzSLJGCfhZq9AVrQMmecT0P+EzGRwI
VNWuzrPXI9fxk7RAwn3wtvceSBna2SoXNu8AFVDcRW4qfPey1pXnbglmaVRk
ZlhNPKq3zFO8eFrmENSNzRZEpJ3q3znRKr0onFu8O6K3Ye4iAm4G4RipWqwC
Pz6ZRe91HN+I75iBjyJOmzagJQzycv8yjPcMWFgJDx7tIzQPjbz21KJv7wgu
yWjKvi9/9nB+LwTmjGybaUcBvFeRJSVI/CC3o1w1wYiU5FQlf4Q4uZY4XNwL
uklPEs6MJ/sXXVZ/Tj8y/3OR+BhSllmgedFNcZxfLlYwU9lEpC0VStyUEYg2
vKG1DSGfYjkc+zwvBiBy/ePV/lG1dYTb6WzTCs12PgrtntGSNMlilPubb6XY
/TL8siWG2Eim6rLES3jb0nYguKIHqTjrYWqPy83Zosxzh/IUmrBm6AwFdaNK
FtbputgjbbJh6/G8cw8woL42myBreHDCZLEYF9SZpb8eWfP5XzG48M8G1g7R
X7njNamH71RH4OxdJfghnhdCQ/RqicKPs/OMhVWL7vsi2HRsoHnduPaObjjf
g3Vakbvy67WEyVdnmRHkwELrIO2U9xxRhvcDrf6ahjSQRUf+X5Q5z0dCkhSU
Z2Ax+tbIUp0D03DMlEk7UiGKwzM7c2w/TnoAwwhWgb6V2gEZqESzxgvIm9Oo
dHReCOhqn2mJXyWy0xCfe7lgQwp/bK+nN8tjpz18KPcxKu+CxMlbVL0606ot
D0lvX0w3A1qDPPfFGPScpTjCrZPYrHnD8Oui83Gud6zJGdqbSPvuM5YtpAMH
aSZp8e+krtbv90SqmQ9SHfkNsMdGfhNeH5i84x7lZi23ume1Hf7WQ0uvDN/3
qihj4IJYeOXv50FAPVNyLdh12Q8hNB3mpjZJapXpslcoSdF/n227nbRRHEyt
VCLmAHoXzPiuIlcc8RmObSGd6yV0ZEmQH1f/jjpABel9RpdihRIecFXYe8+N
ZucVUfCd7fKgOwon+06DZ7rES0E/8/JgPvy+3x/QR2YfkN+Xq5LWqDMu4rfQ
5dW1wiOFk7nJ/AZHy6EWlQlhDHI5wL3sNFZHJr1GPsqjMYEwr7FiEG6DHWIJ
AfwMXzi27YhLwU5Y1J4FJaQPIjQRll1Us6AowE54SWQWqj7K5+jJqsEhvMzP
F+tLd6/ChTBMWd68yQDXz3jKYx/7KaoeHVCgKKxFY2akq/vXredjYaKj0WAS
hLRv98quehegf7owyGplB531pKZtiO7/11NC+VFQp2JFjxyluyqKYLnEopUB
zcDQKmvxhjo/wCiCuBLy2eLU3cxefdCDyhS0r8zM06WC+yLx2ecm5WOTCL8i
KPtwWxiXkVF7zdAaepx0I9B4s8Nu4bMhl7Od3Z1YvSVqXDbQ8NqZ+RnzGl8d
dS99RATX0PQMEkoQN9hn9GXG8N5AOZgn6qeKhV6xGlSYzmGNPpOE1zTHkTMS
+wqud3EDHT+tOZfdXWBuPDUQ2oTLTQHUsYP2fP875ORGpur5fXWR/pDg71hi
y+ZEGJX4Dt68zbwyJdBKdQo5trXTa+NinzL01kHo9O3XNpBab0avSwlc44+j
hb0cdFfgMAIJ83/qiKJp1v9u5ppT34LUdX1PTAaTwpY8TA5QrOHDDJvvMJaJ
V5v7gKUTC+1FUN5GG/PRgfJBBvYlp0iVU0aZBIxfRfnuUk2NZVBmOHyYRVTK
Heec9d7yHw2XnO8oKa16VVlZBYK6BkRG+emIx732Sdq9hu7P8XDHjw+uYBQT
3eSfefCtzwtiEanYyeJw4vC28jYhQs77vLC55UBu8JRcqfCh/GIsG6mp0p6y
mp9dggrbShesAGzhEnDTDuVsceC8gtnJ7s9/OjHsJjbEQDqZP3xYiPDMkK3Z
ayasDqbjJQKEplwfH0dxtP14J2uOpGlBKcgqdsgR0hwSV8fcCYrl7qzLHZcw
XzKwb5Phf2NujOFTpPb8vhmv84en7Epa6cKGr8q1W0IVfKXIXQ8ruJNRYZzc
QtImyXCMtoX1T0ifJTRTu34d9KgZjxECbsEz3UruXI2WjE53pg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "t4xPJbmEH6v4SVL0gN6FMeKrn4IhP8uxgDEXixmWFrfkRmUmHah0woCI0NWn4jNi29PHRr8qC3E+56ObAVSYSIpu2luY1Ux8HxJTmEZp8dfWiQKOAKoquE/rRpOs7kTiASgRERfy/4yFwiIwBiIeSiYycsrshs/YcSPLGlUvkeFONkowA1F3QkwXAeAdMdMqD0IZHCYUiyRDun/uIWwwqKpaY0MedDAF1dXVq3jdOllXt3gISiYilu2vx6HxDBBs4Whkk1V7iEc2K2J8NNlxXSy8+Hhk7DAOp41IwHPNGCAfyVS+G00R4zjqJgcrlql5z5h7QEiiZr80KC3kmWJRiJJY5+aR5FKYm8lG12qxF+CfBA3320/6tR3UmZlXZvNTIxGDAUdFiXAGn3l9vNU8LbQ5M2tUmhtzd1pqXGqtsVYoWwFqLIUlG7yaq8OI4xnPTiw0H15jhYsywvjko4M1ggH9PYfnBPOW9Ru2U/LM5/dY3fC1zJF/25ccMOgzBXgZi77W9wLuVlttVRM3zqhfn0ubEWFVUvKKpgg6sHAW6KT+tpknkDx1aE0lrEg71Gh3ITQfHNl7CaIe4NzRVLmUWQ/PXaN/y783vEXq9xUZYPqW7rcNeeHipOyqYw3mgxXjNHLsQ6HOu7IdYXK8FLrUHLWrvb/LXaTwy/4gcXd8EeZdLuPimKyHktJLPLgq4Yo/6ATJP27IbKi+E1iE700wBPhwlOnjN48HeBzyh6wZMxzZzoh2gKMn0Bm4NwKUDw3WT6N8hFUb1VyMxo7ZBXPKt81B2Hw2clUtzenYVvLcoZrN4Nt15X7NKoeI+0TSUmXkALZ+1VQJZ1J0YJWr7fuzI+89cWeHU5/6kxhO/KW1EbjbFxFE4QvNfuqg3WWyadIuEQ80MOKaRuDB6sfddULsIHoFkcW+3aIm1yPnCqtrmv2Lnz+mteEGgXc30RcfCBhYUdCEcn+eXhBGX1vgfD7gMlvD2GMW3mJ0MqXXt+Wr1vtxe2ute5oBFvwAiC8l2Jbh"
`endif