// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WMPisgDWo+uD8Dcu/jWLE0ZGchVw0RIBmVtrQzJ5AtDg4L3izK/TAeHknlvS
5119XkmNnzzGGXoRADJ/0aA0Qv/wuyhghcUq6RVk71nOuB+LiqIl4TyW48n2
RsxY3F+xMhx88fBQ2Q7pZ/offWHXgMUBmKKtOMvs8N2ZGToan1BKcp8TzcbM
rB2jC0Ig37hg0B+2zbMuu+Fioqo0gOjuz+O10XMDYrNIJU/4LjHQnuvklK82
y5u0KlV9wMU0j0ayDgTGqcLkhUsVXJ8Lh5YfBEofwDgHojIY48X+tylQ3InW
b4tIhYL7oH5umg8wUKeL/aUSNrQ7b+6oAJc+adt93w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Y3GotMuz7swajprIYc78s94nJJLLE7gOJXLqScZ7JwbnqS7I1B0wJV+Mx4ll
z796RUS8KyhJZzGZ14SWdRgkaN9lKVGjHu+ABToI2O4sd9YZly1RDqA0gRmJ
3AzkR6KyXcjZ1b1PjK52JRNSxmtqmIIVXOcVzfIM3OahiHggxRAqE11cu2IA
oTPihwFfRRGtiWbXVVH45sh7g8e/ZQHU+EX5CoP3gXPJSAIL/VAG3HRxgIj2
BJjAKvW3k0qyZxN3hzZ5iZ8UM7TX7EPgdkv87tvbI13+VcA86VyFkMwKf3Ls
JSSJUvqYzJnn2mLzS8OML06iyhrbr3cSUTpqV+iBkw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aDU9qBSZzcwDCcocg3ubIuN6zcfFkynKPzmZ7AiQ7734qamy6UYOC5/YlE38
VgUiyM7L3qV9WWHJb44xlsGTA+rL8L6R3v/d23YnhMy50iA86P24Pz6XRYg0
S7S9j7RltyVfN0FlcdhQFNMFZqMMw208Tv8I9nsUIoBK4geKUj+pmy0NNGdI
0VMv4Ir9CW/cM1imI6QesJ8aUu4bsubTSggEKW0aNrI5F1iU3+jHsi3PX1Tx
EddBYk2uEz2h+egl4ZxV8i1EPo1QutRuTAsIsaIc7nOKbMFJ7EDPKwrQFdiL
jxOad7UA+ihzcHj780nKN9VDHWCnxybR3CDiQ2nnDg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aCZVdOan9cKUPr/kXj+gW1PqqNN3AHMKsEqqcrGnkatn08cimk+80PBXfRzm
eXX+i87BWXz1tDgEJdyzitryPUn2MiVPx8BC58FHTLhWJ1Wx4JMrCdlVsfa8
7FZC9ofhtSWezAJlHtpRiVdP7U1AqGwEg1Bb4Pm47Wyw68zi0Hc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EoLXIKHj4o03FdLn5kuYWYHBnPluUxo9YDg60+UHT1fqkUwSMCZN4xr0et1G
91CTM1ZsvOTk6nvhoyn5/hiEpbgAUeqj5Pi5Jgzy4O0xS5n28TQy8hVfKlto
AaRkDrS/GtxIe3I9l4diooZOaIiOvoutRZThw0vJuT2RGOXMUM4g/zCAfcj8
PTepwUSwhJnMcWBGu3SN213K73vyp8xK1xDGsD2JSqunjVc7zoSN4Ceqc/N+
qEbz9HHa7iNaYp48WvXLJsFHrp+26LbgrbHCaZcRNGoIBIAkALJ1e61PM468
t4/XM7D6dRtwWOn3g5AuprKjUSxNc70ZI4982rtdPK5KE9lG9/YuxWbNP51M
d110Pu1PwkhuAN5zXH87YRg+sssfnPnLhJff+9+ur1ZHRuEUsQ6zRB73Fpmf
IPjii7eW7MLt55EUoGFeNTYZSVcznk6e9Qsu+Iso/6zlwHjmGBV3froDm1YX
DentdUdu4FnFAUziZgYEAPs6O1RjbDa+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cbGPaSrgEVWWaqUj5bSLWLMfDoRplpQxxS24rpTSLeW1ARWAjExmF6NxyZ48
Zorj3sVu/qKXdImaqZRGTfF7mnN8hfH8ZXPQGjWeJSRRo6KaP8ggItorpH8t
cfkft3l7HwaiZN6v6QKvwYnGqhshBJv1HR4GKggBQ56hBuQCliY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R//vtPXPhb2VvvOx+tB3ePYHwhBgU6iPLXjbIkl58MOLDZ8lW+M8TtYqkIdF
5+RQTTkd9va1FCWvlbV//yalsv/evHw1Mm7UFYC3070X15duCEjIzI+rg+PU
HkPXI3QheM2NhpHIoYCcxXWlsvWhGZR5+Bs6nDSjpAcHXgHkUog=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16912)
`pragma protect data_block
L42oksmiSV2Nd7oHEyUoNgpLg01zqZZOn7Z3Juw646zAel4rDWjIOcq4SbEd
egf2Nr/m7PJ5gUJH+x1hUqr4gj3+E0dFU+q0xoxhx11LMK6PXje+qw15U4AB
1C1GnnGpJBQG3bL8VQ6Ny9LghD5dJJPl9fiVhFTar3u2SEuRM8lLOHSwke/F
JzJ9ZQ05qui8vbWX2kIlT1C5yFxDSTd9DZb7BjK8ES56c6YVs3h3nXJSFMzf
gh1HpyVHyb2O8U1Ns6I5fblfbYTw3sN7gYBIhle0cTytCpFbC1lV+MxYuOZg
EdEsvI9zGkRBTdPq3InrhY1erDxbXtNr7/998odD2oQHIUNxVAFVRloxjJv6
GfvytORvZabAE6tFqDx8Nd3LiGAo4J6o3z9MxQVQ5GNf9dG6fo1tgCZoDoIm
Ck9L5Tr7TENpoof9PatEg46NYINBNf0t6nWQU3IifnY1yWdq4LodEJPJmQKt
Kk3SDQvP65fwUUBXpY/7pHlOAEHK8ZSJOIJ1UDcehGEIYKr13LwPe3OJzUp4
7kyUVamxMhYHcNdXWX8qCgLv+twpcqqOkUOOlh0jsjblezJO9rWhM/pmMBy6
2gJ0H6MY4IXrYlGnNPdx8NvygeKqUJhlHcQ3mmTQLwp5PdvwaRBkYD/BboYK
kDSzi+8DQ0ADQbOTA00JECA7/+FazgYGCs2IpPa+uZDZeWmrjG2CMUSygsMc
MUo1HspLERsvnXlB844LR4H3U1jBa2XqA6F2rZS48hjv9HDrE2L1GyeOXVSM
H/mmKcD/Iy6uq0/bmWeEWfa+SvndR5Id5aNTon5RMnWBzZAJpW8laakpHrKA
pXRIfGo3HyCPcdLPDHqPMFN+m/UHlQoS/C8+zrmVPdleGaUGYZxikknZaMgn
YYR4Q0kfgWaMrfzyNNvO+T+Pyqi+3B6lTLRc1pWC+DqONd95Gfx1GK0NGo+b
t1ZBid+l9l46w9ggUHpuZrTMBPUBwASgjPShMUnNB5fnJ1LfRy8k0kX0PTCT
8tiIYxsP+28Ojp+rKsk4RP8LidRZXixQa5qlGFQAVVWZ7XrzWsazzVjwUpyr
KP4vnDc+Y08j9xBx705jO3CiWzfT9DMN9KX5sdDWaBhec9M+M9jNbP8tyyLI
m4tz1edRbNWpSkRdfjPz97tXaJpnQjQ9zeiuaQO7ORf5goEyvNuaaIsC14h8
0mWNeU4jkuFynRrOjB2CFG+MO2b2U/B3QFP8xKjOJRqxNXz6XXWsHMFiIx7a
Bi31LPhUjOnFGulJVxCjTe+KYKCuAeegHPw2wjRlcoDOd8PQ6ZsLJAXmTx5Z
P/Hw6IuS9lJPZJA8gywLDvK/HBU6m2rzKeDCkv6qCrjjjxygXFpz85SEp7fE
EyBSHQtifSkErhEZjpkoizZ02kzARJ0hFHJGjbprd65UOqGaQifvUbQheJ4d
/9ZaFNt88EkD/M/vouzhiv3bqWcVi9e6Dfq6ozZaO2TyoKnDAl1FAN9R8MjL
80YXGLBOmWE0nVwMET+t/i+dZZJgvGyrtKmr+IuixRsMS15UO213ZbvjkykB
8S+jDEQakDIxXuj9ZnkjaUqNV0AnhgviGpfjiUZK/GGJsljl485hlCGiOABR
uOpWb0Wtzua5l96gkVwv3RWQQtVhZjY85eFkp8CMJ7rMTmrwLtq4eeMvEE32
/mK61uxtUsvi820NfZHc4fIdcuEbWQLtR3p0dZTQChAuUgjtOt4jC/w58SbK
0BGwQaW6mXw8/VQUobPRWf6yhGTye2w4YDvTTH+mPkkxVz9BAuktf7ve3Uck
L348sEEZOg8/Gg6UjgfsKpmxFQ28xbp+j5mpGN/ngwf0xWML6WOejP3qdSIL
4h72SER3YIGsHoMTx9n4aJQi28WJ3GfV2kDX/h5bD9V+stD4PzusKB2+gRTf
q2sUPYIh/6U50z79Qyk8oP3MFMWChKn1ClU7dv7IjqgSCemSrSjIt8DVE3M8
/T+X/Oy+i2KWfpnoXBnMb+VWkTSKkUtX4fa7+3AHeHIZvJzdXRNWR8y8X88F
8lp9m9HpXu7U44ARwpTxEeeQOQDdCXy63sntMRNPyKnOI7fZ7s/7ILKL3PT7
7/tfkCaV0QVZz2HLER2Q0PX6G4jMqtGPefGN/Sn80RHgMmKN7LLbJj0m7JBG
4y0Y4mNHKl0R9DHRh5kkkhXKvR0NEjqiQx0b2rVsCYnEwKHTUANhC7HyuFl/
VNtm+h5DuBBsO1GksDCcl3SRCMHDNVz6bFDyVb+8IUrBSvSS2t96Jcrb/vjh
Nls4dNoIdNdFOGIXCZNTSz+8f/k9AFqmIVaZddcEOSj2hZHb/h+lJDRV9Ogr
UunGUATKENS4JagRLQzjBIdLDvFsEhqtauxgv8Zo4/DOFryU5GQa5X6V1UrJ
qjDf4e25ZbeWwYQez/q46j1VJM8yhNGkJYya/WWyOhmKdYwnpA2F8SVA6NPH
jpF0MAU9t15tJNnOigw42o8iTJ85sw/Z5Yv03x+DBqEtRuxi1ncFBXnbndS7
JoKK2jjOsbICrTtfcA0UNeNVu9e90feY85UhIjY3flKebCYBcDXMcvam+U8t
oWJyC/PqF2AdfzHVSu+uHTf96wUGYFVk88d2kB8+dcRSjmK3/pChsv1Hsj/i
/Z8Zc7TriqHNy9KMB2I6HQ2VoZVSIBuNS9ahFIkggpGJdLZKXYGf2IdGdJGC
ZJihnloR9Zj8M1x93qPMn7HFERMn5+A5KOZuhUhuA/Wt7jDT0Wr8Hbfg0YDu
cqwrRt1mXAIv5DxBMGOcnXALRAgQYD41bvE6kPdoXktrm3VYXvYdvLu1Gw5Z
o7WN26vgWa8ZbvYpDL94ncYSaDo3CJ0GLHhkSwtu+7npSU0QTeDA7AhgxgqL
T5TiHdjjOiNWEx+z0Tc3jc69E6G3DchskJTrOYz124OQtz+PNRCsTwhWm32U
iF1OUFacyVrHWjeodHgfX80IilBmfH5jTI3YykzX3mCZvPBr7EgLwQQ8pfPv
SNj13gOFjdS+pzGgKfQWk4mILgYdHxF7JtKhAJ+wCsIr/Z6IniZm/lBI/BfN
zzXHGb2Ew2P5+vIzf5Hq0RtU3leaMXLoN4WtY3WqdTZv3FGavv0vvGQwk8Ag
NVYJbdA5NKctBZ+U6PfUGWRcYF1vqdJmtjFQ18hvvzIJPnEn/mLvrlRWSWYa
GDLvYVXjA8W/47qlQsNNki4ENdxDjdJlIuBYrzWfljGv7u2Js87SeCDOMuqR
6fuFwFFvGrVXnliGcEu2omKAAoZuyx+jC85bTPq141nlYeep0FKJ4ijT+MAp
t7V/a3JpNA3KMMedc1u9cBkilYnviVCNEZJhT9fJ/EnMqUPd+14LsJxkfTeo
t31fm7hMZ+kaouG5pdZpobT13DNafpgughwX1m1wY+EM6v56pk5Ewr3APhLk
jBxq550PEyTIk2STJCugghnnBy/zcz5ZYtLk/7Umb2Ot5kpVxpy8WpJmGP/6
q6btfJ+OEbrAsXv05tw/QUz+HX3eakLPlFyo0YPNDqlUhdmnYBrMK1bMReeV
yRYltgJVQO+wl3M9f/zprsd4DPojwfO4/ZWKtMptZ4jUWtJo72oU+M4Ui3fo
WmHm5dTBMTMWZyKW5eY8sm02mDB79dS4D3EwKsMWjYKj/UGUAv6C4jX1+o+O
YzwTXgYGVfEhtDMBMXbjoFbf5iA/5umQL18+KYZnC10NQGcYGI258/shhRnZ
m3dERPSw740SdkUDxV8yHprsfOzZWKe2qO5JBECGxxYJz+BienJq+yDtR8Fk
m3P7Ix5qILb+O3c1Fdop2jZGWdBmst6FtqfNHpHFUGWzVxbQdsFctpAJrRoX
cMOU3m6QqT04gp2/Q8nsQ/ACzE4s4XivmByjfbR+Y+M5lLGdw2wne8GDW9j/
rqYso0svxo6zTAFfG/ZMjSmx+q/rIPrpd/MeDUKDft/MIfCbENB4OzptVkp4
YpesRaWiaJa13y2NFvrai4Bx0WvGyUxcRL57rrq14tLCYXexI/9lcSNJgqGk
v9qL9/nEMP4H1J76phxVb2UesmnrqIgjbsaza4U6RO1DxgX+g7R1tvYKax/c
/FG3V7ucTxMkPW7v3HBjaBWfnomDXP2tBfi4gRK05p+9T3yJYGWAtoo567Zw
50beGszULUBdOO6Kf88qUNPhGI/ZWuAdIcEZ9wWjfzLohK7wzmTOXkKuxjM1
qB1CecG5KQh5BraeiO0YA088oz7IB7leAZS9Cy7NcdLBePH5bxG7IHXW6gzw
qqT6HcGsSJuTyQ23gcgF6sRNSTi7oNJwgFJv7KmgNWR44yMqFfdIE+/Am4cL
EuRI6qI1bVvltO/x//gwV3CqaOHhxhqHzssBE0MS8cAleEmBfGZ4ZYwg8XBm
OUxmScke6ImbKdFELxtEDrWe+045kko7YvhCEjN7bR/h1ieb97C9Ad7X+dVu
uHQG/QR/zf+0dJDjrAR64C0Ij8YqR2mQsOqKf9nXU1Q4ymq9T6lAy5D18/Jz
EV2eIbJL21ueOig/HkXVPk+sxvciUBIYIP0+KHhGjbOVAn4/Z1ZbMAEw4vdN
QoGYREnpwS4DIcriUZb4euBBzXvhTo/IAoQtyr2+DuPBhw8eIY4wyCMnuLW/
+GRvkBCVrriUL2wzcbkEht0bojcFCT7Qxbe64173XRrGmaIQ0Udg1BPKe7ps
5Y4T+Vlmm+K0ZQWKuh+BvLx4FiBS5IIVy8S0/1Nv/pCCnp4QdqPsnJoj5ZJy
PMJXxPdqUmgE2npSwiZfLGBCiIIb1Mh/E8PjUsMVvZAhBCHY3vrsYEabmDtF
BcdZK2mVjE5gY8Mdr7ri1e7UAjHuzDj1DTHKYrgHI69tyrX9yGK0J48FGZyX
FEy5lqmuFyCY23BLtf6HBKGpb4a2NAmA0i06vgF+Ad3kZZOi1qR3QzHfBBL6
hMcov6bB3UX2evQ/unuEeeYvmmSARmfC1X5vnUdumDIb/HJnpl0Y8dX4ToNT
cDGIJxE2HMnQ2vVHmdwHOSYzLYWpeSzdsuf7JSHiAbvTBt9apraL+NcvvE/Q
6L/u+C9hMbVv57kqWcPF9iN7OgXgexSvNtCmI3xdIwJl6JFq1YIIgUCVXBuw
OFZNY7pyouDGPwbz0Fy7o52AuwaQQFZlMo66A+xKPJGqQrTnamsLkhSmJ2FA
KuJr+L4YF+U9ZLadOuJEqSeDjVzfy3plKkoEl+T7z3vEsqa+ZNKGwFSccXc9
pWNeNhBIswS91pJZYeHgEJ9t0xvVVHHm1zsED/VcelrCGWUl57vqHZ/ufK4P
aZV8UKh7AstritYndsjHhuvJE5pa0Dc9zIxgtP0tTMyZ4uvaTVd5ocSDicOD
h8iY1kjpu7QBDo+S9i3XIGPC0I5OPSDV5TdphLg3rKA50Djrt1kZ+tRJyF3+
XaQndyaGlpAWF1f760TAaCs6yPTUbIKCoMm1L/vt9Mzid4Z/5MEazdD1gVqD
tbiy4zmLoLn7cFtMxlfU6+Z8uE2nGSDRf3zqh8cXNjieLFN1o31hXO27K2pR
s86otCqL9UVKA8RAUBQmOutZ8KsA59xpjXHFF/X9hSQv0CRlPRmoK/pY84yp
Z+fxf+Rkr+3AWtGkDxZ8JXDxvCHsWW7P6TuvuMacv1SeDjAnPw+0Vee9czkb
Y/P0xNCk+E9emcp2MZn1dNXfo0qxRG/oTKH9PP/VMfVh4z2BS0lc0xe8ctAZ
ja0qPibIMtLJlGkCYgfviCHd9PlwS5+ca1cexQe6EFo2E34jRsqFUKSO8+Zo
UFXZkWBFXPVHmk9NWwDevK6rKmuXP+1dOXkODxeGQN7ANPRqDnZBTVPBUDIP
fiEa2So1cM64ulRcytaGv6T6dMeyTT04FxJvfbD1QqVNe/jorFRylDCISGIX
2fcElhyJMIT0HtyySRdrXf78Xi71/jcH5PxBLpbbjEgG04WSYHqs5bvhEfPI
sM/fRO2OT3RqZhyCZk+kGF7xs8CkFthRQTlhx3L7ps2DN+t4CgTG8tRByA/Z
pX82/+s5UdzaTRzf4myflVG7095iNIcOwa8sXYqeL2yDHe6b4UOdaKqRcGUn
lHYCbdY11yGCxixyk7SLJZ3tDZ6dIx3S5dTmZQnQvgkeeHPjmXuEJPC3LGce
BQsPC2gR6EYJIDioED1L5y4yiEt1I7+YqLudWLSjnxqcGdMgY0enN0eZw9Xk
h7Zek9SRz3dJpkkPH4+loWqa7Z3ECECY9VTcRa14QkZ5/KzTi4WFIFdE00Ji
IvclwQ8ZXnRaH6xvl2jGoc9ePkd0Tz+QN/k1PSid0Ho0DKXIAE+GDqK3/xil
+/YLX/cBLtFhobbbjA5fKBeI8XCpZfadQyrQzMD/9ubTkBrZG3jZKjYVBrfa
HSciJQCHYPiqcnT9Bckg013KzxjIWyYoOrc2SzpLk/pVZzbYDPRMF2Xghlph
ZG6jBHB4OglyvioOexBKpyJX8XdvXxvEYu55r/qFZby9czK01dzEtwm2HzUh
3DM1xncvfQHTfFLaKj10TnvnFreP+gfJcb3vYB6V3xTFS6hTaPbKPQFMh+nG
GQ57rWibe98Qdbb8tEDScPX5YnFPNF8gHdofZQVIySjIYtDN635Qdj0WC3oS
wYbY3cUmZdVH8wJIE+KdXKq5nE2TJ9ua+U9csgxKINV14ZLAOUTqxFGQTH6h
vrLF6rFXs7OATZb2mcDl3n1kK2HLcuBdjm0kjJD2hqp2MBch6v/422Re2Bb9
njDj2i622P4WWp6A4iHFTidb2TAIGFlLZIhilgFjweriOsAHXYd9wMtjX1EF
LSw/Zn5lydTaJH/JDiO9dZkw7V7zASxTAgt47UoDuhuAyvVJ82DL+dmSuQeu
/qmNZgTJvvl4DMcxZ7gX5SxsmJokcjO4oZgIIpsjgAcjsZ8cMDWZ5lWaTmpq
CWVvy45TK+Sf+STsQcmDkkAP6uIuCqzpezvJIpT6HFtnA6ssYxSj8Yoioy6L
Ld1jhi67qLGT/J9o4NYXtGBnAohPOJNnzHjNHIniee/dy6CmSnpVNzLoCJ/k
CNn8FJ5LC7/g+X5986ImX0I6yuFHNSW5ED7yNmwrQpDmd3qAAm8CpubbxSt3
8Vm2lCjnHj5hzA+1hV/b7Eba7HJCK0zyzQVf3xDd1CdxcQbhf7hImsjs0DEi
IyKVffzQrXz3zVkhWXRuMNvDXeW2jf0kE0bnmTWXlyMiYfSivlB8ls06Vr1F
DA8ZzSgbkrOuFAaWzBUk9qWEvnLpPceKu5VJt6B/A/6FAuD8UhJXunY0X+VK
RT1E30LWBBeLQuEhJv6p6Ly4esOyE4JCU686mdKJfHUvQaJtWQ7LFQxU7WPk
u5+ypAS10M07vt4covpkBbYJkXriQ+iz84GB8LtavIyMxGSGHRj43lKF+aKq
QzrqK/HfjlRs1DwfNYzGeTymYfp/vppAAtygJw1mHyKrb7Zc7GtDG5nRuRR9
H1FTWER0IPFp+mX9sGWKlZqdnfHzlkz5FbiASyGKadOvyem4ovH7LKgmcLMU
S9006gvZm6idYfDdYR6nfxH3v7IV+83hC3kMe5XPUkJt3oHx35Ucd0uA+Y30
3hjxwP7GCM/t54cCPhHFWFLnOO1sryTrK+Qn3Wq9IB0+UWtd7/0vQHSQlNVW
LZ3GnVQjkdmwYKeYMoCT8I7H1PZfvDEFmIuxspK9CsjHxIgzEgkl1jsJ739/
v19dIhzRrFlYEFK00AynKGQ9TJHRBR+Y2KDDFfrwfzibVf5+5A46hN1NkR1n
RtXPJcC/LSE/85mayz0vWWNaQTH7mVvkqudSshNpA+W8OCUI2Xrk1zYVnrYK
PRVdQPEUIb6gskAgZWGNajpPThvqRIqOLdDXApUU6yXxmKXX6LXzi2aQGUPu
pyfYv6rQyaqfxRAbQSkGlplquVk9pqDHNtOtEF2T3cf+7NiTQuu588EdCuY5
IGRspBJo/u1bHPxkkfsKo9Du+uRXHXWcCZTP2H7FX9cr8by/H/j5fDbgrHif
ECUwklFDEQHN9+qJHmq7K67FEGoPriryxDSHatqM/OrVH/qlt07biV43bA7F
Jl5X0esVDQGryTDfZjEw8QtK5hILMZ2/aFYJozt+GZcLvQr+ln6aXH5b+3c7
25vZ/O4yiNMXAisgD+tmUJncUSz4aM54jYzlZ4EiLQQU0rhM6Ntg3cxnU8Rl
lif5UOQOTB3/2nFFRFcTGiRDscKigJDbv0NWo41mECsfOOrljD+rPKTCVWsR
eDjV6aftTEfB/SvHG1z7l6mM9e58OUPiuRkt7VHjcMxtfCnDeoVZepWadJVe
Wsoc3/C643H++M0FXP3fdw3+ICBqgL5uLFGI14pKH9Hq7eRv115/tEbo1Tap
bhRti6KlsqteUyubqHv56ILZdiednwx4FJy75GQLpT0Bs4gVNLCPLxNO5PPn
NcAeGyqDuIy76QRiuI7YfcAKMbCh03gNtvMpol6G8RoGMV2VLZEPGOG3BFKn
IQ36EpJTowA4ulH9F2AE1sMgCWw40dXZDo7Nb8QhKOBjTZt3U0TrS9XT8X58
C3WzI8SRqtyCBbaaUW1Ws0VumEBphDxsqchqh4wUfXgBNJwim4wVMQSu8MKu
bxMh6Df/Dc1P1kg1oClt0QCGPdEEMEESPfujaiYbmqS+thPPWfK0aq6BDKGy
XTX4lJ4yQESMIZyfWqD/EFCt84bjGzYwR5SnqegOJetgBdi7bly/J6ToKDEz
/TD3JnmEAoq2eKB1LDwM1oXljFtbEhpjqxzwTGAwZmH3rb3Uy04Wd/4yry+s
GemvE9/HwmLy+k6weacCkxYmLf+IEtlhp2IQG4g1hit52cr8AASFCkjGLSXB
aYs8vmZkNzU+O5fcf8USB2DqEuCRnVHHfhdU3XdjGmDv4Tbd8ahkQqeCycvu
sZmGq8ovBuxC6K8tLYk8+RAQutQCJU26CIdcy35Q5JFlAa19Xi7anSxhUMhz
XOqD4ELN2x9TomAWU73hp6tSpqIjQ1GDxPRIZXGaA50M7SZFYnfY1+npV3mp
n6JhlGbC4Ksh6tEph9yYq3P8/U0JxOhlFpN9nEU22a+f0iHHLZFa1coKFqUw
qKc+dPDE2uuoCz66uublPAOpM2RYc5Vm/jHrBfAMQ9mjvxG6NuqWbACvp36f
Sg+pgYmK4TAlBSlQo47robWZqq5ymLq3Gf8PfjY5cyqH0BNEOLVSr/ghujSK
s30iJ7M7Bzr/OdG6VbDEXha9DZq+c/dgpC/BV35SkEtUm3NeO1gqw/DqMcSI
kQcZPe4Kt6SXE26yarKBRS8UyqjuPypPchhBpMYHFheimo1RpOe8+kRBAj42
YO6LaXM8hca1MUkzceVF3QudvfQYYzPKeekUp4zUK9wWWSTXPN3eivflAlMz
AG8jmccsAEKTkgQQgau0QVjJaYAjoEjWz358AMb4Xn32X6NfQwGZKCSc+gnQ
M4A5tqLigZHGaXlOxkiDgyNACNLyYJS/KySzME7PAiI0f9xcS8Qj0MEokB11
utwqop5uXiLYXWNyTe2MLj8lnTkDmcL4Lxua8+oEkGSK4X92aYxn5XTBdpf8
aSy/YneIcs3GtSc5Cj7Fq72/RJfDUZAB12BRCk3vok4dn+iDtmTqPwgtLHFC
L9P/qCNDWn9ATTza/WVox5T6FChanVX9hbklKSLYBvVglP0n3EfFVWo2pMYs
BddQ0EBD/ZeYmkOR2HWKR8BAhT3RWR8BVBZ8F1Mv6uTZrPy49/B9NJwYKeS1
F1+SlZpg8gcIdays+qit22uoHz9aKnmGYf6tcCJiFaBLRC6ALIzIeNPIVWen
Do1+er+GBIMQKX2DP8ALhClIL5QfhDqA/u2AMYyZJWYX8PR33V+jUUwwtNOG
stQC5oXGu7MbjSsA23vxeZy+xb7BNiZETwCpdmXPPJOPLEU1P5IZ/4MWnj0Q
VOY3UeZYqwafRzP+z+zJVS+hdek75QfCJ9G5FTyMVGP+Ych0wn/u406Vq/Yp
3/6qQbidJbuZTqq8RYXBLlIZqWZ7mF5+RH0m8fTlERLm68cotTPGwucLS8lG
yKwknbJRHUEJu1u+nF8laPl+UlgBi4QrXm/tomvKqp6KYH9GnaaPY9yHg/DZ
q/c2atN0NuLbrSzzZgGcEmwAiUAQfBgakGocfDnGOGVhtgzvjQh7RE8e2ziO
X8d0Q2VzlbYdQyayRnp9bk9xghijx08fmFUHwvtSvdvcyZthrOaykVt4KChb
n8rXvxKZgD9NVRIZ1AN98ulI1TZ05k8uouDUVkuUzy4NFVsMn7ZFuBM54wZj
fTcxdob/rCeITzveiQHchD+mzbCkQk7IDKnBxcAzX72rjbRxLsVqNfGxvqLG
jzl/TDoM1EnKkQz2oBFXzja5Tf16cQDOzumKE1+l8bP5DCeIiO24lChSf4MX
Dq2EQIobZHcFOaBKZvmoQzwSMKmU3yBYEhQ1KXZN+IL5iqyeKSqqUVJlI6t5
cDBpOg7lgBpXKt5nq4W8pusqpaerJlCz48PM+sJUeZJUlbW8bBrWSowXw6MS
mONgjCKMC62QxQhTmYceHzYdBupfttaw9VIw2mMXpVdQl6DP0Vj/pw+2wG1G
tKfc9K4DSMOQsbjco1/SLnjdQRMw2JDJnlD6N/0kemfXvIb5L8yw3Wt9o1R1
SazCPE/OZrGWps5V8O7lrs7LR+wa/NDptRvDqNmbHIyY0rRk2hHc8DGAjcvj
dtO4GXmpZQnC6aSeaVDM74iBbRGZSeLTbyJnSLJlNuP7/d9XitOADXMEZcKD
bPZRf5HuZ2KxMKqstp69ACR8lXCRWoqnd8pKEPSzDUluaxTozuTzT/yTVmDd
EQeVmGb1y8B5YOlUrU7mLpJPUXz471jJXFXe0ye9b9eqCjgOt8bm+naftntj
L+jzgmY21VggFZqop4vY84Ou4n8JzA2uk+HxRrwSTiNT6JHNoMrnTEt35xd8
m++aQ3t0fK7L/eXSbj1vMBNXinaM1irEh5An2gweR4yF7wIik6TW6tOwiKwS
U2O2uvMC6ykBvzR9JX85TU9yNBvmIHxruyxyspp2gSZCqUBeThfXAqIpbGRu
CRmajRURHRUhO29+BSGPqk3JXEWhgaV4ZHbkjrJk9Gt0bdUDvOY8qQ4eLjm9
gvyvgfaLOrk3H6LHZ1uYAaElo3iipcHZTKZPK3yjbgnZgeQ2Q/XWysE2Zu/q
9B7OYtmuJmuNJKkif9AjXKcV+T0z1UfXo45vZPnHJeKCyqPzUgieu1u0oC+g
8kT5apo8obgUURx/Xm37heayQ2FFK/9Y/gFlb7m8kwIUwZCXBjjmzl719kYu
ldoIR8CmwEs6mJhsRtLt1Du3cj8eKXHv25yMfjdINPMQdEaqBIvBgcRtWLKf
KXloTpv7MKijnwb6JiP+fXcgC7/jdeL+dHLENflH3/urMzmpP+HHDHtPJ7ad
NqWr0SdHE8jGo/F8g+KRIHCMPqTL0ZVbSGwlwOF0JcX69RjgvklkKLANk/cs
KkRqnwGr1w5Si/IlU76mRxmm7x/BVAQlIfiR/lff2s39MYl1+OOPKeOC4sPf
TOWSGduxumT7MZWdgrOG2DYiW1YtPi+5/Cv0E1mBEmP7rXuUprGYZOIGsN9o
hZEBiwLmlcEHHrhCLXJHhy3KMrYAGjOedIukjlS9RkM6nTTezdot/enX1q0Z
A8jzDhOOIcjwVFL2SjWvHNmqyS0P20Z97v3GetajDaAey4Xhfcxprv6zMqN/
Fb/O0qGiViaBh+ct24Vu3gA3N2epJZvXhaQJmDYWzTRQyZe8D38iMEhB6Q04
Mz3tftsVLhV+HHnaToxAqdUCBhk3aFlRbA8pGy4e4DIyJmINs3GJeuTTYag3
P81JmTWuquhKW/X2W/whED+02bXQyKEr6cTtipA23Fnn+3ZsTVHr0bK+zxnd
DnPxBZ0Yh8j0fSjlM2LXDI5xnhmuHWAIxEVi+I4MFW/PWRcXGdVPz4s38A0c
bf0Q51nhTT3XQ4g88gqzgT9QDp2DlMD7ER2cwe91UZLGK3Csiie5NTxwiSKa
wzSQPDXbKnFZbV2Wf1qnwR5BJXK8Cd9CkgG9WJCPDYGun1Tj7Y39dhvUhl8N
tICHKvensoNsDktQnWGkB5qDahaCOj83WUiyg20zcL5Pg0viaXEEoDHfarYj
VqnGoduA9OapehoCgFPL0Y4jlK6Zfau+TaZGbxfQvpIZ/Nz6nUvRQwRrODLS
PzHo86DQYhGV1Lcei1d7jxExiPEK9i0483l/Zg4IPuoSMAte2PBj8OU2KvHY
A7xOmdnTkCm03T/nSv+ZQU7OB0IqnFiAEQbwYwfU47UtOALTIr1RKGoN5XB2
XVR0maRv0C0/6eESA3RDsw8tuEKHz1QlgrodOEV1dkOeXmJuYPbUQoj9Al/j
0LZxYa7NJAgD6lhg1GugO8erqyJ2O2IauAaE9Mh1BIVywT1Cl0PT2mN5hB+P
hiM+iJthW55CQy0Mq0cNKPdcybUl1Osoxc3KumetMbbWriL1Us5XR3+sRNur
x+biB+v/s4XzzbnFtNDwVqAvVmigLnMQ5kSaZXTLUO2DHeCPCZlkxmHAa6R9
Yw3ax+4Mn6Mf7siEoyEjxSaBSTw36F3MLIY7KUByV5rRXTuYwvfB8X8k0t3m
rufvYX5tLOnIm1aH2MCTOTQyEjmlEM/7H4tfrydlOS3iMestQFFZaJx25TGv
r62BdzUhRqhJl+mM81/42GzvJSgSnDFRM1qxl/k7Akup7LPhKemWrsyre8nX
SFoBK9gAYSTncT7S8/z9FHjgvQbou/2bAcylNo21WyfP4E8Dbch644Ye51vP
K7D7alrSAgROC9rJjw6ZnRFC0+95Qt8wemAHfvXXVzlVCbW4h2QOSHr0gnFi
RolCwD+ZGAPOQGohJq2DhLzDC1UNVcjM89TnPU0Whrg2N8mNCLzAx7sqKqwK
7n0WlDkppQSY0MbgWSTVpAuo8HO/wI5Nj08++3e2+e4akj/AwHy3L2x8emb/
Tp1zWPGQFg3T3IxFFEb3e8C64PCAWIQhqDJEOV2nq64KtyXIdDnNfKKeyWq4
6uOQlNtc/eFJXhUmcMLi485xwrGsNrczfBhiBNyx6lAhXvCWDMdZzC3+r2RI
ic2Nnwo89SGuCdQ5DeHkjJemhEXDK7ycCa4Cu7ckUHcRBJHtZrLbYwi5K0xM
a1+F89kloMWBwAQo0p+n4dbt17q9K/sQaUhT5ds46Ro3SlIUHwR+zFGnK7PK
p547Xf+ZNXHQlbVZF0AYQULe66+Kv7/jPssL0jxNvgexu9eC6q2/a/1eJ7f+
ue+LQMMn5v70ZpA55BM0MwilcFetmHma3G1UitFKSSCvuwgGq+8O9eVaPsKd
+7ihX/g4YNogwg48lFCjRWosTLK8B/F0lrhl6T+aQtPatT8LBgqVSbnSkw0a
7HCwCdsbl3xfdz2f2Am+F1wdLyQqoW9D9O3otkKq4B2H7JbhDndeOfQQfZhe
MV/3eicT1sRgYXyYJKszubft/u1mA6C0pjvch59esT4ITpE07wI1Ty6F46kN
IQjNDp1tzCgDY7UP0PtlQ7K1ZTPA3WCQNurbH2/PCFb6Pui9U3xRRt7lwLto
zm93r+H5j2CDHsCJOOEIBVdVVNJXz42ocdhpu3/nH8s9gdlDeGLCCR1LQx/I
2lXA5Drk39Mv29uK8WK1Ip3yL3dlQWiN+5wToOwmSLm12WrjuappwRJihV64
HM2uS6jfGI88NRwajko1rGnwLvGtFcZ/mkX24NvjzGjteqW0h1U5aaRD1xhA
TbM43Sw3NikcL4ExDbSGsL0pe1DL+hqeNA7Vj2JvYnl7bqXHT2aGe2OjYVai
ZEAHe/KMCQoVgxkXviS1OPVjxp4mP/07diQZf8zBc3Rcx1i5Bgk8xdHKVS34
yvdPelMLlp/RPkVVMI3OaVzaFNEbWtG2KjG5E+je6ybntobOjgAaoMDY/ne5
sBNnieuLzOgWoGVlpKC4QakjfMOEVDnEVpALijh9ssP6/GdYRTsFnrvZUg2F
0PYBkSovw4PBt8opnp+tN76nuvs7GnxO17tvhmU9iEO4sl8ojqszS8WbPJX2
bhTsjEFqaX+kE5LIJCEnbGC4lRQmCApPVFVsaSpOO2JYbcSLWSDaqIioT2P+
YoW1IBPtu6Qkn2nX8g/cpEP4tiE7j/JGNi7zUyuuSHSr8fEjvvfRkNW6Rum9
BwxR4ltpaRCu5ziMVinWJxlY8UWghxnWUr0DkyPodCxKHC5TevaE5lZUDOqR
4P2GbkH/PU0wACI9kd1HsBRVPT/Z5NXvcdgM/qGtDR4JfnO+5UUi2q1crLWB
bQwtOPYGun6693+EvKZ215Wd9QKGBCwugCqzoXVNGqKE8M8UDgg20e+naS38
bI30+rIp7QbJHa0IPRlZWa+59+OwcDB+heA2fvMJNrjy/xn+VHMqucWLi0P/
fWoT+vgVgn1wpBwiRGvfOm/TmTTD3wVQBiADmzY7wy6HS3PX203Qp08amW4z
ASOF/Dw36CipIgPgJa8G99+LSHYjtm5wXQdiyYCgOWyKT6ucRqXxGz6iLv5f
OFK7d2tsDk+VQqbWeHGmX/pb9zlzhx+MaNgUzlu4lr26r59UWmNwrxbUg8ti
6QroHNXK7QhkhrxfW2ma50TgJ1Q//aMYGZ3PZ5rR8ZDmqomMxXC/HhVr7VqP
elU7IuEh9UqpqJWrwIZzHvngSM9uu5WasVSN23HA3IwvtgkEf524BkPPXOyV
RgaID4paojUg4ZwhAsxM5uoGPC0Ns/0XmOZSOFb8ZQthRL0nJU7153FedsnH
2pI0/EDiP1NccHvXngmhO7yPa+cLJguX3Lk+g3MYt8UEsy0JWUeJIKPjgYTZ
/ShseDFcE/wlGuacjuvsUDMFzEal3TOHsr81Qs3799hFuytMDsEN3QrwQ6tU
KxiMrR/YHIR8P9mXrlnnxJnNjPE66dEaXjJQ7de+Vyzm/h0tmYluSb+B44oS
9apv6lALEZJA2EERtQ9On5mzus1gjoFTudt0DAAWEoggvuVhKCFqtxCqi4ae
FuUQEke5YP9R+rEwKZTmtjsoMbEGt4Ix96BCvpgiQ3CXOaLKwNIxVVI685MQ
cUTctp0DnQ4IRxzM6M/gCYq4rzAjhyoY2IzzkW65HOlw5pItAzFO7k0lUigG
TlZuuSdVwISOIsygHZHs06LsJIQwajE1UDE1MCn2mTwk29CU2o8X2Na9K3Ha
X8CgWyKQHDc13cCEW55kuQ7w8ve6FWHiOxCekOtUd18Gl3Yr2fOIe71Rs2h7
ILbeqY374cYi/zG+OmmAo8tnKwtGiVcpFxGVpo234ANJJvhNp77g0mbOHS8I
jVmJelh64yI6Tzzm72h3mHJvcotQLAMAP3C3JHg1iTnmUeChJWQneNrBfF1s
wzsi62guq+eMAaa5SRmJaBLMMA7yLH6mLgXohFl+AmOKy9eCo3wkopFXBX6W
r+k0Of7/R4J2aoNr4jG01QDIP1/PSUT6QN6OoVKJR8tBW7GYn2wd7cFduP/Z
JCp3xTy6LwoJn/Z7MwINCLaZohRm1inB8B7GayOEPHSn2yhGGf8SqQNCPq73
y9IDdb5hU7FocuSSg96ty8/2RZ4Tt5+WVKt0XAy8eEVi85CGj7UBFlL1w/ZA
+qutwtRzvi6zVfZ0fBy9kwKmG47yUXu/Vwf7A5QUvsMvWm6p5J8cDDmpn43T
WL9t/8y+C4oaoBeSWQqiXmKILO7ZWDEr+3lo/la6wTRb1nS0XotBmbrQCl5X
/4msA91Vg7hrDJHKICo8BqKU7iZpMUbXAzvntCf0QaXpZVESMstomAHgR/jG
FPw6kGAxASxyI/FFfug6y6lMYqHkr1EYgxnhgd7SWOPP2Luqjo8IYLIaLQRE
s2KbfvE9l/bWIYtysl998VSF6B0VI5HE5EWWB2mVzFT2iYQnsVn0bV62f7aI
5U65Mf/66GBRUzbswNAkuO7isv0EqyLCBu8Bu7G+FwlelDy4gjBhuzgEskIY
Nv+bFslcSNadpG+BjdyJWeVl9BqsUDmQaDHe3G7rx32N4rTOLH/uy9Z6Di4l
xUDKlBtgP5jdXilaVP9SjImHdzhxHD5Ayc8EscDrDjmVZziYizodPgSDe2iI
500i8GSwqxOKFodfcnrBXV7syHYr2P/KBEszvCAEp4Ykf59cTjkTjh/Mkgar
6L9Jl0HOIqT+/lSqAHWJxHKLHoIAC1GbK0ovELm6L9aZV12Y/nrwFUmCPISL
spMF7dbwcaOXxlkvfa0vVaOpC0zyzUVKZ0ot1wx3DP+KnuNtAXDGiqtZCT60
0OdcdqBLx5IfT7tTfhQlYN7P/qz+a3gRjwj17h5SxlaagrTwhcgl0hdAAyAj
+lLRl535JXKvv9Q6saYZsUWBTwr6RzBfQg3btQ+nLo/B59RHEfkKHOeH6OmH
3kVLlsUrI6HhzZB63RNGzlbmZZdeIeBZTQQHypTf5qqeeVJrVrdPNb6V+M+E
4zUJUULwJf4+wwIGceuMg399QGdeQCVNhrBWpWIzQVHUsLJQAfri5dG+F72k
iJ3LulBuSAFyWNfNHKRCM3Wp0VfiSGTrp5pw7nRe/pSEq0QuMmSJxEY3O4tx
5SrBsNT58Fc0WaD4dW2jofjIaCnyCEN44/J/qu3g9tBZhi1TTvVcyt/mGts4
4Ku1KNpYbFSQi5Bst2F7CBgE5rgclBfCdKgFyfAfWPfPjd9WfxHGgVMo1ZVM
o6ULUTdKdKQtCCdT4GANlMpdg0PjUbO+a4VMR17QAMEmP3eO0NhmEDy3zSCo
7kqbS3ZohxLXvA8aF6TTCKnjMTEKRRviwhrHQh2W6Y/AqvPKvRdXfdap3YHA
NAYQfSejLJiyyLEQeKu3iUxL/EyKybpt1Q5i4GH/eNxeDxTdvYUdwKUW4EbR
2P+qPBK3i7C8dWZ7jfeAPfCPgx93HDSnyvooOH2k4zV+h60lf6540IfNgDKW
YVFk5iKCoclQeGgEKqYfrGLxwFcATed6iEs77lbj/c86FG7L/cgLUjG7g61H
9qywml2DTf1wXgXdrxBKOAXX37IzQalnjujB/QUIYGVhgKCZtDPRGg+EMG5R
3FB7dTOjGg2EPz3LfP+vjcfQzfpi+cKndUCpMDkZP6CIMcw1W5FV9CcdOX8h
9QJY7k3BKmepLXHyH8rMDS4Kd3hUDZfnu0BiZoFV0yltgkFLMkEqaoYPAJPI
J4DBT6iAf0lnaZ05btIhH96z6dfVXCH707dthDi7Hk1wHSS3JoF5tDJ3VKm2
8KgGrspd9z378iLLQ09+3XIegAwJugPTKQMgfpEqMIqtA+YDjNyvzB9KFvNO
C+GmlVZzL2gv8r1BHp63Ey8uQTajsyoMWmXYEEh0Vut958qRSklvbp5lh/P6
mOPDD7vuAuYOGoMaw48AP4UWN7NUvcOBiNnNdRWSyyf0XQaiaeaEdQjvZjRH
Qb82rp3IdeayjuOZ+nkVz+k8A3TJJhJEkiTNIO3sO3eHkve5ev40rd3j//Ub
rto2iFJYulHqr8pc3Zos0ca3S+DOcC3akINhPScizqksqHyG7/PJmr6xPO+r
9IzEaTQF25hTAINcmZuyY9VBmUKUilILEt55DESOYuYL4YUP0lbs1A44yZv5
0kwMRFwEM25WBGRStbLBb9ngufB/RLHhdXnnXxx45p4GPu0TD7hNTIRTt7n7
llZOd3RTdaayghbCyoXuohI9bg/tp2LwfMouitxI3fg2/SFSc8tkDv0uJcIR
WHbruLeoy8+ukWbOXplL/ZASRbpf1ANjFRQtdfzAXgEg72Uo/nsAUYQpBmuv
sZnwaOOI5bvt+0mMxrwhgtX9gQJ6lyfGYU7ql3XdnPaQiPrnxCYlK/sff/lP
10FbOMpAFNTCo7wRa/KYnJf+rIgGEFI+R98HeJ/xMUJikIKCgeD+k92jhSRU
XnfpZyPzsZI4lt4CSDBG8eTmZyWxS+RA5OtfF6vv7OMRbT9fLSPz8sdLdZUd
384vmxfujpkPEAxtRmAQN/WxAgpgKrBKVe74qo3wwvp8+yyOtvoPYcM85YWt
5xA20Yq+dzJBE6Fk8gKGbX28nBLwpMaaw7J9lEHYX86SqPpo8q/6mi1X33qe
kK8meKw8JDlVgkLUaITOeSbcHo7lAaP9MGYcxRBbl40S0OmYX+T4UuE2xOma
9uVfTc5d1uTbsG4gflluNLQyeSWELVjypBK98/Yqvh0EHVwWcEbLOy/ZUZ9A
kSiZjCN4FBkkhcrDLCsGdqzQBL6KVhUob8DBqHXEYplrhH7+Sy8JjvNKuvO8
zBxgqKStzQFX7Prwk7Xxa1nAiiBnQ73rkdxQgkw4dgClN649+PHVyC5+yLe/
sEBE1WqUUkDOICBJoSnNR+3sKKSXdpSN69F8uTK4LdslNcqSiuCYWZluiX+3
a/MNGZuqiQ172SvNV+dqVBVvtC1mMVRl1FfhKiGknk+T1/WqkFbGrBbHCnAO
0WT5VFlETrhMvXgnevMlqi4BcMslZTkOimx1snKuUqv2MppD4Bzy5y4V2eTG
32CstU3rLe9Xly9oV4kspPVuDBj1VK8VOAk6wcPc3odPxzybHEWNnrlpaeQ1
gU0ZvTs3vjqEkT/CmOeRd2sYJKGt2SfyQmry9Ys8bY8YIxUAiGzBrzvyZX9J
ynCa+qU9aE3HuvX6VNjq/m313Hk8rUwFiSEw3zM5A9RvGgbyZUFURe2I6GVo
amxb1BYlmphEcHV6JmwnEpNAQrYg/izIx9+IGV2aDkMBZmcfmnVDQJTtHFio
ZLaFJl0AjN9YpDvjP3WVQZnwxhgl0I0M3BVmaRMpIKVux/4pM6HD538p3ATg
q/4+h0XnCAGA2SLUzg4+uVe63SOpBBXbOo3+NBzlyAyu7oRvyzd5rZ8qWaZV
qgiQYa43hX0Vzb8+f50Z2rCmW6x1LR+dge6ExvIiHivJFKWamUAlIgJHMmda
4n83zvccTNB1sA1+5zd5kLtX1eyQsWgOrvohKeAzVjS7uxADG2ST+tlejrXK
lTxe2bgiwXTPJbg2fo8CpFP1kAnt7kcB5Nz5XF/85tL5P2qOBzHYwceEm9mu
y7u2LkpYrPidvrFZIqmj6zeA2ZFKULkqiFfyhjOLB38gG8AREl1oElyBiQjS
aWMJD+Mb5ysdNAbBK0UnH/n1IqmEWXlI6W/n4YEH71uzAhdB+wEBXxdxJr1o
i3qnIwmr4PtkC/HXbrNdIWwKYHIdvt7Lp6FkbxIG8H9ot4EoDHHdzAzy3CVY
kxItJJZrFXxCdPKlQDBNkn037w3X9Qlj921Lyq+qYwF6W2Irb869i0vfyUZ5
Kpkb2QNeQTP6mPydO+raHbWmZ8FlcZcpV5/SKS+XQ1zg8Z5f5jVLcqHGf0Ut
isfbla2tYTXos6I11vGMqGdwN1pRnA9m6GLeWFBX0c4xv0QvltyEqaaBtzJu
GycZH6fXMCFOn/YBM7mw9eJ7KI1OltZjW+jxNATmgNmPCpXldYsM8eNfsQjL
vUrUa8+HogJhuYj0jSAUVZ23xioA2/J3fHKdmhdrpIhFnyVxTHRxFlp9iRla
ipqRM//dIDKjQ+WJis5lCRvrceEpsqq4uJVvrtYLdZUsccu5Uctzy1XuEgES
UUZMTdai/QtG1709ZoQTs6I30Etms9pdO1XsrxJW2EZ3aSn1BUlQcm00smOv
B1eGfNQ9Ny6BKBq8d+C4bb5XP0lQOP7EgsLW8FqyfXgneA3ehOHMtJwWNFZ3
ZuTn5q4WDAuGeU4Y8dmWeGhRXj60aR0gTI81su7MZRjq8cImimSEJ3y+cLYm
9ierp/moKl1Rg4nb+92RTvrpA83KphRjMdJMUzLcbnEy0Z2TxbVRTZv4EjYw
YNJ/B3Nerud62h3BCAhIm6tcMcCQUJA94SrZ+Jgd/2PsF5bBIR8aWBO3i5T7
jH1sbp4KuJMwdv+dkQ0KRCXJME16LhP7EKDEG+hOjKiMJf+FiaGjH5fZ0xTi
SO8dbLoOn9VXxFNVeiQCHDgZXzfi2FHpvBYazCwkcGB1FTiTkn6s0zbTLBP2
qmqbPE1KkKON8VM9PZPNKbhBwybyN9ntHACIo5PTRWOWtp7TDlt/z4OCvpdg
o4iWXINGHYvGiyIUS0uijjt2QpHaSoCLZ8mi2/p2isdRKUVIFUR2znfvk7ud
9kZadAIZr4h65m0pU1JoAKNfLvfZKUoGDLstGu90N6bbbxj00chHsRNPQybD
8ljbp3Y/fkkFteD+xNTOkEk6HGIZPq1mpaOL3pm2vZY2i574RBESuAjOicAt
XC9yk1v/8AhuF9zogON+TpRMrokWFrFUQ/yS1jlcg22OJhDokXqZE6/2kuyP
xVgu3F7LMlntVFvkCNy1CRBJFC65WTuario0nvto3ZaJ9J8U6p7xJGltMMsx
7aVRjFcogzCvErLjpevNTP1ihwnbw3FYi7yF7DxjiIIOor/MH8SF6ntaELwh
JZKvyHI4rxAE9yr81QAkH3tXfYJjGWUD0i/8vxs5nPix85LqfbdwxF5w0NsT
oZ5Mf9WkzhheIEH321llKp0MHVrtkmjKgF+OUhLG5D/QZ6eIgTkoaQTjx1bJ
f2ZjdxWa7w40TgeCZ0z9IVvLpeXn/j8TE9tCHhL6vFZjD9gaIXth4PCerL7M
7iVHcSjzpnRYyOSuIhiPuWM7d+mUVet/o/X78oi/D8IXkL0/5Gadq8KNWx/n
MNpnOk4W7NZ4iObKDYtiD9VgNb3+o+jLjbfbUuLLC9Yy2sC/XAO1a/v1ZqmA
eSjIzvt2sku/rmBW6ulvYBhb396IJAmr+Ga1SiwT2kDm4NmjWDEwDZ0ALhw3
ac03S33u9iKxyxchFzSZivWRfH+LtZg1LCg75EdFQIHIzJ0kSYNG9twWW18w
UQwzEZ5IlKV+B6+07yI2fYJrgJXI3ocwSDMEDTv7dYkbH2dUWtt2yD5a8OAx
tzu//lxLS7Tbf17DeEtTPkR6H94Lg/iqeVBi3S3evEaFUZYz61FS51BICMjw
9YoXFC6aFToLoK12Oyq8KNU7lGz8aqTYlFqCJIWEU2Px2liES6xAWYFpVX2w
t7qbkcjfP7KNBMMabika7Y/VMmAL5HNX3VbcLJFhkhUl6Zt9IijdRjXHoWpT
pLfKljaUPAnxzdVIL6KwdlPjmbV05V555mAXmbVfDUb6Cg14oLs2yjFdh0sx
YYqjsBavq1IlfzrRzSf2bFWNA3cdyJ5BMCC3ZDZHNdzGIP03clEnr8qYz2rc
qdu8VMaiudb8PDTtS9MFvgU12WxyHXSdh3CXC/MZKzotW8mx5KrSPdUqLXjF
EhFGIkJqypsC80NADp2v6W0/EEESKCPRxTLmStKZCrfNizZ1+LEtpNq4jqoc
+mPz0d9U7YEZbwpxIfHsT0MTL93ktawcqRkA0qqDxFekJp6neNVw6p8zpjR/
b+DKxDrmr7/gh2LK630kgqzCkeLQ9GoTZAk2OaOhXt06wFsO6KfB9n8klFni
Mib2cfsNca5q5dDHR9A8xwMieTQxIAaDO6mIvzCaXSO7NZ3N98qF5RFDHr9u
YSMnVkDMZq/TupcQzUg6LOYl5D5lla7n45jqf/Hpc4f3y3+w5TA3vU6kBD6j
wxb0cVRjua/1dNl+NTAgfgrgJbLToPyb2nS19atatc90Kl9RGQLC9s0fwelq
HMiVRurTFE2THObeOacYpAjQrQiXxDRnc6C0co94SS5HRUekKsEBHuJrl05E
Ewc0OJXcoMFaMN+XRVDkHaSHA8FizDQKUUTbqD9KvHvQwGUR3/JjWRCzFNbL
a1JRu2VOqRhjhY/W9u1V/Y6AYiRBhLDKohIgvEWuv3aTVg/MxYsJLwv+VpuQ
rEQGRg9+kAKL6tVX5Hk34GLmvatECfzB982AIszcfmK01FKEYEHCkxfBtaSV
VQIVLdu4w7OW8TnsjDCIugokRftB1ddJ4VHPtETD7OoJ1XdxY3sZ/ZbKvXhT
48IJEsfiAQsIxb67BQvTS5OlxvKRdiK5RnIdMMa3VnbcRRPvRSv/6XbdW/+Y
zLL9XJiEScy1Bt27+15c6Rn/H75dedwoPW074WGXHj/GDR0mSbKcmyFMk5cW
rTJk61hwpopTAvEiWxLym6L/DMpvwzYEG6oVioELY0OtOZEUZs2VvXU+w5vq
jkyNp9x7bw50Kr9iRX9PWckDw45F8d3QOvxsZ8JuYt8a1ysdw9Dpzq9OeVex
T9DOjKl7UvpEwetVF6fHgkH8JIMnDES+VvJ3DdcSFFtksBY2/VfFissGfijt
UzlUKis1hkbiCgtk0TjCZvnk4YuYSa2X8eEtIbrcltveGHtTQaEFfwg7S7KY
SGjleYQrIA4Ykirm8xVxoT7uu7WF/hNjdTauAOX1gthIpQRSQylKjRXJu93i
KN8I3KK1qQ0Q4469I+6i8Ye6h+tPiHz9xYeVP94O7001Zih9TEE58/sCnjL5
29dSTvj5/Rb9Q4RoJdXKbPcSjfxNqvh/Mx593aMTWDyjFy5cKn9t/gTSg8AG
kQ9ZMu1/dcJB2Xuqaam2sSnJdEB8mGPjJ8H9c2yfKuOk0r2JIGoJdqTddhJv
HeSsIJ0fLc//jhzVuR6gB1gkq6d96jovMfosgGiDsf9vrlF3+Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3HpdA02Ie35ow43/wevt7rJqD0tu9EYlERZjzqrqezvMu36mlWjtkWZqrU33iiUOrsxqVtrz4V4+jOk+MFCFwr9m5fON0Mcs5SYvhDE9RYx4oNA4xT9j2orDlvt6WuFTH2wp2PLuCsaHQUvEh8oxbnvj40vYVQzbcj5IVGWhK82HCsWlYu8LhkKxiZaVaIuvfMVExUoes0gUELVaxb1wuk0RvcZcvFDEu2W8UgYbF6PGUQJ+BcN+J0sQyJIWujv/WL5d30xjIR3ys9T+MjYt+9cZhBds6Kuf46+NAbBiga5zD+iZZq06C2P4wKTUYOZi+6wF4dDGD5/MzuybfyND+3DdfSHIZ/hGSvFrpN9oWCqCbFGd4K3P9S+8oKWUS9bKWyPHIgIrxZ4gRjK0AQ1qCdowd+kLWhAzY9VAcOqnRk18sW7dDNwAe6Xr23AIRQ3vSdLGY5fbsJ9dOWzHEJDC+kCDhje5t0Dnli3BDDMuyydhX6b0iHxKx3mc4U1PdGj6lrt27RSCpyitMMLCQ3LaNQdJzxtIByv8wcHt/QDRfbDTwb4vujPNLwMqMyPjH4yocObDt/LI9OeJ+LAQo7baDplLRL7nEZs1Jy3DaN657tQlGScBCIFXH2GsHWqhxJYxxvVyTQB5uCjoTbvlqPxMuZu8WSzGvyGO1td0lSnOeLt8aAT6mRWMcb5T/LmkvbnytI2xCrQIMX2QbJ7FSw0U1LkTCT1fOSpYRzjiU8/+1XHw/l1C7feMxJGN6DXEN5H582tSjeEnJe4jiEFY+g3y3m7"
`endif