//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GXLrM5tj3WPVJM9GVLSALX+cU/TWiXFJiwz60rK4b6qAoiT8CC/Dbiw1E9uJ
OqFQ0v0pMPxQ5TGY3xtyZa0x9nIUKCC7qEZYzDXY8zth7r1b80Prv2p03u8v
3dXqH63q+wC4cfdE7ISKPdBmJujdrnnjct1IXyimnKWBEYVaP4dt4wN733Y0
e1F3//8FRj9jy8q8fd45DvaRwt+KdRv2FGbxZyQf++gYRzUhGI9thv+92Uwt
62HavwwuQgc/jABFg4lsXk86Hw0Z+guE3NM8nczc3KACbH9F3Lp+JlaV34DP
d5W8WsKcR6GTATgMBpec6TUMtR1LF2jz3eL1kIUPMQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KVeYsbg4Ludl5GqD5O/y8yp/ixiKpj+GaskWOwTYKiuwGSmlEzBwbJfhsIuQ
tS2N6/khZsKL7N7h2AvLvRVB347psjIskaufiXWBFxlG0KQM7KEy5NGv3Yrw
TwgBpL4JnGsbGHI6IE1Vf3C54XQwOU2rDoQJtURTzIz8KhT6//32Oc9d14q9
tdNsuEGroqgD5NpA57rpjx/WeREeFr4Nd5nr8dlSoUJrm7OfaiaNuuXyj6VZ
1eCOzv+LMFPllCwm5nOTbe/8F5HC7cgrJbcFa6+hhan7MehZFMtwA6pGwuXI
GXJgkQmZpE+mH8I3jRqHzw/rtezCYUY2ukbiWcX3DQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JOvyw1aca9GL7/9zFXflGGXZlOEfC9foPzkv/SNZtvSJ5AKXxHzrUc5gF23G
3Q7xK8MrgxhtE3ms6tnjkTgDrO7cEQqeE9MZssH3XFTQ/qpI1+IP2vFSTc1B
Ok1yVpWwXLNQs5dIrZ/7jIMiN/KFMQlHvDabSaDP4sgnubrmBBGAsecYC+JQ
LsES5vguKCsX/aUz/98EZ8pAyuqEtAmEAuHwLvMDTdunUOqrDDeD97DEmSFF
bl2nDWVKaLgPjwsaRmFP8Lv5x6UUymHbVoiHxYW7M6/2LBvqzUUpqoR0jtTC
Mo92dLw4askKuYz06V3qlM4OyEb0QtJHTUulSOIsaA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BOBPXP9tKTpeQ15qRDQOBdmQANtHRxQ7BN0Ds1Gh4JI6yLPwwSuGHNCkSL8D
VzKC1bVUrKVaOEP83Zf9JipoPGhmKN1df4BHowueACmToExD5n/+ZoSXEK5F
BnT8AFCLlBP6/MHVllhqplTzWhdbdGamVD4T7wpgoXF5QJpUZOs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XQxXlok78Hdgozj+BNTS3PZd3PA7g4mbiC3pXs8E2kTiorFDBks2Has1hghC
ri+MV3gxzphMgp/dHPzCh6b1x8wZ5KX5cxVK7GjVAfespO0hxfaOCCHIa4Ja
X5l5LCUUk/iMJIts+HMFiFZ4ulY4U/L2qCPVuUGUjpnLc/8N9beqU5w8w2rD
C/EBuNarabPNFlI8fJMz8ANYWM2vT6kv4F9tDx1RsZM69Vg7GWUo4C1Ss2uP
udFojtW6ZQQBH/By8paum+sU8cJ3ZX2ykLbCAGlmmmgnI71iwaVtsVjS4vDg
7hhtY+v4r+VCGITaxmBc5a/1DkGCExRvbM6dyrItgkzvVHUY7RZNKBSbU0ZG
9u+cHBt8aDKaGTk5bPlQbqMtb0PO95qteyuKV/n8HWbQeWTIa1uhFFD8/law
0aWH60t1fGdJDv/zs+A5hecvhpAZFIlzHHO56HViBcO2ZLeieS30NTg5aF+t
gji9T5/cRoFRkjPAEZ7eUkFvoQwaEQAs


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VDMMyIAScMv9lQzsf+pthjwoElbvqeLKqurBzsruhvlmgRlfwyUk7HIs+AiT
Vp32rIC9C5NmETFtSf1m7hbdVnOfH2nbG2TL66zm/lAeRDQC2YP8xjuUv+9t
SjV3rDm8z6ro7WUSRH2AY784w1R71ZyOg5s0R300iojknP0XBu8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XJhZsGqH6d+bNGZUUwiT3+I6+C+l9QCaClJuJjTWekYkR3LBu/HUk8Au3qxI
sMSfDcLACZo08k9eU5rfZRvzqudKBGyJeHgHElDktHcZHcuNtuUzzfVLyuF4
NsWkv0xWawCvzQwGmnw5O4cvyByQyQnPSHXcsXl/D6b6zA53KqM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2976)
`pragma protect data_block
nFFlOQSKo3rHcitzO4AjuDHxeFMH08SIP6l4E+uglEtwotMy7PvIAcuQsfNX
TMyPn+rOJeisaduQk5BFDfSihQ3aDlW62Y0J+iQqzkmvWlhqnYThBDdwnWsi
6KYgWqlGEXZDS4t+His3MryAHoKQKDbWBML3c/vnUC/cIVhKITj32ugwDGwx
yxkSF2h2Vlp1A1IhOSyANJLB8t5FgHuXkNJxN/NitI95Wq0xfBbXMQZp8TT6
+UQGXJITtX3ztKQL3rIk0MdlTBWRTx9gakdXSGOkYSvjxuzpTGNIzrRg9nSH
ungAML6KZb8p0UN8i9xWRf13XOTO5bEOLG7uQmI53rweK/aw48iZg3SuzZ0q
9wj0GvmyOXWUSZTzuEGfn/z2W2lBjXXPGQf0lFyjlwGEN1nnZ+VHVWSZo5qq
EdRBB39SgHgHI5ZwLoowVzxec+OWLMooMvxJ5wVsKbHhChOAju1B6EAMgfar
57ZUBC+1si6U0G2RTbWEh5QJvlS75G6WC95aM5WH0Kc41zdXu9mFc9uQIPxi
FmugHD836MKd5IXfT9lB//KAqPOMy0xzmvpbcSvmMLVUDTPpGRK2N9vXsit2
jSHZm21bux26ez4ZS3Nt/S/t2RrRv9JO/m2npuKuqutgUnUAMvpJTTQTGWqJ
ZSd7CKyBW4tsNHu4ErQD0jTSmYCNPQhgDm5C3o4sFT4Eg3oVcbGJxCV4Hj51
pTOU/jR20C29c/FD4z0+ohJMln/Qen5xlQvNuSOJLZLwk9fBiPchZOWY7pZ0
n92+z5wUPVXZMXUx0EJWTdGXnO+VL/oZ/12WdcDtnqbfIUUOCgcGNObKvkOm
SC3GLnt3kvDyLfzETl0JKambrbQlwhPNnMzaiV5Vl7DWTJ8m6II3OBcyDc+n
uEgJdZ4RAbeQPVJcO0tI1Jto8XwaNzzzYGCXGRdXrMBE7RPVfAhz/ngHvMNO
IEdtNneqGcvOFNuC+ocMGs1OJQJWTmg7s/hoNrFL0kWu+lfBXET3PJVs9Buz
BIqeLHNt8jBFGoT/z8rG/UwZDttXfo+dkLbFTCpSsrgWrheAzkEHIt0FvWH3
mPSDwqDkpw9DvacojFIOhsfXvXYM7RuVcA5NVLaIcrvWfoKo1kuFZUriVCGL
4AXYH27J1QIVBMdjC9Afc+RKHCUdewqPFGwHVJBfec7uigxz0LMOq7fBiNzq
KjrqNSyn4+bCfP5EDbkrFLu6rdh5nNtcEIYirCTtGm15kIa1KnDwPcs1V4l2
5UOnKSmNmifPkuFWAU8DYgu/YllFkl9OvYrzeXCjFylh6dnfS2GMcrm89fNQ
AYjvusrGh+e/QRyzHNDugrEoI/wo9bnYfIVYXiUlHaY9XdLqa+JUy1zHxYi3
uWeYpZGp9Yj4G3noXzy74wNj6tYZZXnaAnKGOqYaLctTGhG3K1PV7L9YwHM0
3GpXP6t2izhBJxzZtyRU7dEsbchbhSbPgM3kmoa3ZHHqpKwlAsk7bgsGWVEX
udBcKDrs5g4g0gosGfbYIBNUCoQoRl3L2WMsNvBeOJLDYGbTZ7ErnoCXs1w4
g7JJwenhcrIj1WAuiNXv1DMYSP32x73do8iF3rjE9QpKWgv3oJlkwQIHw2wo
XC+BG1OmMB25tSxIlUESV/7qmH4sPFbX+F29euGppjfVkCK5oLVQgKINscue
zIp1xjiQcLVdVZ5nCVLNiHDViSHlYwqZBQ17tECyhWxgLA2qzRsrkMv8MO1w
WYZcnJEKJy6zcEbgPYDHXFqQC5TSHNOWIKuaR6I25ybN2zgJKrw2K7yzbEgr
mv78QBRYngYmpgdcwu2ncrQ0K/76PAbeGVZ9QHFrKl+tTdEN0/y2tsUQWrG3
1QfOtsZZUi8W9vI98ZDh/4hksJA0dWzBuIQU/UdYVV0Wd79YEntdyOFnFWJH
jd6RB5elwyq/w5lLtWxZOjHiKgAlDJhpamdT9BojyP8x0eTJWHkdZVEVwJup
eBjPs0gpGJb4G2UkSfnwr/LAO2RXpFOaL8frH7L+fcXxBn5umtih4msgZ5xm
y/NAMEesr92Y6rw/dALCqKkirJaE2I4yWuZ0Ata5LmixAAC/QN8vcijBHcnF
Y1l/CBOuUNSluSnK9tueccCjE31YhDwv1hTiWS1Hl/z0d5l1r/qxwVurgAeQ
FKlsb4hSemTtajqlg0SnTrkBd7smWDckwxKQRerK5Wfa86IDI3P1tyY14Lwr
vMVmaZDiMmIAObN7KUG7bq45jM2k3PQdx98tf7X6uEBu7vrX3beBRiSW1oyB
q0pV98AqwyzTW5VoCUk6YvE7DX9ciR6O+5FuBJAiEVsL7HcsNUCg8l9LSKXu
qCfkIniAJ4Ud0eOCfTerFDJcxOP3JRH3WrEvmSbBP0yVo3KRcKPb+QoSCLUT
zcWichBDzDwWQAL26FMW5mVQn9afWL2PYQ1YD6PItr3N1xg5lcXClj+x6A5Q
Mgz8FGdUA7pglbxtStnww3s5HwjknCPhLfjNIfpanEchpD+pjVndcxNW8qTZ
rrIdYh4iQU5sP6IDRtEX8B8qpigucgUwR8QiqK82czVVM6nH3T9bZjDRicBb
Fx1A5ONezfGbAuXaIf5BrQ+haqbLM1+4/9a/DTjf8sn4UuD4x48h1aWhvzDk
rLnInIgt4FXwFXsLC+jOj55vmKpNehauHz8rOue4TepSOLpBrYxyw1ZqQjaa
5qb9RJb7T8dlNohGGQy/WNNZ0WGErAKzxJusTjvZiQkgd681Jm/UNC2aVeB5
CqCb0PvyFryYhnmu6IRiKVF13Kvv4lODzMKupicqCGejKkNY+JJcNmg7DIGM
wVjdAuxLkjN1K1gCwbbYoLSmFrYyAvwZFtyCmYtRL540qzGJcCZ+fR1n2/P1
rZdBztWYGN3JGuG8vBlre+PVXt2RW0QaC+n8M4P0CIwhQIZvJy6pFO/UJvZR
RMavedw4+Rnv9yE/KbDXm3LLTQApl93uPGClnAtfJ1T+O/Ul8H2OC7DvHAnU
lwKUKLSiL4NFvalaxqrNyOy7Af7HfVhN8I7tc0R69Nd8ZyVOOEaFzGLrGBnW
FNl+K0pLgwybcsq6GBw6oDnrCCbOW7FDqDCtrRCVURj8rDOeK17VZvYgxgRN
KLvW5u3dfnPFEYnD+TZmwVdxgjHSStZVt98TatpDA5VsLtSc7XM91I9+nMxf
PH7wEGWzuTWi7eg+UdEAi5VGLWZU+1ssDl1kXw6TwKXECrUvO1AIcbChM+xF
v4f20siebL6yYnk26mKNTtC6HHvVovB9pvXLA8orhyYc2yzQ8SQyWl3oD+gr
MwxS+IM0AHLfyd0WxdQSC7zvsBzpEFa1kSIbDjiRXChOkVMDxrm+WFjbHij1
3dt1FgBCcx9YqbV2klrd+62nuzx5bb2QPPvAt6nWa3I+xCTlv+0M+KRWWUxQ
Q271D8FXWllm/uAO9URJzzxJSen6tx+WGf8Xh7+bAIHYvHdgR/JHz5UbEFja
VG150AOXnTUAVevZqH1+4lPWiKMbJBbUHaNbA0oXEyRC/C2byPgo8zVeKurc
lxrMxIBENJOVCxrumg/y5uNfB+2nAkIrzezcwb7cuApquKsnqbyhhfSK4BnG
M9XXTUzrXvkaXwIiY2C7ahRk97mu+vp08YaEQYZ5IHLHrmobsoZSz5YXXkuH
gbQqi4jDwl5vM7qQVwC0I8ZuA4BYP6NOQBTtLpX97wzzNFUG0UYp6EHfAPf9
xjQX8jS/+IeKTvX7aSSXlafk/puY0SI6v2XHnacyhShChxcZfyNKQNjsaFDX
UgqFzNq9a104oqZQZg7t0ohM8120sSbzPqrtiYoJvuXeJKaKnd87UNLnA2Ed
k7hw9JoHILGH521F9ox/7v2h8ytUP/rG1FMACM+mFhFn9n93iMrNGaPx6MkP
kkOxaWLof86cPfXiT3uSqBRd7ceGP57j8377TKxzWt3agVbA2Jybg3LpCcKB
SSukhN2X

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG1xACKK+OH9lXFdb6R9dYWuwD19m1jsisZP/Y9qB0XYJEq9WzwKXMVdjg/QCAWOhS8ahQequU51mJ4Cmjj/1ssJQJut9IRs6BeLKHiSB5bbGJJI1lGQVq0VPxDAJwPexDdh/S9b9OmEHvhFOtnvSkTipl4d2HP/PGv13OQtkbJ1f5ys7wgS0rAFqWZ864oINkra1OibOve653BxLikfozhoAjhU+Woop76mM36aEfBS8q36lsfiC3ArtWe5m3CCe3bBp+dcMlGWZdP5uFrCd/KfWANedZ9vuyYt9+w7PVj9iBPLhG88EL+mzElrJ+vDsWVnozvG56dmt7/phsZYY+PZO2FEJoaLWkIwhPPABH/wVadMv6DwA10okbfaKq0DosGZhh37qHtKzZvz9NJaQ/SrmuKQVmuQm2G9cekbS+Rjgtd2W5xMWPutj1ru1XqiTbmeVgc1D2mdB5Vx4xTTr4NCHOn0DSIy21jKsxKLYIkHArguu/1ag+dSNGoEbSRnW6wgZ+R34/owSCvc5i3gc9YPjRKUfmQyaYDPiBGue5qfWDT4+lA7aCMSI5caxNOKy4ntbcu4n08HK4CwDNYypy9uodJGYylXoth5adEw9M1q5rTQoo+L2eFRuma7i1qDGE0NEmYa5rKonT65RWcsdmv8fN0LW0UjWSSnd9c2hvUA+8c6QgDHzRA3/KMgCw4vhP3Pnz2Y19WntltPmPO3OrT5Nvb6AmdEM1PEMNYuc5yaDpVdB8rRN4pP3q4qqmzDjfjvzdOjOe/zzMPmnd4LZ0Yu"
`endif