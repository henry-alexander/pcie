// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lLarpL8ArFGv6HYllnXFyWYx0bDJBctTVFWns92rYy6iRfAqn/Lmy0uKpxyc
xBRVNMHKrRXt5QcPn2g7cvGEEj2+BwW3bFNJoWowT/nkppv9uzvFlTRYaynt
HCQEzCjVyGs87GC3igAW7WPbhO4yo4I4dT3Q/uDZc8fnGoS0Z50Sez62CaT3
YmBrxbzB+rREHC8QyLEIqIcnLWYeGYC1gViSOHmRs7AZhsaRYq2igK2SYNAR
uILW3D3gxX+JPfimIqGVi+hGgnpWwyZtu9NWBJYIf0XzMbzzf3DNFAoTHKbj
mg9+LqGYdXeSi69aCPzHu4ZUstxlUgQjxAQLecsYmQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eWZoQNk9s8QD/u4T+UJNNWF267zD5Uri1q6xBCdLXeGwwgiSCIxQCAhWpgtl
W/DF80SJsK30xp6yf1kdpbnzf49AYpHFxJp/LYacax4C5qY+/pABCBjREO1z
/4KBU4kAtAmjmzemqm/mcnVL+sGEbY7fkjZU+qh4FVLl9d8QeK2FcSRbUTGe
wzcWooLurDBp+FBMGDpG5sY96yn4fSa8hPCDgoz0ZjM9RJ3Pqtay5DB9hKU2
jY/TnSEWQm3zlnTQvXbKjf/o0N6kqih/XoX4Dieyy8r2b1BE+pwYcikh2z5n
cxTq77VWs0j/C5TGm/stdYu2qQR7LQM4fO4PF6zA5Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kUxTtlaArMu/7xOgaz3KCw5B0AgGFvuRjQ5CNudX1LxuR33asjNrGrfCy6uJ
OHjg0YkzyB7Zhzj3vOgr651JzvSc/uABWcu4HPZkcAAKeHvdzgOC1oiKAWuY
IkvGXsRbQTlWEQZLA8IvardojzPL9xbQrdnmcp8k86lrK+v3xC65oaec+2FF
dRqOyUUbLSbTA8cnluwJ5hrogxh7TpfylMVXMkmc6bDgQWU6JgwLHmzSEd03
oao6KS/PqYiTWsdiCONjWofCzz2tW5oy+LbIiHEbzjwpcLuFJajGGsj7eA1G
u3FXQi6kdppDx0Tv3gRd2U7ShGfQwNekD2lRPUD/zw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nhL2b7kcP7/OzsAfjYtzW9DsZPVMdtEbe95vzjJepYv1IIC6vV7bJIxkov6I
w89XsnVw1c3UMZhDKsQHZwXVI26dq+GiVgDhH/kCzJMdRXCzPhFsPx/13/jH
Bcpz40Qz4Nl0R8XtYcJ4DV0kz5hFLtBK/VABqJ2K+ha9vdbHOQY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
w3wQ32hWrMf9WH3Xz3UPvdPleiaMhu1AxwRUwbhM3QiiqtjDUTJtRjUCcahe
peVDHDP4fFVuO6iMcal+itcQCGeJR0gMlq7XFi1nY6swyvHnp0Jc0ITE5uDY
VgHvcJjng08fQqY2xkYinvmaDB94WpmsC9xHwbHNikVxuZXfb+aHNlV7GTAA
SUqCDj23YhlA86cobDDVaP4yJAljqouddSwtktn1NXhQ4GJFk/SNHi3KNW0g
mt3DIN+WncolXwEGO+IAfe28OtBpFtFGog99TYsAXFEsyo3mMbRcqmGcYq7u
l8JpyeLblqXkYIVa+vPknUmaPTdcoNf/CVdhPvHw0NtQere0a8jVshTHV6tO
R6ScpMmCyAHu8nsVnwkk//wpVezuZedhj01pE017/SRUkOySYvun61p63t2z
Wqv6r1vhdOmHBSW9thF48N2ud2IKcLRwtOct0c9YmnTUzQLGt0hDP6R53Dt0
/kmd2ZpPBE4q+NO9+ULEjlWrZVlbTLlg


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QoDn+xDHGfDm4kDbIfMMrSHMdAhZPayyiOpUYIQNrghSvj4nvHHIvnbRJQoK
LxrOzQ0GYqVSN6yqicGM+noaq3q0csb/eI7DTdZZfE4pxr81Pu7Gqifaxqt3
byb+7/YMiT1S9sBqbPMX4+CaXzrudyGRT30NxQB4t+JBzG9ZGto=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NK5Qs6A+5pElnfdu9JL9AaK9RBP3upN4bpd7wOM0L9yjgNmZs6eRwQp1Lpah
WN7PRZsbQxMBSN4fwGoAO1vazaZO23VAbS+v4n0gdkDdsXmmtquvDAk2YZOM
MlBsY3lqgBQIth3AxOtVOMUgK334e6TbY8mR7jrNqxTUdUpKIrc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6720)
`pragma protect data_block
dZG52pwBvIStL5yUtB8H3LzXQhIHzLMvctYIJiUZ7qGryhXv1tenmIn3GpKK
0VI4jiAjeP0SgCcJQklu9haNdcN69r4ISfLLC6RZHVLFUG0SGEvt78sYbHu2
eo67VqWqDfPg018pZ37gl34vyDUQLhVL6RtuUub2/9yCn8CgZtxHV93HdLv+
mnFMyLVzFDknYC5GMeB6lznCk2pN0nUVQCico9rTXh7xS3KHkVvpYtJgd7Qg
0WX7rj1tFiiGAzV32goxOMhWpCDMDbPVRjBqO8eoE7QMB0oRhvj+U7VgMwOt
fkkLrRinq89R/1lylMYY1oe1+a/owZ20cSdVE1qGcrX5OMsxXbT3Jla5lhHs
6C1VZM7vO+H743PHrX4bIpEmmKpzFFTWilmO+U3cBZ3ylLKn9IrhhihYpRCv
l6XVDLapc6PV4DEPNZ5T6QrXI/vozIvc/iJa83JibJ3Ouz59IjviXT/QiAdT
ImrtcFoekIcrys4naOLYG0Ua0vLqeKOWw/EoxmsMn77Vxzu8kghOLuD7zLX3
zqmnzu6k5NwOh74RXT1dxumQCRGA/Lu3MaFM47mFdBWUlFDnimtUx3F2JXqq
I/kUTzTdDCgmQ1XzslonwVStml20S1nLlu0k8UyjIA1RKXUtMcCr52JC1k2A
P1d2gtH3ugl7zEaGebI2m4cuzWcB6kLy1BVCF3epZpPT/OMOcmkLf4aHb9qL
W4NX6tU9D8IaOSdU27ciYE0ef30QFgX6Y3XfjO7z45qP3Oxe3Hilie0+fKoj
MCpZtxfJZ2qN/qa0c6d7ZqRPeuNz9M1HxYr9bSRQ3r0GwFtps11fd6d6uUZq
VL7qsIkfwYAIX3AMPRhpwc0C/oXqUXL62jCN466p6ct0VvWpX5sGBTq2QZwn
GSfkbqK0sjoXRI8H7G5kbzEj4KY/O/GkWpvexvs8pry89JsN1j3hPv/CSLbr
oEjHJ26eOj5PnNLsDDvsN3DgWGDOTLvSyhJETUQB7btgUlP/5/5cD5a77PuK
aUkXE3NbkLz9dsLATCXffGpDmiG2qL31DqcrLw8MkimXR1UaniHqHWewObjx
tvM1GUb+fiJ4UY4lx4GWv4+w5gnD7kYkr1y9pTBfiMMQrqAFJ/7osDWmeJhA
MaEdQFLrbEgnQ1pfY3m8NzWfRkb1v+trdTrWsNDVx/ZlFVjcOuydpWRa07KQ
R3FkVnq/+Y5ekSZjcCSdXnfnplnC4+5G9DiL/o1DKQNrH3WezmSEAPQGUe5E
6e8yVU2Nw8aMBrWJ/G8T7uKybKzXszCmK64pB6sJkppU8JreYOa8ONQ3BQNV
ClgC0SVPHxfiNlu/qdtDRFAqwvStOGgb8sX3GcQRz/nZUpfALp02v4iDrgaS
qfzk4b72IujbrlTXv3IfK4O6RMgRyjPaStSpiIuD1MOCWFvrlfpI4u7qJIlE
N4qznMLH0aoBYikdsfGH266AS5jJ0Ap1KxkdlDES7J/ZdsQ8WpPZ7g5iaft3
UZBUghNp7WJUalXw0FTVQAJ8T79ieR376gDT+rK4MYf9sYsmpfw4Fx/ZDi4M
Fn4kgSGVQElFSSkjQVW8ojvMlOoDlBiAIveba1tixf/FjLb+C696vAEuO9HI
tGYk2F6FGDyeDOG03VUsmGNV+H3wnYvAAucYdLIrM8dYTRCfXjqqe8Ouhhkz
Rln0bCJfEALSNR0PFBg5JYR0VHzVNNiGaHPiAscdXRP21uap9qB1XA2DAJru
/3CSDFZas5mswRETNCFEFKvxXrtzkEVVF0GDew5V76iYCT03Ta6xLcrCxa+a
TuUIuHktXyzag9JMPqfbuF/B5QX1tEkfwoBls247vO+YCLaeI+72HMNX/4wH
geBmlWS8yswtG9v1as3AAsNUhb58H2O9pcnPOUGufLQUgSYN6RdQf+fabdNH
uXSTRPa5EADeS2URrjQ6mHIibQFfGie/VojEI/K/PxKuLe4/koV8oDcbM2MM
XWj2BT6gxo00O32orzl6sgT1iF1vNs9B+S7nQ805LJ/HrG5Jbfkvrvc3uLcs
9bocjVIPgyS86orV4RyQFChUSK0vmejicaG9feyZvpfcBvzIA5AfOvaXnhqI
b7YY3V5mnKL8uBsqP63niLCKjPW8Qiw9TgJKZXlqsXIZCPKEdHDrVtZtCgOO
wMFQNpPuMI9jNtX/rObmCNG1qqZIWTvQubMl83TzLXUh/xuWBFNUmEwfbX9W
PyECVIqNx6TnQaEQSTTJQBlFvrYdBytWEWyU/PReJXXNV7SxFYhRLfzTXjb/
0icXlU6kynHeKDgOkgpJsD1QyaIPJPr287pNg52760AeUY6eL4YX8tDleaRv
S0KrmQ+l73m6zUGEa/Qgt9F2M3yBWio61IMTdGIcOBDs1aQTxKjOCvHs3CaS
meOS3NtMmDqw5Cw51l9I0EC3N3/gUpgQcmtvd8SW/0tosbHR0q+zsCdvVy1e
MZdoXZB826VFQhk6kXXlfNqVakmuZWdhKolnTUurhaNFu02TRvycVwL59Y/3
7VhvOHUs9XDR1JL/1daBoyiM00dJxCuPXveKbv0ESIqt8if6DSRMldYYGAr1
FXvO+e1PeGXwxkR6ZztN48BTks44lKPoEoaJy4GfPBM2WkZ/71X0Aik+xXpZ
v4LgXcwnaawEG5RBt94v3hFciOTYBVT0w6fS6tcVbxLFv11IuEyOZtDups0X
6Km1IvDleCgnCnPWgcJHgC+Wk9EtYc4q30ku7Z/sajuRvRpYBwLqA434I1LW
R6B7zEkl12p6EVPWtSycZ05hUOhgeQxjxp3H6mS3YPacTP+vTBaLOS8EfPlX
58M8lXAMxmTXuh8N+zIY5fPFkcv39Rm9F8Nl4/T6jfEZ2XALlc86LViupvuw
0ZQxbbVFx7RweMHGtRNavtO4FUsXu9vSPUzmJ44rkab5JqHzqqlRCB5bfJur
+64qBw148OTG1kdv7ULAS6iukilQb6GcVYr/1BZadrnjxNsEuINkJpQUdgpf
2el38t9pduseixpA4UbWXj66ggcDQLpwwtkLkIUER4AdhGNZoWYfywZaUTy8
biU/sLsyeJ3BbO9G5LKjZ4aupacs8ZApgc0x/cv1TMNFwtaPf+x/eF4rPR30
Ck9BK5Uy2jVl9Izn6ccKxPdcC8SilbbrrupE/GnS6WeugEz8A7l+1FvOQ7V7
ILIWcaJo1yvV/eCL93CInR6uP+lInvLssDw4YPLRvWD7IOBqmsqOmdM1ld78
Dn8frCmax46ZaRP+/r2CVd9ix9FFBgDLFnENbL6ggsEv5Z1EgQx6Tj1kfm54
iJ/hOJ31MyNK7BpPWrKITpg6foXjw8LpEVTpXU84xh+FPwG3PlASegTb/6Ll
a4dlxwU1pZunh4VmrCNlROzSEg/EltERy23o7QAU1PST16iHf5gi6AIS+SJN
NHb4458EL0BylmllyR/lgaIAY5jEUXGaCzyOGooTsC5vIXvQIQJpoqvELS88
ZPNRZwTcO87dg1SDv4UrVgv/AS6PM4JxVKoTsy+rDCos2NxLTKxhypBU8rZy
3VUKgs3ovnlo0XdNbK72QCLJu8W/9D3MA6nA6uuYramaF6G/3Gommn+7ycu4
Y+T4MKqCUqofjsvCHQfor79UwzNvPRs/lHfHoKBQj9RW4Y5QOj8DjJOW3dYb
6o2tFG3Xa4FPrakEyxQ0KfzRM9PSdww/TFIIJYA7IsA0fuXs8Op+2QpHMbQL
6+jDrkp3z2X5m+rgMzD4Nxyaox8knTvkxKJf/2ui2hirxNFapmwoSjOO4UuW
qoxayRT6yXz82Gz5hlOwydfnYqGZAMGjPbrRtWRyij5JyKmQEs7xitYnGinJ
tqon44CC15B3aLejLeX94x7VyvGOleCKCwia6DJ3Nht8jZQTVjyqxlpewdjJ
w8hTlRCW8+ljng7b+kwPnJi5ecJWWXWbAeqVx/i7eigOlptqz8fVGdvEYUoZ
TfUW5Cg7oCJcqvl/rmQU/2uCjU2KvcnKM6D3r4/Xl81kLMY53kNbgIZDkVtp
Iv+ZSKQ93NRq0ga/Vi67tc/dEUA5FasmxiYDCG5RtKfwl//X8Ny3/lpdCYqZ
EMxFizX8mJIomN2QylzvhwFviA4R64Bf397xO9UAsyzAwsIJqMwc5oEv6MK1
tr77U8oIEnFmnw4fv2hrEY5MNZkN2O0KpcBbAQXg9MpYQ/rLXindc6OHIzMX
q8/nt3VSrlrIn8/Q1m3nUQ1YXj3fx9z7ytaK5FiLZhpCUuwLP6PqGtWiSoZJ
72BFlZbHhzJkt5n7uztCWGw3Gh4GM+3788H4k5dCnZ2wWUse76sx6MXuDi+k
rozL18hSRLs8I77adBeTpUczEQB8B67t5A2juoE5XVdOdVYBs425G5J5JPk7
lAe6yV6/QwA06oOVRjKrQulMxZ19w7V2tjbrtcaiP9PFBhKIEnye5nsBH7LE
O4Q7lZ4pyyW1dRjBoYNKaL0lVIzCHhE9MsGZ1jr3mfcfF7BBKV+dQarIAd7Z
85QOSr8HTY2cFQyCMlTcZknxS8wJGfWBJWAz/oqITeoY9/e7iu1+Lo6wLJ0F
KpbuNVJ1utShtAnNbEwWqZrrPGrokoYiamKf0xJSXoHLug4e9CVy9O3s5sK5
GEh/j+0tye68vmY7qwh6j3msBRGCaHlaHwBqTBaW+tAjxk68KXYjT6gPif74
oRrgB6EOsq+ZoTyaVyOqW1g8XBUsdTqUQm7/TBEGVhQegJK3mCmlHORxsrpp
v/E3uOrPb/8CPGhDVtFBMeRO9sT47Chm2uDmS0EOfCrD0vDeNdlq/B/LduNa
+7Ou6BoyG0EZ3E1YJzTXB/j1/b7I8nFakfFbCJ7B0ilP8A3SpCxHc7dkWCIe
zUS2qtAW+dsg+RFtXcZSQrNDwRaxbUeSGVJSXGM3BF+EeIPe62ENJFfAbhBO
m8UHpSPEmM8oeH4aXAC4oa6N0HsAVWp8MtJNboG8ceHjTVedpiDkHLTiW+UE
M2HfVSWm3qKaL1gv53CsfnGUUNcqjtqcsHthDQrAq0dsqnjrGVbH/Ib3sMU7
G0ennfhlyZjlQzWVybxtT9fT8VraBD2grUVa4VXOzMw7gITTgsix/BAxoS/q
LRwmBM2jWuXaPD11Bh9VYzV8LGNDP/BINN4rh2ZeH8vy5Rk9ctKXEVaKaOhO
pDcf4VbkHvgsqS6FWSzTJRJr4HjqWMudfIDEnFfuDvV1LXHLrDgaoAlRceNI
LuGo2yIossvsjFxq347qnpJEq0eHAd1IBWGF1npVHRLo64w2CNCEXvYT0S/C
/DWyOD7n88uQqvL2ruzzUu5yMvEMMf/ZH/42/hgpou+Tf/DccB7752Gv/sW3
VDEfPzIT+grZDuj1EYKFjZb8wsVtb6hCal29fPTA3IXLRXHIGbEm1wr4f/xQ
/6ISS4jrIbjy9BUWJmTOlu+3s0Mu/fPegj25257hSu18b84q+4K56GHmWCVL
127jW1FtZfcbXl6AbXKVvttx2P2cG5Ug0MwCLgBiTvkWqvXViPumv97OgYul
ehfm/kZcvUqSDkgaUS3AD5cIhtf5uTOd9ZdBGp6xSUdeBCjrhgbbfi9vDU7X
i4r0wx+CgnLVKbkptBwGogR0dCUQ615nbpwiFbiwN9730DayOTCcTR+yNetk
NqJ/dCgQjEzzQgC+wrZuEloPH7B/Ft1bS2VhFILBkIdS+VvS3vl9K3nvInE0
slJ02Hopmb8BxFzeVUKmSvlv71qFmSPWVDVP0x9uF3VgTcp7wZIEobnqH5MS
+uRyRS8XH6MtW1Ri0hsR85rYpTqomRkIcU1j2KOpbuDKrydrs7a7L97s2xU5
W3Gl1w1CZ0dD8zYuP9UJOn3nGmiC8Z+itRsP3FrDrsj7AJcAhr0HMRgHB6pS
xP8UVvrVwOisPolkMFthkpyQHSnPeytTvlWLh9YNghtid/GDz0iySddTWWxo
mgjBgtv2Qg1CFgLfdgM7FWbebVLK6B05EQ/y/+g5uPMMH5xKn196Wviko9YB
sg+sHxQ+qlNkCKsQTK7NQAC423ti5Rj0cEbEr6aFmRiZYvJZEMovlx+cBG04
YMypQ2lwBbUzxnzFDQUiNbnV8LLrd5SzAV0RrK2R1m8+QUH2g4WSeQh2brdV
XVhX3qlVdeVfSnOPCL7H0/RnX0ivYKIE1BHYYsNJnVyA74bUxnsy/eVXS461
CR1Gytv9h91DcZyKfS+GQUM5z1hOynaDiZIJxn3AN3hk9SF+b1hNpw3a+dvp
teWMtUQBq0ybIqXdacYjdweeqdL1WnuMTAZJnwwsp+xz1aPOSVG/9tkDLT6x
4ZNGLx2TQYO+WWjt75dY5NIS7gSzhhbZJK1xUIf6t4O2M8gjcYabzInxmy2W
5a/mT81iPLSWfXBY8WVy6W35JPSJLsehIRWjepYCAP51cttpUcEV6V+iZQle
3+lznsoSjMuJB3OPhvrkljtGxnpZk54VLtIIZ2AmxEo0lMEoT5LI1kEvTX7f
PbPrjaQRQanujHChMkFe+LzC16jd/0yrJmZELOMECY7cVtsnLj8/x4kjTFA0
13xE84lBz63FMqI3Dl0i6G3S1xHPMdOlTIzc0SEeZay9qZIPYpleRmIqldLC
p+YNHcPpsmympK3t0zKci6D4Z8EE+J20QJDIsCDuYfLD2ik5tK9fm4YShEtB
ZLIdaHwkS4/G/ZP4iTN72TEkb35TDtNU+/89LcOfQWBEH+oHz0moGbCbpPfi
Ea9uDip8Ws1d0UU89P1aTd83OxghUXGXfriLw3jwyf1sExhD81clPyKDBb+i
GCKGXmkjgsgim64VYrXJZWxhylpfGtNvBRcefXt/D8hZj3FDlq/D5UDEDF5E
uoW0BIvSHw2eYMjBowJ3SLFGmKC3bxXwoVPbdhiaU3QFGF1sVGiNJprW8paX
/vrzavT+iWcalhcxN7KHUTDjdOseSwaEpgQJS2ftYn+DlsCOAIkXHvH5FJsq
zdXrFPbku4zpEAOj71tFm9UXpEmYzqfkumS10n3C7ebrnVTH4nWaZHUi/1dL
9eZHJlchfzcfP0v2PESFeRN5JsKzFNT3vHzYrNF4jWtB7xnJPaus1fLOjz0j
vnAhuADqYz1xNiGWMV8jN73G2W+1SLmSC00MMXfyZQPlwLM12BMQBqQXEVof
pum7GsfqjtproScxkgGnWUNt4yw90HW3EK/FEXMrb+sPO40qEHOXeDZ/GS0K
MqT4pMO+SuOZhdwYIOXEFCgckc8HJbBgVVaCG44e9s8firko8NC+jXfiUIX3
DEBKF+Qhb43d7J4XUpQV3e+CVJCkLOW6IOkhCWoVHIWzSJK0MI8Bv168NOxD
HB7LtfTDoL8/nCdW6aEDeBgKsHTKhaLNh0zs6yXGIv2NXxANbxhOPboMYPhR
zl9Z0LZ7nlrahyTb6ZRxa/pTjRpUJCeVoDMBvQcoolDL1erkCyioI8K8vWlW
B1VH0+EhOB7ZwXfiN1uDgozvMdg3FSbSJ1M10V26NRZtKoo94hk0KYldj19i
SJRJABeEndkTsKJ7W/YysASK4aJKtBqU944I1s6zOUHlNtWgctk1OogRt4lj
BBwLCCmwigt2fW1VK6yA7jbRW66AqPaR2sZmKom10HGkCXwwTavY6qYpXrJL
AjsY9JmElXCSktsH5DQQjMgDpR17n4RcBCOxYfz8EA7Zl+rc//Hf2ZhS1zdO
Fp3ZyxBzBr19FUfxQaHVyExUBO+oJdWBx1BWkiqsSfnbTk1hv5jp4Ybb0ciG
iL+1ndjv84MVmNLkq6GJVGBcfA8MHkiKtb1xWOzrfF8qSSmnxRSYzwRAwLck
enIpXkzb+G0XY0uFDhWFrk8Sl+YPNi5HZwAjXGnPliGRvD326OMlE90ObXCd
yD3ZDWQ9Yu+4rgUuX2u3Pm4iZdifPpFHuBrhED3rD2nT5ZkIX3fxYL/tDPZ1
MAdcuclMq5xFYE0z6sQ9qRTrtk5eptnWjGZ6lBw5CItWSOhwUPkgisFb86BC
d59grRh6ed96+TFrhRPaLfKZI9a4lgVOfzzmlpi53X4Xa/TkyHhz58mLrPF4
N3CjdZ1YEiTcHlsGiYw6pESSbR91UKPBMdLfyBpD2X88VIW5BMUMQsVu8D6q
4cJuAd4/Ws3Lz/6+ombJmYITciiyqBQG2tGcuZz4u9XSFebIUci6YZmU8njO
NTnH/B3IRdfgXVhIwOYLkgNG+MIkEcbaNKcSX9HuV4j3Akbj2HpB0v/CCm+R
Wa2CCEsgsp3MHT95u49KSgdr+utRS6YnzITIW5ztRMXBFKyjDP57ctsLCCbK
KSivKo1CHOZdOYjv91PKggpVz9AX5LRZmwfFIEtq3261LuOQ98Y6drj6wpi2
BLL8Mm05vPZSDg+qLqPyGRo50o7L33SB084Tj+5TP4l2Rv/rzlkKfDsrqS0o
IG+wSa2wsE8yxjqcDCP32cdhsRAeOsU4VATCiDPDYJwR9SWoeTBkoDhUVeby
V7vVHp7Buxy7dAFnHVEPa1JehvBx5eHhpXUrlDygmEeuYrSZdZRFWB7d4zAo
oxSVER14JpZg8b6p/mNetfIjQPwvOxXEz2WNPizBL5WSj1YBDl538w3qYyFE
HSQGyxKpG7TJU8fmoM0MHgHThDLwPrIc57063ZgeyN0M3LcXbW9Hbb1jjWDj
J8yYKgBgP9+Nm12shtkxF2zgc3OLgXF0YB67r9JATDpxJY7HXnfU5iKdivuj
MCD33+TJD6+/OeHElU7rSV8JY5pYsejdwQIX6wV7X+8qQzqlCx4x26DrRNwP
ZPEe1KTwQDwP3InW9aRTZRHXGvo4VgU7B6uvYehLP++H0exIC3/Rig68FBm4
j9rE8jhuFXt50PI1BHlVWXnsDE79ss6qgT/q0IWSbA2cSVLteyVKaTsDGj6k
u5phU9FzULP4zD4yJw/DU4075CK9ydHoS/OvYjMgaulW3L/7A1AZzgU7wEY4
JUPmnVV7t5ED+zTeKEec

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q60gJP/cgOAjJvKlql/WhMEdSU1bilJPFldiL/weegtPAtj+IbZ9D9ULnU64CMS3FxI5ZdgikhBzymaKntvxJyauuHNEpHDHA4hdAsRTk8p3rduBb5mWW+FpR9qMrrxs8eEEqG5N532ji3qcCDZeEc7oXyq0htsyZVW19mrvi0SqdY04aXadpfOrx8OKidMMc7tNjwr/eNEU5JOtnkY0N3hkAcNJGu3iHNl5RwD4O/nasJIVtQkmAH05Z6DFa1G2O4lQ3+5MoyllPnouYAYlfOGoZFpAztsIYQVK72LRgRyZq8IG9mI24dvSl/aUH3Bl0Orze8bBtpFZxHIwEykzeOaxJlNwZwBUBCqPqMs4euqlHwzZ3WCz9iJE75a/8fHoc5gUCBZzNIfvB6MNpdPst9Sdaa9H96RUYpnf2ecmtnN5bNdrD73FKGCWwHAGZ+bk1P8ZxTGboQD0w85POQbKKoogatv4DkJsJcACV+iQs/c1t2Iu29Ew+1ihFrJBpwBze1SHPqtk9DqkbFNI+a1tsI3QacfLyOqgdEQQBPNY7oV3lfG4cuU7VZjl8nNhQlyHX4T+WHCrHRbWvMvIxKtzF3rmRLXL1pOb2P3fIkhBraZxdUgT39fzXziOjhLxxtjD+zKkiH1ulm5sosB7euuoI5wwA0FaMWd8Z3u+ixrItJqHcEKAi6gEv5ZEohnZalACr8Dz4VSfDN7CfAu0eYU9ZO8KetFZl+mX4ZDxz4Fv4YLzLkyvS1YTm39pDcGCQcl/wlq9uIYk5nEeSaXEcyE8ZAc"
`endif