// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AuS9ifkIDLRvMugNMJDD4VNWr3lemPorh+z+wAajlLfbYWBjDoM4zEJh9jHe
Q8PP3hGwfFHR6a6W4DL3jo6d+1o+Ji+8WMuM2IZdZPg7g2JZrWFZLazNFHUK
HsnLlUZ0mDPLGqs5U28GpGizN8EbWtJqvuyTGvzZoqsEYT3YxDWugo86upIi
uTSRH9pPpZ1zK6wUKnnwOO1eYRrNdYS8wtu3KaSHuqtDBEuK1/AJ2pCrFiy0
jvVmnKsq7hf08OBlGiaUBEs3DoQjS+TFnMdT4eOl2y2/rp1j38N03br4uZh5
8mZ91us1gb4N4l+xpu8wrQc2nZkP2UPY3QCJcckXPw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Ykw8qmPWjmecftbO2GQyav9QUzgNn87AsxIY6mcDLLb80Rxq9fgwxfnwgnwq
Oldiba0WBbkz/CUS1mkC9w7PkJS2c9XVTyHCm3xLEDCuh5ho1i4Qi6eLpk3S
dv1djJ1VYEN12EH23yq7zpFByFAQMRAJUerDoYlgDAnhigEbRPajBnHBXMN0
okFzWk7OnYp11PGSFeqVXmhZKR7Y0OIMbSRHydGKVU+5SArfhMX87+epl9yh
30bSs31S3Jq1bGJWVHJEeNBGuZ3UCVbqUlZSf0jQcBY4jVePg0iinZTpCsCq
zdnwpoFkCjF833S+RqpydMNa5GX2+zIZ7wkSDQVgag==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZzsF2UCNy2YR8qzNi/p3ZGXDfNjBPrLqBGwQ92/P5zvunAEigDCe3HF4hhPl
ZgdYMnvlgTMvmX7ie2w1Lhrl/wj/DVqgvVyTmNfHEXotyu9Wdl7EHnXZYmL2
U07W85MpxnbSUtbURSUvSfR1JywNWTUIzuU49w273uKuMdo8OFRxWmwj4Zw7
whIO3aRYIP6H+gHsO2NzF9fatMzJy1BQVnoroj8I2M479qMPe3usWp8JDZge
CYQtEWpJU+Da/Q+DxQtoBzEx2KUkHgyl4Dkob0GrppA8ZZ+uNcaNAdcMGX2E
y0a0LAxZosbLzrbdp1/dqkKQuF++QnyiHHAZYGcc0A==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
N5+1KQqTLoxMl2GBiU9wzAGOg+sZycKRH4YnEICqTSV+w34OgjMBVvOrnnj6
9OVSbnhwidJLj8/75uLrtNGocKRLBCtqcE5WxH3/lPXTDV4um48Qm7feZxY1
T9XUq7j84IcigD/72qo1EGiyJry8X3ALBMHNWyEQFflynjMvjlE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XlYDeI9S/dAqwqcIV601/0FJ58DT1bY0rH9WvlYnbnl/W/wM3RX3nv3NDIJO
lx46QCs/QTVu38ZRp/PlxI73hZBZzYTUxYz74lRuDm17bZHn5jECKufd+ekg
HBBhZgG/MTHMQdoYLfRVsZtVde49hFJ73NZE3LqCjhG2+81nREtc9Wpjqsjg
pQXNs3Ek0cHPaWIUy1NQj4Q/wJd9wiSEI1kspNNduOhiMSEoz6+lrFFHk2Mg
d7Txn4veQDoHl12z8TtbLfQLTeG7Cw1icSHNDKqVa9sU7Yy8jGp3/fwKHotR
RV5y1xv+u240smKDtKCcliFnbHmekhF78vGbM6GAf5kwAUc2AOUKUPIin05j
Lf9H4UBTzxjsqNLVMdyJX8ksWIeRG6Hx+j/ecZTV9sx//GPE9gLHOlxZHYJT
nArhx+vUCZJQj6d2BAL/JO+qs4AMZSwWXLexQJzTTeDa4XU8LbIavU3tMZLA
b4h/X5njNjLuY+wHfyZt+yGqnBo3eYoK


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nxV2gq1kYljf2+l4DN/3tLkOPUgnQ6ua/R+rRRzxnjFcmUXlB1IaUiGDcVQG
5Y5wfegGl1nEV66UoKXwKVkcK+g/nlum6Wzceml8oTqEQzNl2THuv+8ogJQP
AMgJmq12igWRO203M1eSjtIOd2s9UaK/6PPPkE+RnYMTvGT7M74=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uVfHFycpjWTKEt2apBu/6Z+2mCvinRaD2T+KS360SukzlLhEbR+ameiuN0uC
njw2VvYxUtJNT8B4e1mbMa6oD4XnKzE9f+t//bfitspj6eX4TrgWT47Bhr6T
b2Ex1NAy5jsCAGTSSf4KUlThIsKeevWZ9t4vSo7pbvxXipU1iUc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13008)
`pragma protect data_block
TxncwEBxsHR9ePk+3WcjqURcSRWzDZ5PCea43cEoFXRibJcb7mGoGXEv0Oeo
S9LwTZabwsP9/LcSGf13793NdzRLkPO36Rx6NvM3fZ/ZBHNtVbURkvzMbujg
/WWiwfCLorOdEk5zlNuRXXn1bB1stHHvjTxE5O0Y4azr/XisYtdzis0ZNfBk
jsLus3B9T3z1ksGQIPO4qJZ0LVJSR/DeE6QtAvk9cFK6Zzf70r5JSp3HWBUz
wmFx2HnuFCvo+Y4OFpurRs44Ouwy42LTxkfvd8HqQ4i6Axo4fEzbHl9iXKrK
mMIEZEaR2J9YjWpmpOpoegIFMsUdOa9nnEy4d8hmsqJfmrhsQQILaetTI8tA
vzMcsrCOljLN8wujtJQ7KEZknGdb3Yr8I53wlkFCCtwXeCP+iLeMIXB9ZA0i
Hbq0gekVTF3ebgMtO4O6HbnpfqRO365xkBc0jC0tQRFgBgUO+d8n46OXIh+o
G/934yNd8jXNfE3pI1oG7zk2+tB3sqd0N8b3lUr3olxtA7xZxDXFxLX4gO5s
HfA8M1DxeknC7qX0yKle/xqQuS8DwRhxz1x9M+bx2oK2jUzQz/Zg2dP6eOa8
NLNH15LLD+St5d1LCBTR8RnOlqbhKTIKCiEJekNqwI8z762ScHmDkGZtT0vw
a2DJduFplO/4ccprDJAOE+JieAYZsMFTs7j+Ddpq0A6wGyIkXW6CYkpoAQQu
wsDikfnC26nBWZHXv1uY+Cd/m+QRDy0PSRwnCzMn9OPXEjqiVVTpBsX17bHD
OMOhTKPlP6HBrY54Vm3FTDSwWJ2C9zi4cAfVtuSNIZapzPFYb43Uo1h3gH28
0z/dEAF9LwHSLcb91b3RzpwNoMvdLRDE0Jo53oLBeXPpTWxDRt4LCxbZ1Ox9
j6aH74sRKNBIRxs/ZKDOMzXzMxwmZ5FuBJYNu9W6TO4HkcQcSAdtu2gRfX5S
jddPCEairY4JP+N0JlrJEL+rJNY+z1qFH3Vs5DWYHJFTfVyLCOy804b2cOzB
+7H6aS7ezE4V+uWs7237PlYBOwZdaG33/Dx1gaEkASWlTN+Z+uic50zEYytK
uTzfyYBWd2WAY8B4WrVQfiVfvrmd2mvrCMFvoT4x3dJysb6od98K0h0WXSZL
lO+09cvWPb4JxBFUq3gc21q1Bj6RpnrVCMEc3YchAi3I9lv7VYsHvXxxjkzU
JnQxbY2ds4JZZKbSLrcNm03bq78DPWw4DmI1Kns2FNzkU4iiVCBmpVaJCqTC
lQl712HYuR5q9kix0Mblt5/UwG1xp08opyAcHXteqjv8Ob7HN21vBtUU+nyY
vbwr/mpe27RyXEbsLdZ6G5rPfMTnVkhkb9L6KHKAYW3Ujz5J8zbvzuHy61Pk
ff/Gj+DP3zPbJ5rZ8SZG5Fy1Y+ZOvz9sx+zBLFd/dWvU99M6VPoBH2VqCOlp
sAe+so7lQHYzx2BzK3llmXKKiIMffo8hn0oKwYgorVLXhHnakezCmP5HmIcr
NZyN7cE41AIlIRFI7M97i6wXbZusfPJP3BeTeh10PpcCOJmDZnRPyiw76Ktr
+EI6HaAPRieq32y/qhaY6GPoyc3414hSjOktI7+/HmdEVJ5h0zmJFQ5jjyKS
POok2JFEfl2HgWfRAS/yxlQRDDDlCXyBh7zRzDSFoELWdJTGv2VEknUgMJ7u
NxkHEkYmDmrHcgx/0I7LS/1dSIiIM2IRZtwTxYzyMH/pAmxRR9IV2iWtQOOv
JgqpUkx0XYU4BNfQdjlrEfPevCsDlS2PgZpDZS6F97kwH+AoK+VLucCfj5iE
NmiRaMC4RLpQBNGWyntZcyVABd2RpnjGSXfKbVyWzSoJjKDBWlKBwpGWQj4p
0VAgUz1yxVFMZEp1QAIzFJGST9HkJK5WmBZh1dgmIPD+NAwzX5gH/sbroyyk
bnBDLpFGnrkMXe5q9GWgmr6MO5cLENhOMnmavjVgJWFcFBDjqAEM7kqrVhUD
7WOxXnWf2bpgOFUm+TsDCr7MSTCxnPt9qD2m92HUaqe84Cjrn/8fmigqEQlA
Y323rvs/JpbVCgiRoertsmyjSKrnvvwbEEopOtHWSe23bNfnKe7fglRu7ceF
MKA+ZTFO/814om2L7DsFzkyYbezxUkRAK4NCgIQo3hgWMsXaRhl8g37N39wZ
DAVijR7/T28gcKzbhrKyIhyvwiMoC79gstMMMSreDJmrgiD0nOffYb7v9xDh
8SMPyyO3XBdJ6+l/jolAIlDHyTmiIUN2DjJmQXgjqtzAZBONycg3jTsLmA8y
7Kc9/05wakqfoBwwKcIHnrpmny24fwMfU/rTn83jAsi8ZbvrDhtQuA5hCyp1
PHWY4aQkUfGCeyGuN5j3roXQRXhd3gS20VyMf0j0BpS5Q2rMYSLPAvIP1xb/
ntEVtoDU2kRVJdVBnvpPQ5ZdhzJr31KnWRO3CXo1q1EqZoSe0mCZHfqC673w
sazADHSF2h6/egFxoCQdP5Bz8geZclPQEkBRIkyT6tNHEr8ih2TyMLIiZ6Hz
0m9eF3n3QTbkq/SFSc5/6EIlblloMbLd1etsqIocmJdTzjPHHZhzD0xUAy9u
w9zJNahY3T/gTHa0QBTBkYZs3TQ2RyRIecSDYDDvFt7N+n76LN5C52c3Khn5
qa3f+96E/bnY4APbBxxID7FZ3YvTTG92oauz0yaQ4/Zg6YOcAtek1g7kyNt2
asBhgtsoPClclXaWmnOJM4UJDuIcW/ApJk/tKtrd7PZb3MLvsyce5TPgxP/P
7IxMQ9FePEyQBhpbLsJP1uElbUgdHh1YVT4vgsS42VEeJ0X4wCttI0CXibHg
o/IU/Pnyba+HvBva7wkPDPrCtPPN+Rrn2n85/l1NQxnoyMxt0G1DTOQMRMUR
TJUvcMT/6lqi5KTm+B7wqB/S6MjjaaLgtmUC/mNxfcpMWsl6LYq4Twn4JfNE
UDTr2YhSpT4r6zVrGlZieSUW5fIJR8/f8cPX3bkrq1G52plRSD+/51oKnw6h
iJ9AJT2W9zoQ8BZv0kJrcFm/RV7qst0yEz76R4C8wapo8kOAbVQKE1SLWBlF
r2S4Tcj1kCNOLqblFjUjIHf9wkfn7edCiWO22mpprAekquoBzhCExoQQq8q6
DyZGh2fFSFZBbKrBslx2rWCPHFqmujjgNhLLgrg/38PAAhnyVmPTdqfhMMmO
Am4qRdC+7H5upmSy9sxL8XWLgJm4Sk4PZPEiO1srS1+N7yGT+JmYblY52Q4m
EbPr6bkdjytHHOLMQjxwCbliSMjcPTUbS3x7eWod4dIhzAQW+KQI1BfKXyfn
i/yWTx+KkH7KATGua4VneNWTi7M/c6e1+INYRvSIjt0QZhYPdbge8UYpYu7+
QAPV/SSfxn+EVUKTvGMkD70RCF3wNMhb+y93O8EYxFnm1QwKIM4bmCW9JxAF
wbrV2J31Hcyw6U11MXa/C9B6ctbnLkV/uDWjtwyzty1TxBUCMvsPzo70acum
qxuleWGNF4ClEXln3NcaPhNfSmqV5X3fxuw8fys+nLXzY29JTSkM8tQTmB6s
klvXln2+eeDUYgbPVkO8SgJmVn2TIQ38H985auoabyfJFz8iNrEK7hXlWNd6
HXNMhRHn/GDUy3x0YwZfDPD4qy5Mpe6MNw/sfqu8+pgb2+AZsVu7wRtdg2Li
/tQC7U1+Ubi0PhdTcCf6NJxu/OPbGxzXDK9ogD6fLgVmJc6zDT0ZC5A4doVQ
zNgcQNEPOCZKET8KGegmRh3S0IlxaADE8A4ifdBuqztLQCgqlwKJceq0GK0+
pIJTsaIUqyFYR7dl9bEtrXUIHImuoDsE8vELQqjhvSWkFi+jNYQeO4ICtM8z
1x4ShGtnKMPxdnUXGpImg1ZwvG1sTWItTvJGpt2e4k+Ft3fRKRNrQXOVAKl/
XboJBnmnqA4l872lvfIwBWR9HxokZ7e8NXDco7PaYWvXOLXgvWvNZ+DvNPGi
aEJIQfNukwHG3KOoRFMynnplradpp6cBty2vCIdLZvG1kSZQrZS0OTwLpNmQ
z1Y23QbsW0Y9dbHYAMg+fGcF5KzCedx1qBC0Knh+qrR8ITjlJeRjJOF3snw2
mIlcS5idkqKipMcdw0CazyRvt0gcySxVt/uPLE3sIoZNTRe4K4pJegPjSDq9
OMjCPl2YAs1jqMWEseA66Ba1yKBlC+vk6LewnNy0iCI04q6ANwn/qVHUCIHV
QAqMG5TyFZrwmqok4OLbQmSvO/+JzCXev+woCc53GmQmhp93qmmSLlz6N6iD
px4kLdnpXoGTbV/f3WVTDvBioqYgNhZt3wzVRYB7JbNeFEhHTxa/08P4QC6K
zc+5X0ZdKwMZ+gZpX/c6PhHihwVFjy2GXZAaVtMvbg/0ggQRKEtBadpS7OTG
8dEJdPeRvObqB9PPLXNWJjsvZlMf3fHmx0NMAV5UP3DosZdpH6bgqapcxISn
F71Og6F13cMe1XZ2dTEWKKL3vMjweH67tVMTY4nRrmmIdFXfN3G82CwU8F7H
lU2FChz7iwOZt0VVb+3g0wFiiZOzOL+aU+/+RSWUMm5oOS3sMvVtr3CUav8s
23b74Rw6nGfg4GGu9k8Agjin2gQN9BGrRRxU/7wiJOh+12wkTilQ0b2CJ83N
zzrv8bhgY6UDjmytkm8fRtcNW/p5X++0SlD15Ps4tRqvePirFG12DVh5za7l
k2621Bly4hNlfkQe0+/S0pGVctZtayd/eUnvsQn6TGGZMxU3ru1f+niPv6ir
UFml8IPVof3gFGATVExmSGRQU2cp85H3QeiebiVooxL5I8D54n8KbwVf8DFd
nR6/VWRu+dPT/xCGoQmTd8Mih7YNRGOaXyR3k2QVy71l9hQ9THeC7J4yNHgp
V+UFBBD/0kTKOY2tTRRSavCxXHs2LcihtkthDR+dCPNNo1Tl7xHHLAaaRmkz
9t3au7E3pVOmVTCgNBVRcmVH0lOEw/6lOVUtQwH5I0yaTXRgjx6dI/trSRiu
Wa5DbDoCqiAy9crW5aJZ5gSBi1/FHNGPVchkothINlrAmZtVMbDPZ7QFj7D8
J7wH1G4XvpT6gi8zkIJv938yURduWOvle15UfDJI2hdCaPHpKk55DIDkD7VM
oEtsjju+NCkQURSvix717+romzOhI4mYJPVXz7UhDu+O/mwVLyFPQkxJ+8Xs
38OvKYmb0EElld95NdQ5ngGqsrPzqzqVYy3I0p9R0fPhs9wTNhQWyVx/ISju
1lUg03iWP5A76OR83NzOSExpW9c9yBlPdBwzsVCWzNZjYnDox5/u/YzoLWz8
jIIsUExZi3K9MZRWsgWW9ruXOOSLp3ghscsGeozuqOBN44SgboHvpYT7ztaV
Pkb53ZH+T+Sk/Pa+5sIjXCW69Z8e8bPe/JkJoDSdGB6o/5KZv21fU5XjbDrv
tL9gt2S1hPwohIGWeLONLiCqlA8zVaWS20cvOor1/hPe2FbZVIDyBsB49YTD
iG8J5Vpj2+YsV3nRQ08ocV+nn0ymcDwgQTicn7ysrpv8q3lY8uAW5fJL6Jqq
tBELbfd2bAafop/QSnLPPHZ4lLIDevwIoh1B9x1chAgsOllfxAST5Yn7oXKs
xhFwOS7U5iQquHE8lLWz5ggif6T5TvTi0tlHbFuq+oFq8bKvMEtPgf9q8g0w
1U6vpM7U7+garc3cfowmcOoAD3NSCpKmLoJmecb2zraDhZNTYqFAjDay1HMx
q8fVlkM+muGFevj3YmRVA4SnlSlvCl1qB1uUNOA8Vet2COOwnrFLLFul/yq+
T4dK/xdkwmTw4VI8PQbIv5Rz3aX5M9wDgbjzJjIlCv2A3dUuj2FkrN/DGrp5
tSwAkiy/3q4SOhOhCnYtYdoABwoz1I9NWqUJc67yf3cr0sBaGzuiET+YEWPq
2XuphURNxC5/8GChSw5ZNREhgbg3tCNB1giOjnlO9KIlHv94P3nlDH/8EqJ9
CFEUistUVDPbBrsvVUSksANlg2nm76SLUNVwL6EvqiE4duH0bqHlmkON+Gsk
bc3kvAr3gYk2t/Uhs4OkWAUu4UPvnlBRkSoZgCooEnCZ4keT/6tomLbREqhG
kkqCWX/XqwbamMAQA0pcc2la+ZcE3J97x3/IT8XfoIF8d+xf06ec2TfPzB0J
qWvUHOKUNtLrMsipYkgsfnp5PatWqQKGWewAArWl6sa1ip8eH0mUi6ErbexA
6ndTjF2UJCqCuy78uIvNy6zOtKZSdv3OOTGTrvGoBKso0SaOCTr1FcqNs73M
wJzP8GLiXAO1vowfDqDc8C6pD82b1LwyvbG6pUbLltHnRmu4VByVBZdz9D7p
06xqlfQZu+VO5VWGLWqurkI8Xx2FZNZDROM3qXoXiuTHSiFA6OU8dU+WmhNv
ItVu76UhvucWkpZBAAD/6remNrkCGYHFRKdf2KsctXmqKAalXdOqFtvbHNR0
9xseLkL/FNHym/zV9j3cow4iF7R6bEfcOnNYffKskaw3ecv/IJdv7OhAhjC7
EeEGdmvISLdIEwFHkD4AUQfHMBOrh7Qi7y1KKlM0Yb9FjxETR3nk/moAjCIe
7WruHA0mfqeQeg4OEXRdDBd7y/J6avMQs+z7iQL8CAhx+KLRVkPJvRS+9OpH
FUuVncLmzgueK+VevLUd44w6Rty1/SgkG0AdzpyqfIWu3XBnktFUhuBie1nw
fFBt8cH2DsRvhkqpdOlaRzumv6SN5+jovXmCk0dvWkw4TzW1PrpflSlMW/ZJ
K6iLimc9lyowYGvkyoPMDMtEUdDG+bYdGey11pw9vkL4G/OdsFHkz6Pl/ZI1
LCzV5GDrAmFdnFHNrAHHvO0mR74pJRNAKOqTR70mgY2TOrVmoqbxl5dsbm9s
/K0VY1XzcUZyN/Jc/TMDn6D2m2wX18RHExMqah6YWtkp5e+H1gsrnZfAHlbn
a5ztVP5SisnbYWyiB6SOo2ra+AEAqF1EANngbJpwLCsTgZmzxvCdATTXFqvF
iwpl1hzhaHmt292PXUnRQIAlPnglnjIcQj74ONNuszyYVWMBsO0Tdv/i4S3s
C/Tuq43hupJkfBF6xbgQpdxs7k+OHFvTCXEn6PLn4EaTa/6AI2UiJl71zCnY
8JSYORnOKCoNCOjyuGq22SGF7K8gri8puilddwBbpHaF64uxaM4duk84rylB
gC2lDnL0nXCUPDhQxdzS1Hg3aLulvNO2i2K9eqJ3sYocwQXiiXygyDYU52fK
iRaPru7+T8VwoYMzei5IRHyzW6o21gQ7x/3AlCxvbKiZP4HWE5QMSSMscW6s
Qg4R4uIPnfmVkGn9xZsYbxiSK7sfclswlKXX/Oz2xTxso3hMXWm/xDSsWv62
258P12dFwPkSE9pNwTehHNh61py+7KHSiQIbI+XEXuy0q0vWqlpr9NFCMx4w
UJAobZKygIil1nJ1EDZAGHXLhR1RcPzL6H1V43f19/4oTQMuoyGGBEPPsdXQ
aFHDCaAhCk27XDQGBRu8xOyrdK92NAHh211s+ZCOgUI/i89WHFB4bgbLXlCf
kuLHTjL6vbFKeHTgGBAZ6ayna2VhcuyvlHDn0CGVGeO0J9NwhYsJhqKQKjKe
40GXj/QWEi2vZhGVQfbi7S36gTmBrG9QL+7dxEE0KpqSN2ea0vITt/vLowf3
HPj1dbecrmZv4Aj7QPF9b9KTU8XV14lhJJ8RirGmsqeV+NWCPLNNyVfxTtLP
XhESZSf3mzw1F4dWpQSAaW1hSuOcuFTjbUnlhVQI2zZAknLEv1XXKL9CMcdH
mOnfJM9UAvWIwHXwV2OdAoEEMbPz60Qfj0A4oIppwVWYq6e8OrM/XcZotKCW
DU6EuLcbKGbNTIb4mOQ459k+rZaefo5sOd8ykZWo7Y7+rZaOwlYTlzEiX891
dLNbui2Sj25wRwCNAIbli9xG7P69AwboZV51nQQDNDzZymuy/FMYFY3h0rQg
xtsAbTLaav/RDbB3NI1gtyHkM8kAAsInie7n4EcJpQV1tn3xH5hNS4dLBQre
1oIHrX3LeEcMUmyPmbvoulN7S6Q+RtlnLyCfAHt0DB7S2EaVMSnPbKxzMDVj
SckXJ7naDyDQOL30nISRqcdWCq4t7M4XV46b74FgMIa3aE9MhPBLWRDW9HYV
3z0879M+U55SCJJ1iUteAaFMTVIKdzbyCUeU011+hHd7fYmpLErBDhUvftie
wGN91ekUnQy++Os8SgSILK/EsqzEGuNvLLg+GfViWlqoGtOB71Uo2dPpEIp+
iJ3mc/2aXzlHrhOyCoO6XYucDrD/+UHC1QCa5a5blCcxo2Cc7Nh9DOa/2vFg
iSEc3FjHng6CgqmmblF2PPXKFzqiChNrvcNT7fP1f+lGB7hqh3t5Bilz7SZE
EyMUV341HyQJToICjg9Rji5zwT1HILcjj0A+p/X9S0rTFORJ1ZUhc8wi3SR3
2wBkGy0DsVOEWdAV27nu+crvCzm77+m4Y1gibypQG3y7ay6T6zkHKgrDYKrw
JVR4ahKO6b10txsgDZls2re5axF9MQEL9NmTH+jOiLTwKZsqyjb4rCvIswer
4CXaCuy+oYTfE/njkNohZuy+9cqVAfFCD1+XsNM4SI5XLkkocyq6S2anDpRc
nO3s1D4SIeJ6zApl9vY7ECHuH+aGv4DJtNiq9un96YY4/3B4kikW+VfuP7OV
LjHlvYWX6hzrv9Iy27A4jKw7WAiqDVodVDrSAFZcFQE1HAvfBpi/Y4OM5JpA
wxwQZ9rC3C9QDQSnpwhzxnatvSF3UReaFy5Qg7Lv3e0DK5vAnVBhgPyKlpjZ
nPRGNr+dzL29BYZKQ7iwWxCXEi1H09EiU7FWFEMbLjYrvYqHlO9hAt8iIHw5
G9ivWApquwL4U+fa9SrPkrkiljuvC8xCNxXHWNidJ2Mz14zFKdvf20zzMoaI
g3RVXa6JFg+BsDqyaZGeylf9zSee3230INOMKvrXMLht3AVfdH66QCByYdpd
PyIKv+J+E6oVv1GlaLVROBweB176Sc7itCyaXzsZlMZiJ2RAHfANQJwQ4rJa
dsWboPA4AFeDN1l4nLnw4nFU4A17pKARSTarnt+G6/8gLSWCWt3NbLdn2RQr
m4rmKMVefBfQsERPrE6yD+3/czAGlFwuXGvxuckwOmhct/dgPHdGUddJP30L
gkdt/qhdrdCSenfL/K2eQndikCAbNhn+kcMmDM8Sm7FlpVCQ+z9rQ5A5tmDT
Vxq7Ny0onjiZC10DnTlqWswveOGKLJPW9oUinu573e+mh/+R39iqLBrDzDDT
NVRGvr5W3OMP9ejR6F4PhxzrkysxEIAaBveon/tbQG78EeI+gKP9O55YvlS7
JHKq8iZG33cRWkT7FjV84ch+hmvKEcSAm8rdgmRlIPdhcfWVbEIjCRbM6F64
CcxvmLWuVktha9p4hqkS1G6mDauj1TUnCWCQ0y83gus87NOHU3OPJjmbwPWj
+y6PYLZTFtFHdLNaz/2yhu7DPz7iHYgR3arXcHtwjlJUVzRyebDjEc2iBKXu
4f4h7I2Q4ulEhxJT31x4t6i8S+ytX0/ifODbTH+h0Lv4pz1s/BQeYlfll2oh
I/EXEB6bRWmm9sxnAp9RjQNor9NmHL+rOAuKWdNlCEPFk+mt8Q6bWpSRySKV
yPFX4LMU9U4hIVonThqiaX3FBiVjoHqU0kKWBvwiAJekOh0Xv5uyYhZ2pTVO
stRfoLPhYHpEpTP3745x3yC5LBKoowZ0+4EZ1T1ZJwezNhH0TOlnlSGiMOi9
9UU3DaGLgTY9ldZdgYlSvqK5lZnjMH0avcBXQ6+qLWJkmXDN83REUFH0gPsv
MieQUEfcuBJBFadKsyep+1SrQNQvXEEnHbzZs1o93MDrNVIAidf/TrPx83r2
HkfMiQp9Ai12bT1UOeiYN/c2kQKPnSse7RjrAJeOvbe5W3HVUQn9j4Ld9wF/
8w9vyExcaovcOnWslEVNOqIu24rdhZJq6g1FR9xIQbjULgV2EfxjR8vm0v/z
380hqzOeyhSUavSW7k9N+Ghr1Ck77UqobQKnFBoFDjAPJUHnjk7+4XC6MsAV
kQfQfTDCEgOV+clDhZpYKNyir2Oj1R5hu4gt9cBcvbGo+WeVQnbXPnY50S/m
KrfVtjH2hj8hs+wztS/rF1b/ubrHdkUkVvrZYAFWhWGHVUiTDon1QXWmIcxL
AHz8ixt3/UsiCRlEOQJ5+6TBtDzC5o/lqju8e2m3Tq4YEKs1ekQpg+No//6S
AYu9xpwQgWuv19PHOXsymAexvB9qM6Mlqri6JP6zWbG4ACweKkCXprlyS13y
S/N2EQbGZnQvPXxp78teP0QMEgoLPRLJlMVmUfwG4bMyzBWawmoAlHU5aZNx
PurayRED8WFLwb0F6BOPBAuv4LG5JgOudAhxvFb0MiGdPZ2DxgkS0h2dAJbH
lBKTfZI/AKAmEYZpWzVy0ctUUvluEDQ9Nw38MKADOnQEcKJudjJVATmC0Quf
nxRyDi39ceGQI7hFYHfkCZ9575xt6G4SZxPl7rtXnkOzcJxmc2GcttUM0v2O
vVpvtj3lTlY5YtitfA47wO9cvSh0/VEbP1VZufFOkEcNGNf+yQSUydXtm9P5
Q12D/IFUUU3b5LBufoSG7QFrS6nrXVt9U6ne+izFPpCuZYun0rSbte/7EH2B
TR8IOgQ1eTN4T/Yb+qPNPI8YEJpmvSk5zsA+MYeFXkgTtUtWUzOTvGe+x01r
Y91N3/SWt1cxHiC6UU34WPjwohZOUJ8Q7Knx1zTXCtZQ6zNELEXuYx7gi+Su
ZYgalC9FNs96AnWpxDH3D++ke78qTHCvb4cZhuecoBJ3o8n36x4robcaj8E7
aMJfz+mhd7uwFKVwflrjVU9EpfapRWmbH957GlzWVD8Zy+pthU9KIgS4husy
qoF2/GlAKZCoub7hYI4tuArMVu0YeUdmnx+0oiejTbjUPK72UBpXuFCwzl50
kYlBKQDKpVdk/5jPpkEpzcXFeoG2frOcwXDKZmzuHuFxOE14pL11WWy0u0Hw
3SFhZ+xIM52adYVO/KoIGny2+1Eplj1yapQuEIBDoj1gU6h66JTu0aOTATbG
A7KOSX52y2pf5Y+MfFAlqDeC2aAdF0bgAwE6PchHEdarQ17z2JW7QXg91WrB
ZkiXqid+FYh0lnwKZiqlW7NxtlyMGy0OqV2nWNLdBXwwwdkjfz7DUf5TDatv
hS+Yk8u3kF7KBp2L7anD/SRQe41wwKYXAtZyBFKHPMBoA3f/fICug76mwPYl
dEXGm6eLlFFOQc/wAQ/ghJskKEw65WPm47JbxCxKYyRCLhYPozgotpOomBEf
lhqg/xJ8HkzRCE1vu3wfkGFRbG7F59GHVUWgfS9ADXJ05NLy5nF0+bPksfyc
TQKKRSVSR5NDTpYcx/6t7Jk3eDv7Vlp5iG1JP/BYmYFZl+FAyrRrJFgRSNjh
HPKIVK66o0os5H5TvqUzgVqUJ/LT99fBFFsCthHcYGswl+x0ZKWOnAmgKZRR
6nvVhPjcD8lWF2if3aSOl7rrBC0hhj/V2a8qZAqmI5ktNTd9ntNRDV3mDKfH
rkc2NaV2aNRXyiY6QJjTupfeGfWft3Eeed2a5OAZ8nZAn4x8cEnLleK0Q/bI
LSFh0sAcgRj1G9QsaOGKZpbf8E/vz++XVghE0jb1nWomW0jZQfABC23Vm8Qc
zIi07HEca2sJAoURx5EH2Z9QFpxE08pmeagtHWWDWhi5MDsarC77+aE4T0I3
ZgRZ4jPJQjSaTF5otwj+cSQykM4r9EThgneKH3Vc4wnMdZd5ineA8YOCnAN0
1MKhSGei0mJhUX3Wzcr4QRg7IRnkPa7TtA+xfjBwsgQ+NONTeTmFvCpOhefD
jydbtWY1/QVKuuXP3cZbKgK5mepCoQP1dmk9sH7E6TVXAJP15BOHkpxStl5T
5TALMKFbkXRlZoSph1p3SS05OCfJ+a1k+Z/2PHY95YtafWGMO/Qs2F1sP7tM
Bvc/RtLMD1XcBoKaWDmE8z2F1VHj7WdOD2U7tKz8Aexip/MTUpXnPExDdHC+
MBDN69mhTUUgQ0KPVcNUiSAbSRDn2K6XIjH0KXWtIW5+TmV2Ryq8Mn19GGeI
hLDgOY8hBCK9foVY57W8M5JuXBxcAbmxtgB6VqvWih60YPk5fd1//ts5a6b5
wB/2cCdhTVp4A5x496wiK6xeVJUiia8ZeIYNwZ6Zi6AuhZtl0MS38l6cWYiA
kHYBxA57Ghqwz9a58JGUdvYh1sUyh02uyCy1Uf34y2IDvu6z0hWIwqWLTUqk
h3brcytrF0T6foMeVVMVFdaMYRoSkjuCzX5Yvb+/OsrsZIc82Xu0vVJ+Iiy4
WX1J7GkzgR3y7htKOevRwNPOcV9fm5eoo+rNEBFf+DwmtqPrNKhDvSKMjHry
RnLXyiRZF/Cplm79bu2i/Q3cXz99yOjbEO4R8nK9YMUfMw2dRc7/Sa0W1bNd
nh0dOtFfjSWBbr+UUWIbWGDH/w+HhIFH1Rr8cNn22ElJZF9YXIpFesiTrFfy
cgRw2f9GoUyxEG+Zy4XxtPXPT0aaAlUfuRaguDADR2E+6DsIykQoQt9l+b5b
e9+6aR4glE5vFcl2Gw0YHdo1f1sNOWJpDAYZIeYjcnsDc9pi2ffwuLnrkZwa
LMAHLfRSzRvsv9iE07zSZdDfNCIGwQaBu+Mm030k1to//uLl2Tsa0+53VzwB
lFrQNEdv5pX4RvYJUZ8r6jcM7cvPqlJql8DEiPjIoVud/aLpAuJyMJCoCqNx
1rCTe6+uz04rsgFOpuW3Pa5Xqvo25X4eO8Km/5BypnJet+lJMbUilaTNQEaa
a+kWxo0wlh55c0MuEgqPBl7uRDEKeuU6+tH62PnAamCXzn1HbXGHqpYntQ8s
r/w+zuRuW7rOb7jJsMHIxEVoW/n6geZoo4RibhUyK3Vor7vTYXBNd9wczmjh
2sjco7i1bCU1P1bIY8U5PzUGehRmSvedcT8XrJORPlBIhsXVP//La8n4INxr
oTycJuFwi41xwAOK0GDRZyeM3v43IQwS15XgGGs+lh79KbAAz5v22a2saWjg
fHFpZNVM9pyvBbMZ6zSe53+JSdrGnO7tbPoe5kYOVdJlNVjr7BsTHKrlpFmu
ND4wOXtptaKgDLqK7ZnHDehKrmp+xaJw8GET0y3RMkKy9wHRYMCsQAs7pZPn
ezpzn0wD8ob5+zVT2r7cR6X68WhY3REvrnemyBby97Lj+2HVFHSKUsjE75ZC
mA+S9+qtlEfGlO20HVDeazaNmLGgKr+XZx46GuFl/4aQVTu67gK3Rq16DpWw
0nnHZGma0OcvmMcnCuAJ8b8/eLZDAuXPp6K+dlaonWseff6FzIN6ffPpnJEw
GtrDWfRejH37NyDPSihmGuWrlaHYoirVa6ZtXtoTbnmhkUEBQDMBcrCRHSST
r6LGj+NfBt6Bn92iilyNacm1YjOzQ/UJhNlknujwIJsTZ53ANhumH3Faopze
XyaFYRjhozCYtwOqPGcbfZUMP2vDssl9qOZWsFxzgYYPJetyafM80sm6pL7y
ZXfNxM8vAeERwWFP+ADYgsPA+sJvXI4y+D2FBxRAceddjc6USSjDQVmgEyn7
y6+CAyPsDCNAeGZk7c6XvtW5Tq6TaY4Lnx/+6l90tz+Y8gtClxQgr/36zzQ+
E3Qv/Kx50p2ouTVwlJQQsDQAFSB3Ce7H8c3+u9m4Nlk2X8j3bJZ/MgdZKREA
FSwQhIk8LSdP5o4Xtuvk+dZikMLPT5QrbibzeO1HijpdlwKYATdCPhZ18Jyl
vcpVY3OeQMAdJ5l88PWka9FfecIuYPQ30u33Ao3MzzHcptTs96UEN5AJI+cq
4UTQf8r46r7E7lwvx9dilZn/bSdHBI8w59HU4syQjRIWppB2+jkUfGOfWD++
dt9uci+OdkE6YIm362mS3AqFdRxzrfmtKJcWxux/eZ6FnHn8TXX9gEc79qAQ
yEv4yzMG1F5KTqyY5CHjJ//6cDeaJr8NZMB1mV4tYwZildXhQr1xiB7TaCOJ
XcLOpWKUbLC1jjVzHSRxfJLFVscBb7KQ7wfKO/AAZ4Lyv5/89U/hqJbCrdaf
11jjU3kIJFZYpYBwQLb3q+RKzC185duLwj34P6x8uDZ4cj3TBk2BEfpADdu4
neZdApZWCmfyhLRK7OFaYSicqX5+rJZ+wQCDoNqyKLDZH3lXxP3rA4zZ95Qb
uWNWvf4dfSVw7gHJiAk4XrZ/zZwjrmSjsLJMTFJSIyGPLY2cgKLK9/GDzL8c
sY9UzbaF+aqsCHYpdJEctGcyTADp+DXDh9yGbOWMbcjI34bsgdt7ezR9zVvZ
QJl4lI2KDraNlvCT6HvC9Q7137Ni/hiVQPFPzRvxXE/yX8RNx2iASIP+B0dV
HfyCmP8onImDPr2fAshYF2vok1xRpV0m8s0ZEIxFVtmGLZQXqDKpbNFlgyKh
iQMJijKGQDT8h2b3s0iY+hpkfmEICpL3acy6YOT0Ex+WtBU9klvRsYgUoDNc
R60peWSZ/iUnlsNqwnxiRhEjZWHtxG2tbCXVQwRVTOv64HCgDIBVlNlmBbeH
cBPbXWQXfNOF1RmixiUlOfA4slMNW1NTgTS6BcReF+0/w4DPycXNgackhB40
00RF7y4YKoyl+GXHcICTNpm/g6n1ZXT5cf/wqrgsBABdmfA9xoPW5TkoI6LH
u4d/hkJHt6rjCTvD8+OMfK2psP7GcEfF3IrIRfn2TU+//sh0qIBQkZmLjDo3
eGLMAW9AhlZ6pBdamObIU73vHFldmKGbDedFUPArY7FQebAlmcHSPucqT2Kx
UjZ5eABPcjVxxpvh0BnmoBHyPFpAE1yZUci70Vlq6gCYOpasGTxqRxO3GshA
ICspRXHjeVG4y0ikEsfXMzVUlxrfJrdO6q5nxMFwIckSm9VpA7lTGyztLn7s
KuH9VybXO+nnM5tOKa186MZ+RIDv+ov1iXUcuQ9yMa422kuwqT3/14H9mns6
lhSqPe8vWr8lVHIG7WhTTGFJcPABRbrWBaXZpzwRvNLX4H7aJz6fBPNLaPnY
sqnLiX6ungT1U2MhwlanNpjF+LHhfHgTRV98xfi0a5wiJ0KhO4wkDtz006xu
wJiyYHUJpTWe4wgJ2vA/UMFcjQl6q98IH5aiy4izK1CVyJMD+rPRNR7mIQAG
AcFwU4b7ckLhBP7ZILQ7ljO9dMqOxnX2kT/9Lq8FRk8mxBlYICr0MHZsoZkM
7JiES4NvOtrmFebzm4EOUgmATepx3PBM1Q+PnBG1FpD5t8SdEwzu1h8+u4hU
FBE1p/mm5F91MeTSAV9qeaDfxT/ISbmWbz4dcYh6uKXRWn66ZcsdCNmXIEZA
A3r91NBUdDsVUrLnTD4TXyh5+NR13oiOcS59Cx33mHPqCU1H/BYDTpBLJ6CH
hbZSFHzM9K9pp+5n1YKj1cmwWvZwtTjIrDuukGfFXkHG6SifcDInRBIZ8A7n
VUtCL2m5wp+57V+3OQAQoCb9maj3zIA9dmLXkqrEyhOVtS+GuUs91HJ4SePM
/gAo+B81FeFfK0tUHoxdBAQtBmaumT3T/1eF/xQeyNkUWiq5RVUh+TNU0RGz
Vbr130JjVv7V4q7g0wNi2CrEQDFDQRth/UP5/1UrvVDJqLjqKObm6TVPcRO4
GmkNp8L1+K8tkOfmvF1CUvzG8M9G3jyD1pkX+6Tvaho1sZmqh/eMukqPedNg
Zu+x+XUftCxOeAfjFWIcKixX4gQ/qFUIjqpnbb2oP7vXEawS493Kmem4Lqn7
BE6+T1/XqxDZLFmdGjPG+JKqGnWuPZ8AV9fMM7dX7FFj8sQTda6wN6a1SFuf
rmnAx9FP1woavY0Dg34k2atPej/nDUZ6I1hvCXt+pwuOgVifvcDyOZw3U9+d
1RicTQEQh2XHL7openCZOBWv7qjLwMq4KXYt8ed/A7Gj/9EJ8qRKNIfLGnAd
YjUpcZPc4ar6ZaItcHGIMSc5D3uCNiW52ywySPS+kAMAGedVM8POWun4MO1W
7/iHnErAj/3Ojgmsym6taWeCEWRFjDce0q5gTExoMgbHmJe6DqrJr5J3uTiz
qylZU0uOaJzj4EXXlm82bHRTGZihQBt4KNx9A6cI7iwerTfoC83dI/4hfUaY
isHsWnrs4X6HpdgzmjOh7EPfWTC2boLQQSr/u//PfeMmpZRQjvSiN0jtNH/r
oO44LKqMU9X/nXgol+0QtSvpb+znmXTIht4wEORV/QRvKRkTOoLa71yhjXHM
38VWOFL32G8CdBTkQAVlyPbX1DVU6ru417i2GfPiEmf7gK6etqacoQcdeGAd
FnjUi5VaJ3I3YU+/Pr+zZBdIcmoLH6wXf7blaqOjDF7qEYoMU7aGVpFggWyD
AiZk4ZnLzL0cDACvgS41tn9yl7hXkgjelGLKm7XUg5rkduRFfC+g2f7OK4FE
YooOKAYZS7GO3+k+1CH9DUq8kD25PlSK/snyxqyN+snOxQxOjimdvN2yq2op
Jm3r8zAY7iq3qcT6njoUUrZay3Gqv8sZqnSZuQjhl0ffq1HM1uNFv+68evpQ
wLqRKXjgcfEQAbWyORJMrnT0R8jqbYGy4Zlju6z8FFjcAtpKELfRDxhTDzL8
5mVNQ3ckp27uKYJi7BmOmg6T6gbiX6kyVd/YtUwUsHwf2wsOl8cyhLg3Cwsr
6ZrCH5Jedbw2wqBKPxEuIQD6vtlohy94T7DFM2fHSydo9ZZMVvYkW5x5/nmv
b0o5S5wKQe0PD9AK/l5UnM1Qpm8MHpP7G57f6HaHGNoZKbvrAFuGq2Ttbg33
47mcmSuxZT6r0A4XEIozOJcdOTAcik6juGdByWDkEDDxvsNXBotCEtQ4NA8m
DzDdckuJVR+xXKw4TacE0vVm6Kid0fredU/cHsIgDGFFkgYGISqe6IJ9Qyrm
DKbolanE8gZSJ2RZHsswV47nP6+Y/q6rxre55/LS5MohiVpAVRx7zx2QzmCw
bI8CHEh3G2ykEJAxuZ4j09M3Z4FWhXgjJYnOTpgd1EVpz45jEXRAbIu3Ql+G
i3JtTokdKfueS/SOL756ALePM36Kq7HJn05vwce/PDiy3Gjn4ZHC4MPish8J
6gi/ys7niz2ZZ3ELyBeNBABAIXBOgCss/WSkRNVPryGpomnBEfEzO1+YUAk9
CMLr42pmwxjRUrKfzkOYX3XEvild8iY6RF/VjlQXVR4ZYynXK9bOx/pyBBoj
nOBIH58cQnrMtLCVDQ/2w5uSueNaIVL2cN807BkgQjhwfA6tC5JVQssaTKQs
6rwGcrrRLSGHSEkk1wa4g7tgKksL8P9tzx5KIt80rQ/oRkN5m7rvvYe8paW8
gr56ZiLaS64Ru7Ly+DsXh/34U/+qrvlj71qTc4A8fi8GlW0tG7jbxctReGpG
Cp6Q

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "t4xPJbmEH6v4SVL0gN6FMeKrn4IhP8uxgDEXixmWFrfkRmUmHah0woCI0NWn4jNi29PHRr8qC3E+56ObAVSYSIpu2luY1Ux8HxJTmEZp8dfWiQKOAKoquE/rRpOs7kTiASgRERfy/4yFwiIwBiIeSiYycsrshs/YcSPLGlUvkeFONkowA1F3QkwXAeAdMdMqD0IZHCYUiyRDun/uIWwwqKpaY0MedDAF1dXVq3jdOlmgqv41XH7qi1niJwNQojSRfAV/c0bLm/XAAqpF1IfAyYaXMSoZRDyjzF+YILciTg4Y6TaVLJxH62qYe+2qIQPhdIsEko1zL/QljXGFqB8Kj+dOiteXOvUHrOTrWxkQnzAvdAXFaWyM0d3AhMe/tVKiCbq1lDQwjacrmXgJ3Q3tSnQEk0rLrfU+cOlzuyUVI7RPmBBbmAsCA6Y7w4Ylj4RnQ7hcZcr+dHX98zZ/ln9P74p29aQfZD5rAxJIvFw6THdRgPWviuNj7WAlhlIZ7+2HT2zJ6UouYcN7K7Q1CgQw0FVwyVJC4i38KAFOGH919/gQvvxL8TMaZPMuLQWOcrN04NOicSrpw1RBudiNhNexQ7f2LCbVIQinL+rddUHBxzEAG4tV13BObxCFRrU/XpOI0RZ01vUaQDtrpLdhv+rjmssYdq1tK6SOFWP7HL6qT+w1MuQJqV4Hwvh3mInTpb2ih5InNP++CvkS3cvovTrtbd5SpssiodhypQk5Y7gUk5cN4xtp3VH07lFki5JU/K+CWVNDZGa+Nyk8plT79wJRoeN1Ti1eMme3e08uARrJuR5yQ1R8UiV3PRM4/+1B1ZlwjP4USvxQnXrIcrwmIM+X8sqvRYlKaORmFl0qzjKsE7dKjWoHKl2UucAFbJOnVD1cimOHu3WSfrLAwep946PovrQ3kqTKYW5+OT7uMIJ1KtdgS+aWJ31xo5GzUUVMtP8dZlmo6MCsfOu7qlR3TTXnusI5U4cIu3N3B6AGmc5UhuYwRWHKQuDPc31EXmZpP7VE"
`endif