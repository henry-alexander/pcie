module system_intel_srcss_gts_0 (
		output wire [0:0] o_pma_cu_clk  // o_pma_cu_clk.clk, PMA clock from PLL for proper calculation. For simulation only
	);
endmodule

