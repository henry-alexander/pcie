//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k3GfNTO2mInPCGEX1mjY4FcKPiEu9IU9emiTq08URiYuGp7j1LzScKAhSPvo
YnYOjcBJq8aqpRP+q3f4V47Dt/o3P7PKHa9Ah6nAoK8jNT6rirnI/BAfDWU3
hYXTtYww1FI8NUbWgrcG4gm8f/QFqv8ZAiUqhRn5mI8D72TIaTMxsihQMmp7
tEqISFUIWMI3RTttWM4DViKB0ufHU+NhATUlbK1pwzgEuq0sDRCcJklMWP/O
gj7sF9oXCdMrAN7mPWK8LZ1K51wnJz6uDdQSoz4yZIrcrBqtU4cJWfrE5e4c
VP6L9AYwLXcDEKpSqANhBiAAhxj86iSRnnmBf7W0zA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hxfwZpklrfjiX03cFeS3w2hcoFwvkcu5ESQ/tSY2Yux7/NbMp/CZoNOyqZK5
ZdXKXa+TkTkjYXedcUhjYEiRocuYE7vjDkr4tCVM4T2H0coS2XRirLj0MXSw
7fK7NsNxGoo0x1veSHKXaCyYph6BUJuy7zDu5vYIxFJ8zsF4GB/2mGw8jBIl
IrtJKUOVwO4G5l39NqxFrjBr6sRjNd3ogznbLNxk9+4bMMxVQwrWfvLbn8Ef
0oaOUcSfBygGKltb+kNaujalJu8enBf79ka/UDRkk/OE1FD/o5mBgFB6gFUf
t9movvUOMbbXUt95+HoHWXrB23RagrySB3pc8qDJMQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dvMHDWM/WydZO1gbvnunW1AAm3/zp6HzNu6baIOaLF0HF+EEeY4dvO6EYMF8
0ZkL+fe2sPtOyBWtmz/aW9M3kvWpOyVCPTNTXf4cz5zIa/uwPt6TGn4rM2PD
nZ7J3fqTZmy+eUitkXME/rEltQUD+xn98NGYHUYq5T6HwO38LgAkIuucTt2/
UtubTUry1CpX0kpHdMAwJezCrsIwxIp7AD4lLZPvwifRRdhjDTAo9Kw/ZLhN
xs8LxKA3Iqx79KHYcxtv8YuVihlAI4f5EFNVtmUNcOdwbWGjLio1NeupXBS/
IlGmI50XPYX8HvjS7NDrJn628OCqyi8D3150tgcC4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RRI1S7flOd3ILWrSVNphI6lCBSJaahNi//4fXnlN92fEBm+9GGllZ6YH2zsp
RQmI0XUNs2J5B+GST4hnCowE7e8af8+pRRbhzsd+Rj+jPaWo7z+70awStktI
iwdgiTTtJ6bNo1d6n9KvfOZZeHLKxnZIXzOeV3V8HewZ1/O5dZI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
RltVN/zIHkHiaxo7bTWFKeVXHdxlJHFLtW8d8aakAd4xH+Pax7eDGLZDDFUt
lnWEX2iYBVcjYXh2pURsCtvwJihKEy0ET+7v4/cFVnoMgD+tBmbpqNdkuXiW
2K0mIwRV+Sj5eIQG8RmJQ2ckhxWcnRSX+880cPU6hOmm1cFZqyB128621QkM
NSEMTW+5ESq4O5EgTveZK0nDBvREg0X0ejxrZDiqb+arEIyH4Nl7Vd07RzEo
JzSRC6x1CXnkNx9l0D8K09wt6Oh0Hh6Gb8SUCbHHzw5YMwYKnzEnFdfRUrLu
wA/IAzjDUt0fSSqWFTnFbOUMkFy2QWhWKXtOAuRJ868u3zgD/D56UfhZd/0d
sqc4AxkoMmnQv9QMpxjkjHThS0yWNA5zw9yDwlmYIZ3G1e5CPmy0bK9xEqMO
PbFSndTyba2JVuG1CBZfo1/GllNXc6HVvDeRw35dv1HLE7npiR8rAyxONPse
k/r6if8dZcOuwpwaR+XnZe+MdSY7Pffm


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
m4I9EYD6yTUu8bvCG6W2JnPn/wRKFfev8h9xNieE2roiW7KvarJR26MfCaPg
FHDee+gUQIuD8knjjTa2cdErAiX+euEYmjOp6VRKm2VjDjbDsnst8bcl1Ukt
UYqBpuN2JxGfyFF5o9EN7tGGC/tKGwL5TDM6QPSf55IRZCq4WYE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SiT7cCf9Dzz49kd2yttgGV9doN2VWBSubeCG7TzwWliryl5JGTrdpbs41Hhy
/dUjyw4lgS7QAJBnlWnz3VvITEj86EC67Iyx9Y7GWFyA3lRZstJ2Bz/8Nl6p
KARNsyT7z/ySk8sp28GUrr08+SFJ0abVLotMEbn95rupDxUBKeQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 44624)
`pragma protect data_block
rIR4AFlHraZOLqJ2b6hGekaa5+OwDLzrTDt+GmInbT4KotLaU7eiIV9eERsM
VdRueIXf2ShIpFSMY3n0pY406gJQEB34HZj4h9KeyqA3dcxALuaO1NLX3RAb
4w9aJlUhecASvmR0mmNW+PcwVWw89cWW7DKEWcfIrrtX5lQMMSuC719xYYd8
/kbFNe3AOqzutpl1AdYqsLvN1DCIHY3NDexJsaE72Cdaa1fSEM1dqCOvptKe
3aWgp+wFkkOGPOBaH/oBde8M/OPQlveMjOFCk8WbF09Eb3SRenzcRbkV/xBW
y/KB7ZS1Y3TyPh+4bUwFS+Do92Cs/7SvO7Kg1aP6qWFxi5YxNMh9oqOVakPx
i2Z8NlW1yAZMjPIYKeraDzuOCKNfVnK5pSE9w+uTEPtX/UifQE72uU5X9S98
hPnbZ2iJmX8M63Qqk6XEek136bv6MMZ5ZDbGm6eLJdg8Gkk9acT+eI5E+mv7
4+1mDstDzMNHXsVM5I99dBaUKSB0CTRkHvJ+0STmRIknQ7ArOg7vIHdSQ7KL
37UtZZ9FyQ+MpyxjSSoEjSU7XF/8PgErVBrzUaBzp+BumLll2XJ2xck1UrHH
Umozk4fDOHyUmB7fJv393gbQfa+2xmmVsOif7rRt6f93oNfqsCTAKlJELEYP
Kn521yq1HON4VF9nrugHKqucuZcPqI+qKy3ZXl4k/hGCBuoX6oAl52KuCvww
y2MQK9ZMsjHh9NIjQZ66K4gEakyvkndhfX6syojogn0Zdjne8dtmrca1y6Bv
IXD7jADWAVYTSZKSKChb4uiT3PcH65WpmcqDs72Gt/X/HpswCPHng5KZCNqB
cjl9m4ekTe9P65oiQXBHntKY7iM5mwcz2EAgN6IDUpqHjolNiELQ/9KaE3Tf
Rxi5O6GF6zRCX2lOb9fFMUzsnkWchZuNYYyGBaqP9Q13Eduw97fdywpvYffF
NsU0/+1DNtY53zZeB1qzM1QR9gJFxuq8O+QmlZVfb1YJR2ZbgVOw2sIY9jB3
z7ZrgQmoeIV9PgrB3UhHMMOb7/MjNThq4Ui2okq1Du9ZokSHP/OO78kDRK48
aF5M3OSKEl55vOmU1dYZZpmB7AVU188JjU9VHKFS29oXnfTtwwoUfBf5zGpe
bNfqeG1WIOUQ74j63erLKkhXogbBxqqU+xNFQK2YU7pLFbIxZnh7iuMxyjB0
vkvISsmFPQ64vccj+6hYrAGUkHRolDWhTwuA/elZhVK4zbPwyi6FMntXl8Qt
RcFQMiB1LAgf5EUdse85gBqLJCpEz489CN2PXPOsccklNcXxJ6gwVlJWY21p
Ayl9cG/I9cWN6RuWagvu7Xly2dXLmDzCPWwk6EHpLhqBR+VzVSIQK9nqYb6t
BMpqLO/cKLDybIUeqdlKZP5yG5sTzd6nA1mmei8uYy8eHXL4e83j3mCeJY6Q
qXH2eNZ6cpSLFgt7H3Y6WGVc3jksuwDs64JX/VWv129YDweuEGhLCOPuoCTW
F1Qqx++cV5LTOo+m3qyEOHJC6gQVeVhxatle9uyslfb1PG4rPmFq3qnBdsks
lVJKp6i3GlTK7mZySxKaqmL6p1h1z8DUSkaBbsLapuLyjLuiCKfJwDOylwgc
Rs/t+7n1RScXTW9WbeGB/aLJoly/ZSWjbBteyZGxSXgm5tbZ8xLaS0zpmwgy
YKgvCC6LvVXrEClwhBYSk/YAVeWsUhykvg0SNVzDv2hB/YS9ThLq8u777Nhi
LHfuyQJX5TPbPtABtQaMo6YkffagSUBDMi+vLio4uY2RFL/zrs5yQBMRiNvS
r2bgLrgBL2XQdZLRHPINaecE8kKGhQ+s9HAN7YYvJQ1BARtkaKQ6HpntEDe2
CViaNzS+MPFvao2jVE2Ngp1BMhB7aM7HMbtCcmO6XQsJ2WZVM9azrhZ42VBi
Y7OJ0sxHiNsOyc367w4LMyXQPS9MWEZqjuLNHv8P4NsKUsD0VYCcxRgEo0h7
P/pYgoEfxfdmR+q23JDlt5D/BLrxJ7TJJShUMZLr9c2+QkQVfBOmLivU0YyE
6dU1lJoDlpVqwbFv41reQ501+USnBT1IpEPz59i8hApXA20vAbubERWiVGqa
HRHwTfZil4zMrreHB+uS09b4gWhW1MZZw94NP/nUD0DeNplIJ6kPTM850t21
tma9Awj7ndD36GMuAgMxpAZq6lUrEraYYA0jVG6IS9Lx8r5T3uwKmhcQI3OZ
+04/LcgZDQP1C5AWzn0kftkmooziVWNZOY5QZQ4uWIe/YbdWdoSBGy3joXIN
X/4sSo3ffozJdx6dBvQ09eDiZTs9o5+I2guVXx4ICbb11FT57cbIXeewCKBi
nMKf/DEOk5f+dW9HutDgerUStC9POidTvHmGBvCo+MVSkqYpT562k/BiWpGp
etzZKTu0nC3auaIw/apVr1A2E0cBFg1H5kBUpcCk/YsGFbADAuvFaDFatIt7
CiyWhIsqAIMhxr3O3djKg0nfng1lhagzObNgRU5xnk3yZwoNu74HNPKSOKcB
HiLXUPowj2TXMOzZ9LlgA1xUhhWEIKy5Y26hYlDvkj/IZPrUXCeWckaINZE0
lS2elrZglzDRG4XenF57nz3kFrYDtv1dpnTIJMwKCYaIDLBdriEOnW5SwGzJ
qs1eflp9Ahastkaqy+SKoRte19DsvUnBjbeLNOIRUsl/1O5Xf2ArQBmSsdyq
CWOj0RL/MH77n1c18RjAoGDFO5SD+0sQspjDtuNLjvir9nHtjhe3puAcQczz
jAD7fHrefqXUb1cCA6WjM1wR5/DVj+TwN0zytogcQDxwHW/T9op9554ZiQz0
pDtKe7dXo+xBplGIHsxM38jfQbqx1k7MqKzHM0lziPZF27MbbvymKSxXN7T6
ag6wki9Q7BlpBTEaXskA7yYYDRlpBNTYEsM6Pa0mz4fQTOBOF0N1L+hO5ZcG
/JtL7fA8aIDWivsP3PlBx/RFJ49yudK5gAfUCQPwg8s4lT5LfHjOEbl/nBCF
bwhOZl7nJrt35Y6jvYripW9+kYCGvFucKMcLy+A2cEMHqaKhfDlrJRbfHS2k
MdlkWHeDmU6PFtuYIv2ua2Wf8AnW1A+iUkR66vSqZnHP37gbgLmynvqvGZIv
RPzunh/X0iBmDBph9IP7wnUtBE/0bQemdPx0U3caUM6CUc+9SosnuJUmv1lc
LoLvmzd2L0fHuYUeWbkiPQZGve8HbCb3y6IevzkRic3KbHhthj6bN86Xxbmw
wGaVCS2XHWGQMcjxtNH2eHHUx/AIhqZwaikXmyjCjLUfYahffzhtvu4Z34YP
4ilW0KwAYcvvOVrH2NTtppIgIzV3N0HIW30XF3TS70wiApime1H1GoDxr0Al
cfKr/8O4JhwAg01guh6UAfzN/7HPTwvRvDxSRmgd4/+R24ZRpc3mnhWlqTIl
naPTCE3WwTpCfSSWSF44XybM2O+5qCLNfFWH+iIjh/l7DnPwYjjessWh9T8h
IsQJJJtyfVcDTfHV8Ll+dDy8mRzQimkrazdajHo1SqLv0SqCFbQFNFX4GXse
BdP7u+/wMn6qM9caeKSVvLGhskMbqkKdOLtkq9EGn2X77TPWmXvfQqxJrwcu
g2RITwDWlZaYg9aY6R67TuZOzBU7BimOcWl3ugnj4PWnz6+6FZfiowpYI4QF
PW5NOe3Cf2q9vBh4fP/Tbm8R4gNUvNgLNyPrHUM6CH4IbPT6+4FIDPk65k2z
bSUOcIAGPYWEEpF5C8JiLXfXcl04K+hSzFSexaX6QVVq76766+PA3oYQ+ydg
3+MvJvpcIGJ6OaEtVVWTsfShgEEH3MA3fQQ8gOTedYhigkzF+F0EmAp5MwG0
r8Xr9KdN+0o92Y7WTdRXkQonxvH260ihEJHmG1PYHb/e6xNuos4YK5pO9CyR
mnWD6PKOoU6raPbmRRP+Hwkqoe23rC2CN6ErM/6LuDBHnil9fRrWz76mnJJc
DyOx6eojK4pOvwyz6EG9G67a7tR/Fu9m18FRiaE4nHQXm4jH+a8b6y8Y/dwX
hbPAWR77D/xgr3vimi3ZPpPTgtY9aDuKfzZzdHrrwqdHUabei4HmrwtDq7IN
GTc1aCsZ5MjZDArTgeqP7uC6eqBfqJ/mtNguCqLlbv1D9bzp58nZT2AeWYKS
qG8QAhQVC0ctM6c/1eneqvm/thmkbNIAOUTbZw6JbaqQ91iZ1NrXuGPc2BlR
zksszr7IBj88aV3nrme8kuzUSs+KZOuMOEPEuHcAmR8z4/+PKat9m3IYkBU7
LPdKo85xZrzDS+hF83xoeb7F7GU9PL1w9w0CSc8yhBkQEo1y94DZ7Xnj1Tv3
Sy4nkT+sv0KomwBYGqqtKlZRJiTkvLJABkBGYsBMJtfuLZ8sTcUaRA4abXE9
FTMB7sMb4Ay9e6ENoPeAtYIzoL8M1N87Pzo18kVI3hzjvNUQPphhE7gaFBr7
FX2f/cZAXyGPVY09FTkoPxetTIm+AF5CBHsKWWTGvdZymmKACbPqYhAioL77
N5KOEIhao24VCj/o10boqSED/qnaLamAh97nDhz6AeNAPHldvvTROC7ouFJG
KxDiXwt22T7l6PnFVoX3BycieLBMH/gHswwjtWDWL6GLMJ5ZwjssysK4hssP
S3fBR/EuH0CDhjnGwC7/gyMUAfGe40ewlflWlY4OEgky4IFkEcMU8SPpXnMj
W0uK4Ud63cE+LbotmxQK8hUTvMhDK6IOVQWwTa/Havdgwur/Kvy4mytuklkf
JG8haENiQa+GMg89VYfVG/vjadWW2vWKQeX2aqpf8jTz+hMQSuefmtcZ/kBB
ulMdZ8BN4vSMu5XgCBDhoGaSr6QziX6eAtAmutGWfApbLBKrkuRpWRnGZuO8
+s/FsUguL/jqnykvlZNgVCkFrXlT5E6jaTBKKkFHK/bxOuEz130iIxGM0Boh
wI7nXRG1KdtC4p6pBDlPPQaQOwE73NIbkru1miJXjzeyi9gqgb+4C31AJvHj
B8OQUVshwM38CJ4i0s8Vzdiy2TMZ5wpykJBjS60pgBj+3kUQsvz01yfhAKGQ
i4/5aVhrfcWN1uIYI1xiXv6o9U/2ypqmylXqCudAVcxOkgHgumzXUfUGned5
QQzT/SpjnR2+wSthA5vmALtzyGoYtiKXHy8J/y49pcKGni1DHLDIYLPW2/Sq
GUXLIUtZB3/fyPN7H0mQ+xArbjffyYytXb4/mny7U0CMxFzd1sQKlvYlwvTK
ghHb38LVsBgXr8zBC77QJWMfe1eSEI2vIb+yr6RRDEWbaO0+uoqQsaMS8J03
x5UXMkzkT1noT67syO9KBE5lkDC5cE6JgJiDk+fnqaozaFx/Drs2SUGHB+4y
TJCwuFHJ7+35YVghMhE1nG2UJj8+derXojGksXVHMXt4hStHIID4hNOYdSq4
lvnZBD4TC2Ec4CrOJtrPPCDZMydycqZhdIRKVhVUoxajukXJHfL8YALGa+r3
qTWE+3selKkMP4iyLu3rfT4pRhQ83R4oabi0y8wmrSafkcJCrU39K8GfTo2X
bfg73qhLejyR+pZTx3CajBWOcZRBZJGAjFxhCatxTRWuS1NfRVlSPNjIYdfE
lm0PaVjlHSoZlioxvBf+/J3xBr0Jsbe86cZI7WQFNOnZZBqciKZdfpYklHni
2RVE3utimjUs17D2V6QBSYV2IotcHNOmtsfsTvzMqTFFwmWWC+KYGT4VBKuh
c63k64BWRMMJw9V1pUH34G1UI9eEleh+OPTGh366mLr8dw4c03pLUQsJJizA
UKF3tMmAjIB+szFa/+drdiCs7V2CKHMGFqgWCt20ILYcua5D1ss0BrnScInd
LhjS9LviQpToIkqUq9odHiz2tCSGlrDjqqnwNLXlJiXZCrYzq5vZckA45LbD
/z5UpTXCtt2nWvVU4LOWWrpkrL60tHxpvUY6kVaZJvdn0rHQXO/ZmbBlwKoY
fr5noWWGEyeNmTseaycvKvIB8fbuTmw0JEqNjfozzdr+pC48loSbcLXQciZc
QcXq2u1Kabe8/+O/QTJ6nuP+nVom2q2NHq0V1ssVXfJJRGQU0zlk0QtSsaJH
wZYr7gFU246wHrmfQ5TIWjg297nf22ivrbQr4L0/f99kDcfCTQyYh7X4depJ
h0oXNu7+EqGVI7RfxpF5NXy04XqLBiGVi1akhWgOop8LS0Pa8dK1LEAF9Een
FHVhgkNKCkjR4SQUjj29MQvYlfSIr90//3yz/nyw7+k9JduaR0SeoU2FwJeq
DPZAJkqR7epHsustoUiF5AvQ0azelmuWuXkvCPY4v7kjwC/KdTmbRFEFGsdp
dypxRmQX7Y5m/bYDG6+A/nxb24DpkG7fMOS1naSx8AedZI5fpkSo/8aAOXXI
HMxlAJBx6DiBpFr56oMaLE2kENmkwlWv1gKmE2L5UQpX0BTfPmhhgOjE/bYg
ygNoYKezgZavuCJsxMUFT5Ha0KWE4ysyQTptafjlnulGY0qM8tpZ0BJ9W+x4
5OImVTIFQLbhjcM0cSRbkFt3PvGrcxeUWZvxfc/9qIN6vFCXaEouvHUHcSfz
CqtAHIF+kLgnYX4kP+1peXo0JYx72LuhteDmT83nUn15zPZLJLdhn2m3X5O7
FB7nqnixyMhR22Jmay3uC7uSBix9WKzK0tsw68aW7lgGvebsN3RV2jSt/ckG
NMVTy9E42XVOAXfTYiiut9UYlQSd8PHoOARyn2REXE8mgdYIuetNHnkoLt4u
KDBSZ1u5L2tl47UGLFi1awrI5anAy1vQ2+dVrx750jxjykHkFQbqJrPgcZgL
IcgeOXLspgKOG7plAzGRiWdiYZCriquAgnNGq6YujD0Z72vcoa+7NF2BCVzP
xwo5JEDziyUkTxx9hvtukCEsHgG/OTYwBmGxTkGqLl7Iml9q9DddoDdKggu7
zX9OncfsNQqTF6JqjzNBcw88S7WmI3boncCJsy60tT/26nVnaWgfZhtaC9uD
17tTzDrSbwwGlcyf1UMA771/C/ZkwauspZ13rgEEVMDVAil4Ru6wuty5i/FW
xQvZeKfZ5UyTKH0nQQBHYqoWlQOZa12kri/6D2224gAocdhuEarENZyvoZLa
NtBiZtIMcWBbNkLLacTFwqfoh4KSMjI3Juj4jl8N+u/4zcQgtZ2WRLqV7h8q
mEk9J8W2lRaEvari9Pj7ZuL70+vLP4MFnsMDYwC0Kg5VqkmKsG+zvJskKoFB
GCFjeLUYa19f0jj8ILlR5uJZit4/NzZ0a6W0cQgoLkdF9O00UZrLGPJROYU0
MBKp8LC5mkSxO5kAkf0xRexHIAPI3sjfDu6UPtAAx3OJ2jed2csxcTBppWIt
d01LKk8HSMCHCMpc/OJlJrfyXgVDVntzgPWkVQet6frbabdcXX9slO1MXk/7
LRljNcgoux0yhbLGTfmjOqHEqWNkiV8SJiKwi+JAT3JKKVurEegB93O3r3PR
my507WA2p8DKByVdHaIPJG8A2j20eRukHKmS4/Y4vBEWV2C31RteJSeVXfER
thst8TH8W1PSgMxZYuqeOKhZuOwYFX1tegkfH+yTz48zm7YX56l2WWLLPCpq
qHAmlSRxrGh1ikDd8YDmmJRL+a7kk3bjFLVTyOZfyGereQYELeh3sjYtn0WM
i4wB9lzfTVY+stmYr6iA0wWiijHchcC0kfaN1iwV+YDQNB43DLEbGFSh4Ren
vXRpmdj+wcsqJ1BoFCxfIIg7+1XQpTkeTr6Wdc1LjHApcvL0Eja4nroG7g/X
8avprjw6EjHaRdwqPu/XzPCQIhR2Y1su2+YiouByTROTWY3xiK4GDO+OVgOl
RntetwOFUJLjG2glsfg/oHE49Q2n8JVK6P6G+h+gJxLzRQUIUhBgCpBk0lp6
39hUtqGSY+UI4aBY4AedMr1XHXVu9acSMXYHjwZIpTS8JiJlNs0UbhoW5QR1
BZlx1K6+QergR7ZELZqTvzLYGJZ5labhc9/kfes1y+f3RMjX8v1Yx3Di8Kzt
YnK5z/0495lsMz3jHSoL9izkxXxv2ORD1OK/SDDo+llWYrDa+FVyuzPw56ur
Y+8tcvXwVEEJotjNii1UWVclPEjFMSetJE+5alnQQEUGY2jL7mpFFQ/tInw/
VOXmIsVBRmPpiLNH1FJvv6nJ57UlD9W/PlU4ImTsXKJi7s8HO96CA67Ivo+l
3EkU5MH/HuHf4Yuv3nG1gGbtjVM/aavHTXdIH5kfeaC0/k7VMWuYRndff9fY
4MD5LevPHGgDLVdl2/n/+mvuiV4ueRvmhP/KEfi/mI6pzKJisD7esWJ9+rmw
Lz/a0lNdi41JcKsweyH5mkcy0hl0as3KuwFWfeAw3V7Ezw67qld++khXYcM0
44YoqNiaoXPd8aY4z+PrRRwq9shrEv9A4ByrBXUe2ruOSWw5huoR5nZFIT9j
iJxpXltSC5HTC83dTS2ndAl0LdY+8gHLdiktukvy0/BA946UdcaYKDPt2lGy
fXkjaOEunZ14Os3yU23aDu2/iGdHUsNW5wjzv5cCalGfB9t8YE3lLSbG3Gqr
8bjd/lNS5r43EM1O4S0U8xM80uktg9CVesndZ/viTq3+IoI7Ug9WKyb7pfUA
I7iwrhVatITvkizjZ2faNoW8NpD/B58SXIJIfx7rZfwxTaiEs1SaOteq5KRW
NIt8iT4JOnj3qVzR2PJYIKAOT27oMORvMY3cfthDuMdjBAN+q9JwHOQBEmVY
StpDYEg80YV6HNdS7rPW1NMl+AdQhpv3fVvAPsYr9HdcVq+bApbO3wgCkqhw
/ZnSNfF9dw9/deQNHkHaHZdsX7fJPnXcqxhQjJ8ifTwMh4gkkrmUdYrjNPPZ
MTHDPbxPxt6YOkdjTOKX0sHjEpvJU0fk6ZYFhehR/F8gtKlY5u6eb/Nsn9YX
+j409QsB9ze0wmg7GKLHd4O9ZQf6w5DtfqbMKQAhJMUynap5wplteKXl1hNx
6tT8ElZXv6aRfMSOaR8Mt7aVUMpQ+NPFwuf2NEb7kU/s3r13oVXboWuYPcP3
HHsO9EDkKYerDU+GfMPOiUeebxMGXWbpCLjupStVC7QuN/bL8z0Ke08AGy3x
FayioN+q/CEidMxFPOulrXvOWuaIE/wmnMBlSc/tBWCIfZXIDT2nPrDmwMRs
1ghFGlkE11YfiRiZKNxm3cHMoPH4QhgvlWTO6LubeK/YmKEcdozJ6F6ZL7Yo
oKkivzkYBHVHD0dImAFpaURA/ouJRCjJTTmsAbUTcVTxSrgNbSFr7XZAnQRe
Ny8azrBQn2X4u7RfL6I82sPNc0Py531CpzgOBEFCGvcJ/m+9XzW9gd3mrClc
hiCQdVdFFaNPObL3dHmJFJptP9jcIIKnbI+eE8o353/JkOvcVkuzTQXjCgQJ
Bmt7cs2mIu6EsA9HBtSpIydvB6Jm/Sfnxw9tTdIf3RN+lbPA9CqVZCkdflXP
h7bA0hkf8Y9X4W9lHZX/xO4ug73XMmWWJ6CgHp9yRb+DuvUokjmYfG9ZJHyn
9Yq/yXMDvoKO/rXNtSzyyjZ6LgA+YiEYojhhqjqONOt9EzS4U4LBUfcS/Ivo
KpfCtm0+b6dk4mKc/k0FBQdd5chpimTszey3qdeimXJ5ApaN6tjGBbJ4Go9O
PC1hgWW8M5U+J6r4VMy7O5wXPGH7a8dzHU4kINc9t8fLHXojEl55Ssyv0nDc
gykwtz6bjXlnJ+ov7XyROdowJ2PWe5QpH5yEmqMoNqUh/X/cjp/baSeZ8Qae
eepwFJCUKQ89oj+ou4Uv42CV/7Q27yp9Lh1/ZNdztcgdAtZPh5rapYwgrIFX
6WLusSrVV3VqJ7Q43gl52NAR80JxzbTCBvdEsWchdpNQ2zpKjQjDppp/vA/O
hFmEDp69DUEcZpX+/043b9SH/uov23oH2Wdjpo7HBEXq5lFAVI8qJHgnahER
bg528SGKX/5rsb1IHNJOH1nXXtqv1AemElJYvCK9tOGMN/KhTinhdOpqRAJv
5RaYm7t2kA7pBrt9f1BnVaQhYEjK6kshBy8IQiFs+KVU7Z8shSiTocWk76/7
QdHKdoFZXd1bqF4MiUFY0afipRaJC1k9h+A2yK4qwPjTnKv1xHgfXKfxPuVf
t9rJNXNFsIPulWcA7fKefh+aALOTz4tgcUXDMa4weZTmJ1Syaw/gdVZnhE/M
fsI2FOz72rtuFNcCBl3cSt8qY38wY/zF5acCrL5ABvK4YzAcNirwhEKlJX/w
vyV9prXSy5UrQOOg0uT9Oh1tdE8mt+tMCHzchZZfbt0fuz7p5IZ2gaGF6x8Y
igL3aTsNFo91U0g0TeViQLy+qKAe5z6RgQA4QTpPmiS/3NVeNOC+U3YglCHL
OuFgQ718OGJIlxkRcSfmZlwNvG0ABNDuuw67NCzsjbU+lEaqCDFxJpQpv+uC
eyBrQlnjmgxdf4sbdtJiiQ0W6clU7J5/7DesqMvl7KuXVGCe0BO7GjIa6yJ6
/MC2IjKpjEecTWzXXbYyTKfLR7RlKMyYUB1Pu2ziq96w07AQ0VHaYocNCInP
MiY7k5mHFKdi2Weh3muoQL8TFrVimNhDf0sGCS+pNrhKvd6erYoucfICxaj5
RWHyHmAnefadXf8XwoAXXE8IlrllpDQGSWcEdI0x5V3gfrOyPLfXojqUZ86H
vO/JYcoSFtGrmEPcpDOO6NlQGDRXBagAi45q4VugNwTSju3A4XilsBR8kaqy
G7X5CszLpbqBW98Q2jcgQZytHhbImCxh2Cm80gL21FUwHo172gRF0392hjEo
/SGviU6PI/plzB65mbi5d7gqz3KKNnB6mBM7KbJu4QI59hRPxE/8LO80eaUq
kod92pEVewH2cWhDLB2ZObiyI9PErj+kfo8wATlpQDlC+DKwO5ToryXksYuB
giVdXA1IDiYLHXc0ouEdna/zHgzbh3S16/w5uzPDadopSlVtihJxlf5VLry0
Phn6eDu8EtQbpzPQ1DIGyxgmndZudD3cuKxNsKjGWO8/df7cEfH8mUqB9KyQ
4NGqIJNqfpSLBInFs2zvtVS2yswEdEbnjEAqVMGkgy0UdBSntp9snSuJImzr
8zmC3UwGMiFSGiQ1X+erHpSuq89elQxJqba5J+T7gBC0WzTe88mVxEIULClm
06gxRVpx0MGRH/X3sVWFX5qmU/KtqqZ6BrVJhevKHih2+MEkRTmolbT8gnB+
Yi1nmMuxZF9XK7KtidVeq25SmTqt/KcUiX5DavYTGm3qxCA/jpeAFmLYfHDE
4K5GYuGD6f4pXJdGxxlXKn+vW6Sfmc6eDi0T5C0nhtcNycFmLiG3T37/FFOW
JwbNYj+RPaxirw2SxqubBf/VAi/FSGxaHDzOV8Lh/RIIWOtPTjB5NogJLR0B
L61yKag2dIWtc2WRN/EXjJiE7Dp/n3BDP1HohJLoGHieCgS3wMh1msWVRGIP
wV6ggE//JJ46L+yqVpW2+onGAKPXzk0G9Iok7ioJP2/D0HR9/nqZUsrxf9p3
96/ayF3VPADRDptKSCeWrmUQ2qZeNjt9jeGBYFCRGo6gA+xb5jsjtblQpmc2
dgINSXPguS4JFMqaDsSiHGGbuq5r0DPM62AsxXS0FL/wdgE/2/5XVZoQJa3V
uscBAUf/NpNReSFKB3MLJzGoPE9dHHPDonnDhxicvVvrZx8iSl456G/8aqKf
ammY8EglC/oJvdMsk9T9d3jHOrMnwqhSK1kdRIbkNLxPuGmzALanWu7DWHiB
mo4JUb9drWxP44J0ceNIT5fRCbUuQP0LV0McojxmV8hCRoisfE7Uhr5pUnCQ
pbW/FPIjayAxfeLdUxlMQV5q7rsluudfv3n6dt9rIwiVmoIEcTrAYH33AX8N
rOjeQVJQ6N4is7Qhz+Bib0RPGZHPnZFWE10LcMU89/oismiT5bdMQt054VZw
T8m48LYOt4eGZTv9kUGbkto6H1UxTphJe+qg2zwlnSi70we0N+sF9qZCG50C
UqiMwiixUzLrAi6xT5J9SF3x9Cv6zUKG/c3LhwJs6LYOXfBDn0lNuw7QY9B8
BMwfdGcP7dBpLPMOGmdA1W5S2RILC/AXlOYm4u802sDLhSM/yjoE5fuOsee9
/aLUQOuXMsFfA5A4IxqFOQMPzRSZbn/IkNvHsWzNQk/psZ09+kSOSXVSzA8+
VJOTb7nH5FwY/+ssmO/rHjfo/QT2vWhZzzKLaEdn27UyUH31fzxxQOuNMeha
1jq8hyTB+wppKCuKWmz4tJsZArEZtRaPNIItZ9mYAi8i3sue7yw97FOuHzRr
EfOo9V8FGeh/yA4Rif5Z/OOkImHDL3NmLf7JJkTpwdqFDRwkhpr9G4qsBgXM
AzelrOjNW5emn5QD+JRgrlhghLMFQbDiV54GNONI7aMxzVNY/Da9vuaTvshQ
jiGPzP+9uB0X8WGYlCKAh62hK5cOmHS+BdrGn1+w8iebtPe7rFujIS43cNWR
gF6HTgqdPU+D4ZiIw4lNP+SoDoWPaL2WLZ4z2BKraxKQZGnCGr9Vvzp98mQM
rjqgCS7t7Z2cpnquX4YRGbOL/z8y9rjA/WI1dAXAknKL+EyRuOq5S9WbQ3A7
JkaIkExWN5deU98i6ehNGeZ6avljawuZuvnBaof5zE8z4YUYYPSwpXmpwyMg
/8TSA6rHsgBtzHeHMWteTs0h9xvDpCweYMXkNB9tCfSD2XE8XK/3JO5ZVXZq
JZTxOm1jukhwj+d13sizi6NV+2pra+32yVNBGVls9fFkG999dnjubzpPpS7A
uU57Tt4uwIrNLXzjd3Mc3n7slNOQXx7+NNKmEAEpZJY/vGeKUyfkDpbWlo6B
csG5ROURPYzki1S6KtbibLafW5RPLqqfBOeRwCcbqWqDkEQeS+R4WM+j9WT9
KkR4kPbzF/xpWp0J/z8XsEjDZlEqbwkxq5FPOTSgrfEFB4f3dQWM8l1gHmLC
/J2pj/4ASFg0Q5Ti0Dr+c7Xub/xiLcNMb+nlIJWOSe56bFUHZg8RFhDP/nw8
vVe55P31vdo8jzvDbBpbNCDfBuK6oyqSE5WIMj4D7/U79qsWoRKS/uE/ZBa7
QGW8QKLHJLjcsM6UlHftC47Qd/UKFusekUTM9XLlmY2d//rZ3LFL89WjV+eI
k5J1NxgkxC7fYF5JabYWR5QPr+hlKJBrfAX1jDynVyUBc8u225ikGkNhlyzF
RsGhmLrkjxjRQAcRG2bkHqkGhKGsxB3CPYhseDXp8JyqIaQoQjBcSLO3Hzja
iLQMWPAd643ateL/x8ItCPzfsHslWJqrarD3zwI+zWTtgs2h9/N7VHxu1/vF
pHOR7W4eNog7cUGvQUe4ysDEH/ZGsxA0tZ3sTtR3+68Utjo/KUB07Sl85uyR
2IbjfnAR5G6tEece9nBC3skL1nmpRfYQeSP5w5qT8/KKZi6gIQgyn1OVQT+3
svxJtVwl/p3szB2n2VsWDZp0wukKvxHtEShlkuCpqr5qjzz3vzEWJ+F1RoZZ
DaFCKq/q0WFQ0ceKaC/pRbjBfHfEKheyHGymf1c8UT+6hTBLkdcdCfjpgSRz
EUvfTRiFYsMnF0tdBHOB5rouhYZqBDJzv3hQvVmHcvwcmqxTwGoye00+nU5w
67Dg4jZxJsUbmwR6xFoniUmx6nRIhSdXQ/21+QP3J9mwly3wQbL8Z9ISHUUE
iBAU5v1GLYdu5iQiCmeBztuCfP8sbAKc+NaBGf8OhwcnxONm82DFXwe4WW6W
ueUAxaNakO0oxBEQ2EQsXFK4/1lb4IiNCzaxV2Og28LS7Y96QYQ1/OLkwl3Z
Fiin1gB7dUfC1SavMktppdMdEyVZ2VrmTvWeOKWKAq4dvB5LTK0KUYaM/el4
DJ7A8yBIpG5JAZ5NED0HC/wsil6joAGEr8sZHC5LJVrEUKlfrm4vUWrL+r4q
UopmJvd0kYirws+lx7OyD1V88CaOiHUIat8lfrM3ZCQaFHUJP3U7c0fJI6G0
FVi1igxaifYN45E4rAuSwGeP0yrl7KpMqaF1Q7BDoLoF+NJzeA6ii5jsgbRN
EBnEa8CvbXnrW9Nem6LZxjN0OTkTf4lBS0JbgFHv47v2W7C19T4xVpkFPoQY
NUn1dq/y1Nqp1lJM2iY1g+STWImzIf7Q9Eg1uMsNNE4S0ht8y29QgUlInyQk
79KNjBjgimFYetGzHvsx7I2wubk39Dbw67aZu9yTZY68wMwXGQdIJawOSXCA
STZnfYw3WhIBv5T54eTLiLYVPyUO0FpvY444DqNFruQl1xzVGoQyST9+DeXm
vhMVh4j+pJsgvs7eIFFqQcRGG1N6BlIgGGMQaUYX2IPFsEQhFgrKQSBFwJwy
4yZkpTiqhe4rPPJebjYI2dLi4cupQXP6O5YZl/w+h7lpZNRgxGPWaKAIlyYJ
TT6PdGQvq6Gji/lVKZ613f3pcdj93Ogf5BVnUcTn8sl5udNWBMBov9K/h0Dk
kVDIRQfkD13PbzmtUeOnx19xof8XqjJPBVDZw+0R7Q7jpU2SOVR+E7JJhbl1
GZS5ackvobSp5V60szEMJyJ5tV9v693orECrw5t4WBF/j9/eVlqxjaqWXM+2
IRjsz3ixfwUpPlttqZhOUJjEt+PBfZvI1+upAckWNfj33pKVNyFRdjXt8551
uc417VRGm8c8f178/7S+/spmazNMregoRm/OIpoitLXXXP1NAts84n48mPUb
3RPzFD809Sd8ExRf10dOOYmlgfruf+h6YoeBrBHK/5GCQjVP/zEajKeKpYQi
mcAUCkJ2+LScIr/hCJEQXLq1swJX/Wj0dNcAGLWE3JbKh7tWtP5gF2v2Y1UL
2LAhoPfgFtV/xOawHbnywbpwznxXnFjIphp8LoodrkG/dwEsJdjAS3LQoCLr
UtdJBqnQG0XCA54MNpOt3BEMdB/t4rRZ9RlNqmxC/13m+4sBLbY11Yhwu9hX
mKDvFFKQ45Xx72RVaL7XlYjYS4uBzpVoLXAkHSqfHN0WRvF5d/bVZlbWceWo
HvMIhHLrFNai7MCO1SnEXMU1ns+KOApkBlFdVZla3VAlUNSEnHCg5r/k7/e7
R/4VPoA4uAG2PKD8t2wbFLLk5Oj+GurDJ8TCaKw5UxbcdM77de2Vj0UlQV+H
yDMVUv42AxU1vO0gYHoisaVD2voVBwMuITpixgNKa48ytKwKTlgp7YLU0mtB
Y6gJn2CKc9oet2vMqXmTRdvFzNouQpldALo0DRLlSNgwOXcFiHgyq8HRmuty
9Ti5f2jvuqyYbYKHbrkShziaGZF2ZB01wcHPOQmLp8zlisBj3ScHU75CbMy6
6S0pfF/Sdrivkyvl0W0JGdf9STGK8+YYaS9pwLJBZwYoeIjDzt7k57ALQP7L
vj5lkxZ4Wtn1W8yiJEzlrrfEkZs+hRzVcNCLKR2IsZL1L7IOPvFvhVi1NxWK
xW/457DI+TbyqI2w/ECXnoXZUEGl0cjWJt984hbhjVHS48U77CoHdSlecofE
Yx7CbOimGmQsGWXD4mOTZTyOtp7lJp9i2usAqtXI35ljNFt9Q4ogZ37fE9iO
eZdR6vC+Hl2dgBCn7pIi0gUbZLuSUE8sGhK5LTNcetFHl2MUo6x62GWHg6vu
xqROGg1/z1GjF4F4VwGGMTT0MZXAZTNmN53Jz19kDTYSH2qVmhtuTQlvHf7W
l1vaP6iEQ3hLVwUDLHLLR6uM75EMheEElZy40wbQcHRk+I33O4feJ4x9bqRC
ceQL10GqpCTYjX+Gkl9facx1BJslH7FMvujE4F1/Yp1JppwqKxfUQTOviBEu
B5AlfvTGqnxKyFbP57I69z/to1IGMYtUTZMpQkIZYfGiXqfAVCl9qSrgVzKg
e6LEzXTH+8ChMQNG+8Je8zK5b804v0capFHI5mAmmY4ia3NjTC6S0GeT77N7
THneUEpmC0dUtj3rmmza4GnUtV6yWHpNl5C78YplQjSZIPnxR8Tmj15dJSKz
jHJIC8c1surNwkwjuBg1JV6Xq+1NBEDFNr/it3uaKTfYv/TxMXX2E2VOOS0j
AG0b19wm60pf2GAoIxqi0jdL8qOF3pIia6xFzqrcfrvpD1sjBxUYVO4QAjKP
AG416zdANATp9omfJfCui0nDRICTr1oCQHweQYrSi/QQY5ufvrCmtLNK4/a6
P5q5PxfDKConuK60PVdHV9wdu0zmz/PgGvJP5UFScWgVcNcco/NKhriEEO79
r6yNs9n0RPfbse32iQAtcUAuK2L9P0YEk9zu9gMjAwiHzgnvigO2UoyL2EHZ
KypI6tCR5C9o35c3MrgnCx0eY9sad//Ip8djsdgwhmv/Aps9oXXXmRljYF80
M496VVWZXuo5TjHMcscWnv5xGvP/vi9inCPEslPq11+h2ZceCEmzSJh4ZPoJ
GvWKWlWHwhGifJI809ByhIbqyfkz1ndzRqaM26i2NF0u4mJjarr5PqDPdmiW
c8E8cp/tBfnlbEnpGwhVLuenDjOIQknA4ZuVviHeQK7ryLFcxEK4n79S4tJb
q3B8l0i702SGzyu88I16Lw4UV0i9VtfGZ0ojTdAYWbZjN3vdI0hLbc4WlI4P
mStTst+KywDjUIUKNinEuuwwKi+Iegl55H34I7yNr7mHSvzmrB+BT9O3ZDi6
1zI43zFlh+7phmA/2UCwbm9hTBVCSSZdnV2X7J/bTg3bdQU0x+9F5MKt4G3H
lxhkfOoMZz3VgNSguhvHW1J2+njVg5hI5WDq5sk8DW4ggQ858Z6R2wCh8ILL
DfzOjdmS92PugBzeTFkOyRu9sJi6hTpaSgbeCfuU3ssAnV/N7DHC3PpO0dH6
HXD3qsjXof5NQ24yS89lXpZGCJv4ZFrxNxWS/LASdr8Q7Wz7jL9YDxrpZQRn
usOuFpFIXk7DZ8OzAQ6MClBcz1hRL7mg98O+fL3nF9jCw6XptDe5HSTRMYI0
wAWJuTMJy7TtsSqb8ILoUuEnIsIWqUvDBpizRcJWXbA5iKui750TnGtFvFDD
uIvMyF+xgAlplzc1IFfKtkXYbZZnQLmR323GklXO04wPHov/UAFQDlhHHrkE
ZghxAd2q6yKopFCU8L4FlCe8YkUH436hsAGjLsWjeapvP2QKyi8XQKAYMts8
DsoyH1m4u9+OtSgGK4kU96TWs3SsobdLJ0E6IJgD/qU/u+ZHipoArzoUWklI
H6Z7vrvZgRPWM3qMBHXZAJSSbeprby8DEouxNznBoSOqX24AhVjOC+Qu7xGI
VAABQLRetoY1vKQtChvfDfwqzoSJ7q/e1llomSgNpmfV9CQP7NobNvsHypY+
cXGNm/oCQ2UUC/mW+5PvPSp/DODLlxLUpYWD3yePRgD2qdnTCAE1Uq5kwwWi
PVrF8yzkYrpoCxXiChGfYA/EpPCD8NoU9dMyZyPayUGUTZhy3LNG1EV2et9F
lUTW1S7Ux6h5jdYR+xwvZM6kzotihVXw6bi2y5bYbeBiujOoLeKEmf694Zfi
6MO1nU06sOqPGjXxBbckzYD0Dyct+omZKBz8nsu6jCjFP7NWzBwzIBppcskd
16LxgYiyM5QDdtT9BdEpFuJluJktoOUnB9rAH73zPAqiok98zAj1zl6mKIcJ
+mm4SXacKrSU9hRxM0exATHz0EGyR2jpUwscHw5sf119kGWAPMFxmwT1F3jy
gQqgpTgWLM35myzx9NrFoIpJNylE2YLG/cp++gGrvAWm2dZHrsxpM8f/pWgW
y/E2sSG6KaH6jR0BCg6WS1pQwtNLk+5Ya5Tpzlk8bSE56rBQNynHsaPAQEdx
/dCT9U/79sxxZCrxzg5RdZS5tG54GZcBKh4OLjGx5KkBUvSHQu1cDFk8SFrY
iH4tKUOKKQGVsOtcOo70TJ9RbcZg/VjgTpIP32GDoS7giqjh/Y8PBgKI2IrE
Ix4tyB113EtE0MaGVtVHAAuxsWvzKyJCou9UzPnu2vOgLI565a8B1miMSzph
2aczuvFEeqTm07bFzI9b1vC7ws1oXKVbSZFqZJYuGoMKo9yzWlMWEJm8vVUx
Y8tSElxB08Tqa/gdhjRHolVdIejjEY6v24bJTSM6c4ap0ZvMsdiNJFSBpPaa
7J/dJh2OunI3zHv5OQ0cIJgcE3WtpBjx0rPF7qtwuJcFQ/H53skkGkNFob1G
TvzBok6EygQrnon2A/WsmQK6pmbl+1O8UF1JsnU0KczR79CBzkN7FSZhjtzY
vSCsn9bq3BjjnTVHbjEUNiI33cQYEB3njMsBDjcydPc01KZrNwmz8+4hT9g+
6Ew37fTkrJ5VwPsCDYKEvGyW9A6zEnXxGPnW180bmXzkqPbsLlsuzv6JQj4y
KXNfQBTDCQE/7ky22j96XpsdLE4bHfT9zK36tB4qSEgXFXI5EVPUvSPs0Pjo
3qiUMEO9zwErp/hzO2hvBBTY3/SunXlx8HUKIbRp0Y6nF19+d4HbHBH8lTt1
L25z5YdDmysK1FzNKVmVphUUmyny8Acx6tVL4bAQRNdJ8vZMi/1rBXyjBrIh
ISnUR1TZq2cbejwcWGp0Hlefg8ZIMlrTegn3cHmRAIP6oSYjn3y8lq0RkxR9
7iKi/bDw2R9IjlkNHKFvUBKqE3uAszYE4LFFbEABeRZwEKKOI2D8BjEFHbcx
aCygLkjTMajQkDUonKqpo9dJJPGT8apg8s1+exb0v85mM8dERS93xUfAoT7N
pRsQKZGcPiG9/n1XR1Xhwa6c0zGmPNuwn5n4NuJM4Yj+bSG5laGMJy8zZgrR
TZKvO5OkURP51OmciSKOItS56lm1CKM0Mu6WDhiiAP04E2SrSotReanPouhk
qBa8NigtymLLiEEAICbuqSu7rgJQIUlBVSJRCcWpjNfT12VjKa+ARf1TMiU4
3dDcd+hFiYAgSsQgMgz8lddFGy5UURJGDzr+Mpf6prolPBt5tbZX3UtKAJX6
bKQz55qiK6CvpwrHYnjJR1cjNLwSiN6GoA0NJJLrWMOMV9ZbELN9gU66+Mmj
M/n1m+/mKaplH3WdEqTfRC9TdrY8HgCNaJwMu9MMJdXbgSpK9Rq2roY7AudD
kNYRsrudgunhPbDfhoZE+sprAzKqAATvuZ9jE/HtPfP3owfecRsvYaJk9HH4
q1fzORCaWjajWkuUPu6vERTaXC3kukpiVgyyzYiSqGjL6XoGytRH4xJlx/UP
ieyTZRKwHM6ZpJgY1JDhnQ8Sd7aj3RRrJunM2bSpY5AJYdoW9bPB38Lrn7UL
S/272sf9rEjEifVVrHdLcQWy3h5Oik+n7wuD/7Eza3+V0PQSYzJfnbY2nVyA
STLZ16730nyI/ong6/CNfoU0TyAOIWasx18DE4KXzQWwUNUNRBZdY7VvON/W
80wb2WyalaKoOczV7khkeOqcMp1uBSThRecuejheGf8tB2UTJVzAq5/v2qBT
VwIDLgX+962AM7qQC/Gc6mDVg5+yOVP0AGqmZk5PFrrO9WcFxtDaZfyS+gkZ
1ufaKreyyZsEYAAubz8UDXAOEoRKrvFLMQMRkKvRdoQqMdBuGm8b2t9t+B7f
u4IMpIIjMWTynTTvmlKxFy01P9Umck1rKWTuuy0e0rrbMTg7w+bJ0k6Fxpj6
T7FvLfcOs40yXRyUn5Q0OcwoNIs6onLHcAf3hlEtXg5qPAmRb3BYST5MrCmL
cnMBA23Rad7+AbS03p28aD4hrK3ttvtjO+HupJvLP0KJ9w8nnxsrjCwSYtxK
rDCLAOpaV9AtWpdGy+LFSHWgbQyftVhrm2bHdf4L9sZ4otszeK4ztEQUjx5u
HC+VAKpnjnzwaxO26D5YFfJyGmKHzfQZhm5djK3HS0KJbJfrZI8QaAgkewA4
YijDjp8q0k7S1dPXsMdaaT5iLn9lNTh0yVUMiy9emy3AL3X+QIojA4looSBq
b2idDrf3E3yWreZEw8DsVDTqOVlYrUP2HwSmnnZHV4RfGhV+k2bitF9Guo+K
ZRJOeKKrfVlTnjm9PSdoGEBmUIRxsmN2LWQJGiUvmV7IL2jt94KubaqTYH8F
t0dq8A94fkNUVAMaX/s8awrQuFZXLOG1OUW+kZT/6jcnTsl9KqdCMHksA2Bo
ZLLkAotk2jSs8GM4aRoQbV5jQVaaZsa+GHuYXwBiN+aW+e2VBOwpDMucEHiG
6nqM5yAYha1VcyPlCm2npTltwirbPmHh3rHnijq3qllrvI2K3Pm7th6pOndm
8gDV2sgXvLwntLE8a1BKWfvydLB0KHflMkQjobecBbRMphH0o7UBXyr4By6O
lQibMAgxUS1dz/tgsXd7ZFtH94R91ztCowPheNlqTQYhKGtSfRB21NMLdS9n
SCqzLMgdRyAW5mCB8vepfXiPDCAQ+MYf302e7l3cp6jaFnCuMbtbYKgYHLn3
x3fkAewB4ZtHyBnSfTxxXhEOpnqv/eCDaDTuUi61Za4MleBYTM9gmLxqvdwN
crtOPicW2ubZwNJmNnHiTMyaOCQHKfDerMhVTMddRGLhlwgf5fBpChWWpxJI
VA/E6E21yCRZFGRGJe7yP4D7nbdDFnBjl5YbeilkKryd7+fXXTgRRTih10tc
vtTdVm0Mmz7nDUvZMmTgJt3oQxZ/RKU9PPO4eGmMK8MqYnhZY10masNHqsD+
UY0/m5THu4DAP3eezK676ZxWUNcIBDj2NzvR1iRknqLHTVGty4mANkN0CtzG
uKJABtIuc/Lvil++wReZY5ADz6tJYL2uptZqUgzSyQLZotkHYR6O9Vhlelk4
0JRLLJ6lLjHMKOTUFPMGwUe4bVXOjfqtI4TPK0hHHfiUR1E3BhvcY4/VLuq2
a/x0heGhD10bJnkpc8YcUHwI3rKqyzWXJWKOyJHynTPbTOQgKy7g5o9dC7dc
2OBOlpuucspdSd56KkmNUc4EAKTpEudHQs3QyKsb3l5eFBQZKovZnkJ4Uq3s
UzhpAJwQ2VpS6NNI4KCjpgwGBBGr8M9Ai3rUXicFgINsf8Qfmmo5yV/8IDZB
/o+yWOUFPmrRcTB/R7P8YLNYYIsUjJSrLcqtaVR8D5E32qnxxWtkc0wswNro
uIJC8VRKWXErr2YBwq6vhjk9nn+k6GNzqQFx6nYSreVSuw6e5j8UEcBrE/JX
yVGDSKnnzFRiOUqrfvt8wandvBuHr6AhlfogKz3jxnWghlqznUORG+2mGf7P
ZUdN2QzyebvHbkizAptEtasbrwb9j8qk4o9x7WcuvCAGQrDiFpBMHkGDmlKw
JAtuCb3ySIq4bfn62nLZukXSEGoFI6f8jfg7E7AzJviN9FuoW4/kJ39gdNk5
C4L6Gm6F4yDYUD9CUWRIl/Vi1QlB5mTSFhZDswjfh60/WnK1vZny8gTQtwlC
9+wMMbFHZxiXCoeZUfL0VDiT51WmFcGhYvFJ4y1WD9WhVtY8pUTGEHk23HhF
na0RE414vUdsq8Md+XNifUSWJMEKCMXV7k7/6tf7VyAUrsJsmU9Abc7E/Hhd
obzqdMUN+ap1U4kRGO8wiIxXKi0HGoo5SP0FT3cHh0IMf1dbhi787T22Jee8
qJ9EwZ2bxJM8sOsk8e8Rgi0SSZPWcl1FvLQIqF/v/ohPCl64P7vAVxUKLSqV
Zt3RRhxfMLKq98MHh+U/czxIP8U4iSocBqbwSbSjCLUJj+Aem5JdO4C5g88V
umPInhg9kb0usfMEZ9nsXougQ4zhHz3c1ESqNEPZsq0MsSrI8krCHC5O8Mnl
SScL2z5ry8RLrLnuBPJ8+uvCK+zM9/6w9fGOghchPdUNUOCiUOjdA+RaRljW
Th9ELZgFxOQKOcsTFnC0TJwpZ93USu3AjHuQcrnL6lw99SZEGW0zq0j8FfEt
C85IJKW8iq8fdnDWhbnnSeglqgGCIxataKTX3md3d6ynkZNvFwZ0CxkhsG3C
gpw6RtL14HNO/RaGq40fW7g+QeLig8lYdNIkvCqIUm+jcph1Ge7WH+4Rl8Z9
cN9dF1Ap/mkggUWKmHg40PjULfpuS/xh99MJeMjOO5tFfRvZD7tK46okAxai
wZK4XhGrXJjNuC2us2Nh0RE4t8iIZal1qH9IiveYluZUu7I5j2c/qrCyXezD
WJCEvVAci3qT/vlgXyPSX6UWD7v+ZEquoOgi6IMGnw7t58eMzallyoEp2GFa
wxQs+CfnnHe2wUo6rf0077X278gUcQsHeB7z8BZJCKfNNS8/n02zYFNhrFjk
f0MqCv7deZuTrWiIFXC02XjraZfaMuNj1GnW1iGxkz95g4DhhHCbs32sKm8C
cW69huViFwMCFakHtngwFFQJUhFGGnwGRlRIT8wXd7R2U7dX5P928wq0IMHJ
nYozELr63wab/esx8TM6VGYH1jzz8l7Udw/qBpV6eRJm3LK2o4hJ8V3+0Av2
Klrqof82aHuA8PWgwvcQ2VqgFS3P8LSMGu3LhJwtakaI2kZ5KRRm93wQAegz
3afEYWzCYBs7/8R8PxUdT1anTau4zV+hdhvfYVYpzF41Y3LZwIs8w1o9/V4S
awxWKs5TXC8er7LQNUIA8rsUOWId+/g5Q9Fd9PDZo8ItipIbA03pgZ9sSBIw
r+2tPF/SmEPAtmNjEqqme/iD4OWSFB6skpsG7thCRbbB2hoYjSfpk6SX9TAT
9XDCVNUBn96MhjXXo9bX1OntzrOtZPAkyDxMXJ9Z/XFRuSdR1gU2W8gBBwKN
IHOPsBbKdJ2lWMJ6ovKYw8aP4DvB1nvgTcyXyQmkUXf3WdNXocgwvDqo6PeU
p41dIy+MLiK7IUsye5cv++6yVxLKSyxjyjGsxNN0e7DQzqwKrTtV7ZjpHFQT
jUmWeXH3gGRH8IqT+HbDFfAlA3iv6wehjNqyBE1CO5snWjVqI2mZheqNbJyN
zXSlmWcgvmXfFMKN5QZucSrLzHfyz9+clHSeTc582Q+GXt94Iis2MnxFBQeS
tIUrXFyldNAC8Zrj4EsSNPc49srnirPNwFhsPVBO79ytYutcAJJ0t+OBfudu
bEJJgkiiyUkjOHDegeroAqr8IKuVbGKM1mR7zezMoX9HHxDYnJcHq0UItQ9H
d/BKOslrhqPHx+zhdThSFLkjGtE/y+4oDEcoXN8I8lpLUOdDOZUjk0cm6gt5
3ihf/u3kISKcOrxCw+L2xxAxl7+Q6Y3ZkOEU1R913YhOBZ6tEy6P6kArx26t
nTvKPRkqCyD3LcAacDBaZvqY3Z84p98FZYS4Q5by/gLAtjoopleKzqdG1lZV
S4bEMsrr1zfaU8J31bHX/WnZOaX0HfyQFsYdtQC0VU52aC0ikLjSQTXWc4df
bt9jT6/BBnIC0uNMAOEyVcpNXE1a8TX81W2+GLfcyiCt/Rp1P9eYLelFQ+KE
yHPaCpomaiy8+yRwF6+/gr9yfaF3fjw0pdXXs06qxaJRk4DUZh1GMjCFORKk
uNkOVfGXWOFKmd+nTRdAm1D1eQucxuIQBHgyTd5BTK6Cj6mibUQnixSj0EQ9
LhOW0svtljAzh0a07bM+A/KxD9w1t01vIW0HJ/Mbjm0IPJd+h97Ucw2MJnqh
cL9eI4vkGo0gp6R2/xL4bcYjwP8D8l7knB/WXCmnpzD6Z6K8w31tR7jI4dch
iu9Pex34dI3WPrkIu0/YVj+yvOV7KEEbbxVzsVccRkIzWgjJOLp8ePoF3nGA
iInJnSt8qGaRP+sDGiDGZ6VsrvWVEYEaOyYhKtZgFKG9ZwSIMjWRQH6ZhVNO
tHaDDATgKxJPp4j4G3+MfR9CEshIu8yEf5SZFiFSa/TtJmKnT/hhZTDHe6Pj
LJutTD60dMAUjz/LSqIkuP7Ji9vT7hyCt8bizZfziXTOTMwZfs4SGaiy0sYG
7de76MWCG4UPm6sBnMLfIXTlx0mBgIU5moQOTZXTbKaDDIsfa9MZD30l5v68
nTKOx8+gcqt6CYFvmdFJKHzE41G5rOGcb3rcCqEfw5XB0Py9WsIcEJKjWMjt
487nSvC4Kz/AOjaMsILv15TYo02Ypq/LcwqpC+sPOCidMIgPnl3kMEDryIY2
55m0eKg3JSHCZ+8WDT0pFg0gMFL6DZ+HxsE6JpB2rrHrbvMmlPHUW+VuCesT
QggCUBrYC31E++Q1caaQcExkVELU2MxK+xiRwzgwnJCaFszeVwX9qc1QzYLN
M9wkbC7x+Aj+VlHXrpm7m1qTRVgVa5HQxfjK2ITQhV7sdCGLeTlDR6q6/3q4
x8sQ72TfwfWY6dE2Y6ERT3wGDOwZWDAh9m1SLf5AvUTvZ/xzf4glM9sZEKEP
II6ZB94neS7PTayOWplTMRimS5BU/+WJJWNRHDBCD3OVlQvkiKV+njrkwLzc
rt1hOfbfzT9Ejpw6L/osjh4Zu2geTXLOhJVqDia7QIriCPcIGNo2HJHXWmA5
H7IREcRLK+o6uC2A+BGv61M4C56hUOq3T8vOT5+l/tnpyhJx3YgzMenUZoIl
LLvwn+CnwPCq7f7uJC2SLRxkVylZwEmausbG7a+Dskfciz/pp04tuEZOsqMd
XnawLTQ5Xifa/MXTjpbrKyWTtUbgNCFwbqCchAoYGRnhabP+RMEcKr/RBgO5
7bJ0UTUC/5EGsoHEmub4gg3W3zAhn5cXdBFD0qfLAn/mbwTeut0IGFASyltg
RbqJQIaRdejV0pskfixQIMT8ufi4DsuXoyHBAaqNrPx8ndFKjaSxhv3POfEZ
LD0jTFUKFfokCchFukeSsUOYImE1i3xS9PAfNkJc64CMEO/PAZOR7Zah5bdG
7Nd0/SMVzGCXeT4TL6Ey+y1mZ91OvecJvQIbFDsP3tLh7lbT3gXKj7oOg22c
M6ttNLKdZkMaEvc/ou6mzbMlh17Ea35O9/SdkY5XFOT61aq/DykyExPbF2UP
NUIBZHGyNk3jg835r6Q51Dy9SvSxt0PEeucsM4YWzIofyeuED9UQSqh412fv
SVtpo1+InNJQnbDiVg6Poc5PjP9L2IzqD0UVIsgo2Klp06oOr+3IIXAcWTC9
fZbjh2zqEsAC1BTSrgprNdS4DU+Tm7ffQWa3TpQuTQZNSqcqQ08SSz7golQZ
1+6t1VFbHrrw46m5JDuYneJ/OFgCqCGkpLn3gNizYpeCAM77QwORFja7h8xe
Nuxti8JqqEbnGaw6FIU93nkETOf1piAixjF6f29/4Zu1UgBs70/rLgNE3fRZ
q6KHgsNOwsDnC6nNY/2LdW7VQNmaLS+Mn/mGkX2np1YQvtIKyVpSF4OsqLGy
8vnDYwUoadypy0cuZ/gwbGVQKmjklnPC42cB2o4n2G1yzWCmxSJZbs/wG/Ut
E30YShi742hghicecT62LTL4P/1Kl9sKPF90krzBwTGO1gms8afLLu8SVYfS
hlqb6IjZfxvGP9QsGQKH1EzDHYLvh4ieir5JgtI/IIWtUorjzRREo/z318LP
gzRijfWa+QVR3HAJg2f66LuBZ/mr8rogSLJjE0SDZd96F5vJThO8qC49psDy
iDEOIjM8CHP2aVBs1sIbJmMNQL0YcbseTAN+2OSgtszTS/y66SmCpPiGpM21
uUYiA4ctG5Fj+KJ4DsdHMqr0FUgWCE53GZT2yh8Nk3Rz7IZjVZVNn8B0xdK5
p3V3nsvcmXipswrhID0TB88YgqwkMelvbuZfK7shQGbCs6S29fr5Ifi5jrXW
IzZfOpECVVFvD4S4FG5JbAAX6JMx+TNFfnX3kEhK4LHK/Jk1bfAMikpSO31A
s6Px2hvDxh/0u3wW7XiYOeV8tZMxY4zAqwoGy/38wOcMNJ8Ud34wgTZgYYim
LfqKuefAAWbr5q8Dim1ipTT2FUi/6beNJWhdmuMuk9/eAh7HupJ/7xO9N2Sx
FqMzA4a8sbPVJl3Fh8NuQ5WPlKQ9+datqiNH/1wlAi7vk/S6C5bHsmw9Xmxd
S68/1zsp+J+GBxA7zVmM/AcarSSufgwgHMzPiwnVzB4HCvl19wJKk8J04z1u
gCWgv9tEUvk13KSTbGUHcOvEyAMBG53AIpz3iHfZfgPVgkeDzh+nxNyGecuN
EXNWOYMcwqqmDYxsBAZHjGMCFgGDNuS56c1a/Qzt6SKiENLDLZ1o2jtU/uds
pwZYCecGxa8uLDdVtFybc7ebUS3kzY0FAtRrhw0kbVrsWZl+A0dBIzJ76sNQ
F5+GcE3JFOv0ibUO0/6UI+ow8AhbaC/VN2Eq48IBbx2TgAu20g50zzR8nq8K
B3H7oz15VSLMYHVnaksJ88uf5ymOEoHBTjg5XQcQtgVoEnj9RoAyzAELMGiE
wYOp+IbBBk7Vylj/FTny4syyunm+MO828vceMAdHxUI7yoI1pZN9bK8yLBDj
Z91eVQHeGzbRon1/GelYcSM2VdL4SJnkqv+++petL22DQE2E0J1Nxh7pDBca
w5ZLDAY4XZgDGSeKZaIzf3fE2IIqq1XBrsSHJeLVloHBAFZg0FOcCZCy+YlS
9BAuirw/GKrrFC9Qo2fT7VJ8eNHSmmTFRTKDTMZ/bEV6RDkR1JAwc79UWmJC
Q0QULlQ+AVUPHUSsdEKbxpjY9PVu9Nx2d82rMQcUjHJDe5qEScWFrEC6TQdW
83XZaXtR179pg8XzsyGsxUXaP3qLQVn7DelIhdy+44yXhScF5WuKn+KAD/P0
oWQuvkKLzOeeINm5Q7h/rEKVNemrj5+XHGeMAzvUY7vh8lWjhlmDRvXQjHDm
sNYHsGBwopfmKvuc48G+X+zWiV6M2GZxiO76GOQBS84ofPtDBXYoK9e4Rbkq
EwrpOMEj3WR/VpFY3mF3/ONpoloaEOI++zkf6Fx5ceTKdxsCQLsQGVaQjmoh
oPif7tUGgRIu29bD6fMuIHetNdWYj4SvrjXsbQRzLY+2S2n2jvH0deNR5Elo
jB7qvj18LjwT/RwaBgI/gUlMfnbTsVOwGdcDim3Kh5hhm/ejYIh4ryfsuczK
0XvHmwHH65Y15VfwF1wkvtSGhEKpHft6lIrgQb4b1F86KVewBhY2xGOBCbrD
eaS2J0VeIaNjtAKuckgW46AURCrL8KRdDa0ajkZMKEfgEP389EapNJaCYFrQ
HYqofsp6OGa4ggN5XrKiCfkyaJpGtjrzVwKEUnpZp5HJhof5Hy2tN1MjoYsq
GJv5DtbCuPvZVWohQ6NBHvaJUF4g6FhgmnExgj23DUxmc21pFm/NxtOCpbof
ppu2Ssdg1/vx6DUXzNQ+QiN2JC7ozCvM0X8q6weL7Lv1ps04JyhtQQIOb8V5
X0rzwn0QBYsRkG4SnQ+wkLNrBPr1xYWYyRV40+6CdGynqP+GRrJJxipzjcNl
u05xn7UP2bG6aEYFQwWejn+k6hQ/jpIg8U+d2WGsuWVVG/hHVUmLH1GSjn+6
vE3eTAYn17v5Vpy7iCfzhdakeM5mZNzus3M8r7h7VsRvr4s0p7V/+58Z90sV
wwzYuR0knm2QnXSa7vmUJunY3Xv6nbf6VT/L9IH4z1uMkk6QSKz0a43hMOhR
0WtiDLqSyEZo+bCrRH7WrR96Ioo+vfc2A1d83OUZhUZcc0e2U8Gm6PeLaJXr
WsQRoVj1OGZ1cFRu+j6PkpLdPdiw5qWL/qp9sfEw+ZeGZevSfLbu6AQJEnpi
DnmOYjIUvtbjfqjiaKG12s06WpU4laBiR1v9WYfcJy40UPqNY+yki7ZFPXVS
Ums6Us/u4yjc4BQ6SL23eEtfwsViBb27VCUJrZtZwmfjh9U72fjdbSuUvehA
6FXsq+DvRy6QTmQpi4diNxoalIRyGmRVJXq0lRN8qQU77mx2hu06zkFtXXh6
JNZaLh96CVkrh6kXo7i8moaLufTIVWyfNkO1f1lqU2kcwAU6DFudD+MkqvqH
MPB6g66b0MCbWws9rv00SrMzeHvjoZF9dJtpgwgpSxObidiceScCQdpbrddF
FhpqyCLPzUI6+AlkxNTZcWA25A6hLpLqwcPgAtGNwQAxXdlDJTzDn7R3fSFe
Aipm4OP4m5WhnCspC6Uu5+BRXhwycL7y52ZWoT8CNgLr/gHeBt7ZebnX+cks
CRF1aody4QVRLjYAI7Na/CkHpA50yXgErS6D6Ht5UFtAY9SW0I1I8Him/HWj
dcYriCvuCOdKi/6Qpk8s/xjl1ARMCpU8smOKg2kry3sZVXtbTizjMwwL2V7s
L9wRxmZrBxtj3YSBofCyH0+QMh/fczWXT0/A6+Wyd6AvukxbnXieZc3jeUaU
AKCqG1yycqVPxM7mHxkzh3RDrp4Kqxn51nLvHuCSFZjASdBI9XhHBlHQUFfg
tmSkEF4IQU/o53QG1lRJil4m+/902LpkUjcS+o+Jt/4lsRmIo4nyanqLYEB5
wI67Z04XaLqvtZCMzO3Z1ihbQegC6lGjtc67H/KVXhTZKcTCy0I4mp9cbYSy
sct7TXKz57f0CQ+ClRR+4DpycRu+2uXvg5yRtCCDKMpZmnepdqU1qAVpf0Uc
ov2KLiJ6s5+iKCz3SmIjjVq/1GPd7ZRvgdb6hpn/DTGpvFRVs8OJ7Y/2zlmK
6r4tK0wrZSFg9Gm7IvnBnYPp0NbFK/OauWnPKwlrMKml7ezsZCWzQuAFoaMA
6x5QVM2WCt8oV9qyP1zoC97iJFLJZAncxi997QZeubWTAyZgj695z3ayzqND
FsF8M2h0rfdHrGZJ9LDttWJ12xXjUm9N8AeaJI460G3Kfgx/Hlz2j5BpFR9U
G36C4YFQXquS3QZoOzcZukXzeYvPGPlgIB+X9C39fqL2bPd5hr2jgpEOwpqQ
tRxAknm5vyD3DQU8ZNrffL6l6jhbRtm9yFJDY9ChY/evsW2DTG7UgSFjy5I7
wjq8XLbboTzVj/LONQVmOcp+UfMhe9i4IKZirmQGM8uE1695tMhI7qqKvPkd
tM5S4cj8SF9I08Bnr/jllgFI5PwWSD2esXWaPTLSourseHQ8anKucCnDf/92
LxKJnxYZHApPGLhH6uPiihWEHorDZsMf2i3XTBXRguBWBt+C/WWu0ZuqYfpj
IGn98q+ljzd3D4C5OPmISoHw2WyC8/F9gf+n/K8Xz2ohJwMbU+OBXwvJSzN3
+ePXyMNtAdWL8jF3yvo/MfckI9X7HzAC1cc60fnvLGwQs+ms5fpVGBsBvbLZ
gXWc5dFtDCfLE5sBSVyg5dXn4Ebjw8Om35pe+ow2Er6DbR9Gy1MzVhAr+rRq
7vrJkGOgNdcPWd+h93i3nUy/n5v2gkF0bGlj4cH0qK2Z6ZwUQjwZHsGoVhdr
6JgDsFxw8FBAyf4oxm0ldBjAfMZ4ht/jjzHuH1DlTpzaXV90t7YhTkQTAX1x
dnhaGhsiKgBRbe9sIkE6AjKZzljlbDUFofhEVBKHBwXoFRjxC6TkNb6Y6tXh
V2jb0QvTFEiQBPSOqlVrivagoNEpNBt3yMsmsu/1sc/4rxuTODEzPg+CTviA
v502oqQwlfk+YNiahZcCU8nXI9WI+W+p6/4pBUsi41JtAB6pSKcFsWlsibLh
owNjgGd0ebZnHXhke2vDf+xOrbfkS4xcJDCRf9nKJ+G70vdvs9sFopGGbAZR
wYCS+OCfUsowOPRhTytAnATmdsxnFsjGWwJ3jO0Fredw3s9Hu2f7OH2I7Qvd
9NfOWOo13jmMJlSQL8lbbU7W4MQew0PUF8EhQUXr7uvpsWgJ45asaEE2VbAQ
YzeWyvUgOWo86FYZNLHu5nTcfynJ8yh5yGVdC+3Um80kc4lUHbePvGh/3foZ
y9cmtO5teF7xuVCIkOz4QzAFl+eMhswPrvaKhMoWs11BVN/pCdFBN9ga2AUU
Ocluo+Bgad4qs8eos8GkcLO8MLKlpqTGFmk6Qa9BUrur1VLszkSpTZ0uROc/
vrqCfht8yDQ/WgOmTxFYd+SwfBs0DlrUC1N49jsYtqlZNR8arr1B6yzd/cVL
YXPzEAY8aM7E6KhnQDsmE0kEgLzBaY3wVmT+1pDvXc0DPK7/QnyHei1yhiJK
kQ4ANVFYg0mPTaYa8Lhr0tklSvSNe3cT1aY2P8GPbEYWk9wkohiZOWSH+SUl
3O4mKdwc4koHBlU1GhlIUpT33pF8FndIkJR3c3siFCYyrktK/Xx56Lxirk33
kFWgAIIlHYXmQSROgGLAz7FcFv3hpY9OBKD5rwWqtwghTa64qUPH4OfsfTqL
nnlkN9v5p95kGXRuwrzgsCnmggjb7ioe0ILuYjcebbifm1uJWyh6SBEGVVJR
84yxOiayOWitUDZNZHCzdKldLHiKMchhWUBDS/NIZzIyoMvwx7l1Ndwh+Q/s
wuafuWB4PW+QwYNlNalX7QLc8p2SOgfS5hn3Avy0NPh00xdF2feA1cE07Q7/
3ZyctFhYt8VrY1Hu7NibS0DXqTIIMt5CthxEptqBGscEu60vrjsxBl8JLyXK
njfWLWzD4GCNJ8v8HcMJuVszTVfOno1H/DBNT9l67qM4M82GCJHk+UlSzvnT
LGS7UU+DbW+ywUdfH3uOcQFOS054LeWNRrDqY3h4W3esX9qTZefNhl7FmlCu
9kJvXN9UQYT5nEeLby/JJMj3HzjK2LiXfctKV82U7eSdONlFyDwmpPisV0hV
BkMFh99djOGo8xXjFDGwKkmuKIj6CjFKQo9+PBKNZLE8wev9/6YRh0ABLpVc
Mp5tuLKFJorlnfvdnadLc3cU+uKlEw673fXQ4MeCXN9zObM17HCXjmteZN0C
9SIvXEQmTTKhqpu7N2S5M9RiH8N0s4AuF1/Yod6F1uJRzkTZWMuY+hhgU/Gl
tLh6Xx/QlbKp7erPgGEk+ZpYlaTPi38yxXU/qO9U28ENPSlPANkz8lsT2s3o
SVk1uxpg4du4dK+Fi3DG3QJ7krKhbWAouxVVmGxWNakSMkaCdEew2x4rUGM4
G32kjKyXzBXB4Vm06CvesFwf2o94cMIFxTWeMnmdseF9Qd0+uuOEEUyXPclP
Gwa/O8cgay0MwfqErWntaf5KFaz39yN1GCKzg75zFYY/CeBpVoQvYyetnDp/
f2M3FGgK+n3GZKsZ2bNaWcAjiYckGvpjZHttUoXpJ35K51D2xjOAh7wVF5Ke
eORxncxwydyPhhVfLMBcrl35/NFNwGsnzKPY1ytko+9+njZqL6lv7HIq7FHA
xxy8HrcFIbOqvSmeXKYaC5G2mshSj2EQ7BZS/jj3s13aXjwCjGAtnK3OF+24
kX/N8E67aQ2JNh8NwnH+MJakzPpBCMdphE8JMfISZAYJufAiOn+x/tzuRHI1
50hAxaBESjMo+DfrH1qvfluaazDxQkS2dne1WizRtQc/OIYzaEmhXzV3xFGv
X9t2qPsIUvMCoozYm13lqPWrLE/ngXYVdwtUe+KAaC0Oxa5q3x0nnICYFfyH
p2nkHsMHyeCPWoWUIF/Qa21zfUpUirSx8iLR9X//3EFpm0biqHN21H8yYcxg
CgBL1/LSsy/iSP8bEGrN6yyydgiBXAXERhO7Va9MVHFjPtDJPfjj4+r0sj2k
GNj/Dq6NdLc3XJQHwgIt/zLJS1gGYcvjwT8JneOWPaY5GwL4fJtkx2OmjCZU
ZNz1sBdTsd2cHM6ogAWctOLfCsP78PByDe9K2/X1+JnArkUNeA1WhCeaf0L5
QIdqod32sSajEVjmbXZ/PxLfdif0wluTgrTAuVbW6r75gj1bDT3Jhe+kcPzD
448eJa5fe3FSERJzOtNTY9+Jd1iLLG0+v4LREYIQnp1Za1vRye8Fzeedy6bZ
bTApY3XJQTMueQOEEumhAYCYjFjei32AyYJI0/b+e0JTbUlgOzBsk8ycSP3M
f0KC7O/TPcuwuntUZRqLgjjRyawHvGi03BDFo/SyWofnddN7Bk+DVHM/tpCs
mz6FaG8m6v19gTuxKuowKio7ZW1/aWNEWhshjxnFk9xqBL2FfM6RPINGu3Tt
HBGDI+/fR9dbfFOOzbJx5C1WPTDQxuKL1lBLKNx6BInNjx7L2Zh9wUOEoMZT
NvJFLV/0n0yfT/d4MgDZ/oukr1QFtYE5m8cG1ff8DgZxDzq87Ye8jWqZLS+0
lhcGgSl9ZFqtLkV8asyGzitEjYVIUyNJ6vK2ifdcTP7HKU6bBqYd90VL0Bn+
pnDgci6gOFRYf60KTtHo9Fyi2nDMDP9zcHQqyhUUC9lluBGepfmUS7e8FTkm
Cc4+wEXuI2UUvdu70CMZ/A4Mh32RxsqvWfp4XTZSnzD2yLXAlZCvbd9WSerY
nYmosQgqrGo+uUpXX3nbCOWmjnECrFC4N6oMt7Pd8iJRY4rmJRk61Jlpjq4v
hiGpwl+wX+bXWS3mGUJ5UXpCSbH7SogAPJ9byBeIngTUMgN+idgxolpmwNG4
O2HsR0QFUIniwJzltYFDKOtWIKjPfmOYQSZ948uzDZ/cAdtzP4ZzEab4LPur
q4t4vuPG9s9Xvl47kGVYsC5uXkpjEHOpspDhDPii9hrTfzfISd8Qq+RC+aEg
0Kept6Y5Fbj4tG28qYaR20hx+4cVhDcy/vjAyGSUT692ng7U65+6CZ0oGXnO
ZwNmcrW/SQ2wNzJAMSQsyT/zJp9MBMkZrLsDZy3RSpVl7DhmVYyl3BRaTaQl
3WD5Gte7kgDM5pPnYmoCs5kDsu/bvtZvuUbPWddtWMvqBe8BPM53mU6jxltc
YDPdzbtdWC5RPb38oXRnJ8g0+LNEOP1vVdis9+c0zSWBGg8EETKlY4mjzMAG
xdJss+bVDXyOY997tMaqKrHxr3XfbcPBjo1isa0HyT9je8NZO4MwApG+juyQ
FJ0C/7IqyinQl2GDrZgCOj1rZGHYPYimRz0fGbcM9uKuXR15I2eqgFVhE7Rt
+nYXGvOE9ou0LTQYlxIdeR0C/PNwkuDCsEQ5CrwBEEf2LljQchGWaOWjHSqX
NGwb/KU2piKkH4QalMQkaoCXgxUPlnjsWl7UDk7V9eonW3CCrmxY15PQgnqr
Dh9wiYZZU/5kUAE/1KmWWbzgpbEadBtSe6EVvP7fiaAUXCeE3JbXUlu4UZ1R
cR2cWddRpdI4mZ3rgKYF/R3fcWUGQfeufk0AQ9IE5PlcKf2mDJbkZ2z7HQNa
3Ac86QcGfa39c/Ddu3rublla6xL4ZmPfXg7ottvbQsvs3g7hKKgXZqbRo326
gBHxG0+Nd3r/qI8xNXPxsQ0T5N90xKGmg9YbEO5JOxz4kXPB8L2E0iJ2cEi5
9zA9uC/fBmD5Q0U704N9ED1/kGAHcUCYu03vr1V1gGIkdSIB4M7PDJ48lJAJ
gQMNxUPrm03nNIqwq8Xzt/TvvPDEHsqT7+S4+DKx+Uow1rLouARMV2DxMIbp
snU0xmT9tEDrr7lSdzx7MMcd1HM4Mdqz8ZBZ9XJlJEh7FzzdM6MTL6406EDa
9ug4tXXIR1Dnc8QilXr8R9vrOudb+3DPaDtcVbBcEMS+/VK6L6D2RN5sbbfc
23aLXsjQyXRP/FM8BNkZrl8IqIHTdU/bm1tZZX+s5Y30/tJ/408Vw3z5EUad
mB40qkAi915ZsCm4HhGOPXe3o62Sci268n434BOgq/vaYOLwCwHXcEOcBFKA
70FLTJ95mi7MRNmcG05wNKAbmATraASyP4kJBcknzP2uZ20UdWgakZlC+gb+
eG+sd4eJXfkMV+zzky5Ol+QNqQokOAsgghiHGmA0nQ2cilssec+7ZiMuINXg
b9ETdhPl81K08YU58q+VJAc7NN8n5YbIoc9wGvz+tNTO2skDqYx1SyEIPHXp
396qzh9i80Ab0Oe7YzTgYoLsEeqwkBkp5NFboqbtt6w6TCs6oD7QeCumAKNa
adfsO7s38oWJTWdFC+PXrvB9nllZhJCMDKHZie3E6sKj7qhmrrvy6eQTgVtK
VXPAis/NsOaZDsO/kQfhc/dpZTbZLlsRQT0IRHCHIq5xBATBHSGssyMYuRn3
4V/F67rZe+wx05zNHEiNzBgcAy9+z+APvkSbUK0LlEME2Po+6wNQNfdt/7LG
oDvnpKhSxpuNPOmWSTXUfPxNcjqwH2N9JFj2hYxGpqvNSCNGKC93ILsdCXG3
KrZTkLdHV+C+QoafzFpcYfbURlO/hdupwXg//JlO3IWULDeUgn/tocxVdWk+
PK1awNE0EWyHVmds7+v/xxNs1qrXf+y+VfbtQNLaf8wyirNc8wCDHcxUMV/G
K4Xnqglr/RXr8F/C1/yTsATu/l5spxv+0bmay2BdiNLiEwMdZYV7/T/uieAb
NJs7L0allGoGrZdC2UYKFqcDQFCLMoDGIrc83hVurtXGJ3xDdhPX5GGP5eta
Gtd7+4Zh04NnX5lxLtwSnJ3Un2XWapZC42Z61B9KqEwWWyuwMHPv511tD7/i
GmgJZC+XlDAxOeBk8IH1sHKOPap+DY+udHL0qvyKBpLIZoC63Xqk4H0biTAQ
tz/o5djawlJdEwaJY7MxLUYOV9QJmWYCaBQgWsr2a7TwOxRmT9qjKkLYRpCO
eB0ICJ3Jor96q6oqvygV8kC8H2zXUR6PRwuoVkFtZYA7i7k7GY+OuGbMTL6k
ObljgWIpIgksWht38X6z1RN/BkQOVxR62dWZULOw7fseU3BF43itNVQNT0Kw
yw+bMzGS12vssww0gY9LMgmU2poedn5babFocIhfxAyfk5xStcgYWaM56TH+
Lu0VTuayvu/IThvNiAdREOz1kNDzN391Bg6CCEFjgF/ONU5hls/lkDedGPWT
6acwSjh6ATyLD08KaloEWKqv5LTfx6g51hyL5O2hrWfnl+wTcn7SQr2YJXzZ
SO1kdEhdZfOawDpb0S7gsFt/7AInWi5dfRCeV3Db5e1BdFIOOxobeghbHAHL
5I6BfWjvPvO1pFx4vrcHTG2IhwGqR/kTqvICO5IKV9B49vlAj44wvKj8JFbl
j8Ea3MnbprQlHXppVLF1g8MtGFpDEiaAaGUpGaJRzE7cnsNAAM4gWFphWJeL
rHpg0ZLBxd3jgIZ26lKyKr+5aX1ult7gpOgrIVEtanNW9jgMEe0t1LCDTC8J
6AEzvFRPeEnQaLHCCWNfWPCW2c9FpoXRGidOvP+yaaIxLZAmtR36e8vacw6X
xebVDYxIr+zJmiJidF16nKfyFMHsyQZWmtifUAx83co1aJxq7ksGW7oEKqRj
d9DTLMzmY2UOmKpBONKsUDLEAIRThYXmlUkYfdBgXKDTp4RcGDevt9dL1Xt0
31lHCNyVU65DWjXciemHC9SK8j5enf61wTvtf3cbCTgmnwzDJQUkAlHPBwHI
WwrCMsnAOvz5iblJ5IzYD64jpPipXpkzrAdZJn/D62DDpUsdLn8WzLdtOCrM
Y2ov8p+14Gk4oBKcDZZq+rv6Js3xTDtRA3ArfSodQGyB/jUukRS9nUFFXmKZ
6bFCLVFnzEr1RSbza8l6GXiFiTmYBxLc+ItfxnqmAdd6uPxxJstWngu0VAlS
c3wzetXRhDVvQxeO80o/18IKA6xB5O4m1xGHMuXpwKDY/lflW+thd421j4Gh
J0IO2OWrlsQrQqOZqQxhneh+9wVImOwlL93dUopR5wrTWm60mahU9HkfF1OH
LgmHaoXCzWqdpv/9/93buziU9OI/m6rqD2yEZOg1BpPnnGVkhRoOwoqP1cvW
MuM2dZ4rcfNyRXMylFO6VuSxYBCxxcMYgRZYS9OT1VBF13AA8J+xQEXsFIc+
w1MdqozpkxfxW2hytVuZJh6Gpns0U5RxFo3L/9D2+45Yy0q0dJnsuw4tDsVL
ddBn0FpmS6cx+/4i8XaVIiUUK9O4UwfPUobf6toXR/GFRm1suYo5KQlvF915
OTF4qUTMHMyBP8usdrw+qgI8+onRPt/nro3UUdRpUQ7TQU/FdQNL3k91N54l
S8+HkIbbmxe8r84grBmOYWMQ0VohYSSq2pQX0khM0qxVlHSWc6Hx7rQsqM+E
ueKclyzSr3SWLSDRHRjR6Kq664Mrr5eAFOJnhqMOB6KADpecBp5Cs21Kfrb6
93qQfRA/TxOC5viueVeGH/buhZGLctkLGe3xaUcBjqsW8X5uLf421W7DE5QI
Phzz2zHOtI7amiTNHFlMMa/c7tvXTA9STd7k77JZRs5swKFel6h/Cogo3aRl
rWDpmxdoxVGZ7BXLD+w04rGAhSmlemvG76mL/earKch6vTHOo+/Nv3WGJr3M
DBF2q/UtBv1KA0Yd/Crn3074kTUkk/MqTg5q4Y9kjtFCeBuVA6O95uCVh5C5
ML56hPJA+qcSG3odYZuYknyJfBPhauBIWkO5JZosIH5IiedkASb2Coc7JvTP
HglbeJCB/xAuYZ4vKHQk0fuBKPWNJb5A0DkHz7QOe7x0QRlTc8GhFXDZH+ZS
x5yx59EmxW/Wa/04QKS87E24j148JrI16GXJg7qcNKnZtDZJjLz7SIxrb+f9
GlSLRxg2zyS6S9z8vAEVuMUIeKwdrjd65kQ2IaRJPLt41MinaO4I6NcGpaxi
2GNr5XS4vSQ5OlGayU7owdpAzq3IOjXDKouj4gmBo0QH4MVeYwFtHDZbcfFo
ijeI3INCpvA5xsapAH0fod9P/Q995+KY3Bdnvq2SSwC3Jl4m9Pkl/VcdSerT
QBpEHWd/Q08NYY9jIIeKXp7Q6l/+lIrD9Sa2h0WWcJZsFF/YVVcEfPXZDaEC
0InGH3WFG/X3s7Divhn5wUPmyvuXSHNaDc81P9ub7JO/1PH8UCS2WVARtn8q
BggwWOveNSh+YywNykiayk+PhH1fg8wkFhXjMvycspvbfPVhQ4g7/pZgh+5s
fAPn1G/yrcijUeyhcUDBZSxIEXHiun5x4a4ax2saRZwUmRydZxU5XchncgSA
H1zAMR26qg0zI099M0MFvAAeWpQPe1thjyPVk6T6QSbIpwtFdl5tGZcrVtk7
ZGSoNIMPWMDVKbBJXb0Mb/VzJTai+sZ0BNXHpQvezpnZebVMboPhVkhzgkva
0GFPD0eptdTmBIP8REuLSnile5E9r95jV2cC6DyAPC4ILUE5YfSswVs3mP54
C66SypP9kgfj/fzOmZAmVkWICtNJKgqPd9nTc4+6gBet5mxj6BAGl1x5n6b2
eSvh0RM7cXwxJHlxlKDJrtB1nFCFRFlj0M4UlxmokMfcutXVmA7Ybp6EdelV
zyFfZeDUm7JmWxVDEDGxwy0NUdbs4UFLIC+Xjb9a5ge0AozLn5ynV6ALJaph
Suhmmzsst9K7nSLbqoaebvG5z23iZO8CqmzexLbViTQ2P2yjVlqcu9Dp40GI
7KNLpv40FKnS6BNjr1nDChD6/m9LS6eCeEcn86Jv3RoiYIq1B4uL8UnF9cl8
tKETMhGZQ8+sciye4Px5TjsojEs38vNGW2F5RscyNAEQtwmtNcBBT7jwH6Xf
VdmeyxOlrc6MsV+0PETCLuf/KqFtxH1nGKKBJoCGkhoaqF249vaxCAUBCjeH
0HRjKT8bf1SqJE7AMSrwPBXufU/xaaxl7pTvjQAhMClRbghaguN5Rldj1Kxp
3o1l8jPCRm7GK3UtHk3OVDq3RJmyj6D7306lIo9ksRaldCwCCGqitRSqmgjz
/7xnJ/bCIAjl5SYZ+J84jWNmyodK4SfCVXpS58wRlCLXgNGwIZeuJw9aNkBZ
amFljxSPkumCFzHxWjldP/D0bPUYY7YRw90RtR8W1njMrZvClrooI6cPgV4C
28llODyWTYQYzlWwQWw4iHDnZfFZrAYxfOBoHIsqrcpCEbWlhU6tFSGMXUKT
DUnUlA9BjCjbsgP6rQ2AzL1j2LAP5UX46aJpWuXJPytmnrQb3lU1ILIJoXUj
GWHRHzLxO2KBGtQ91rBEjUFTQ8HTDxbInkyUOgxz/asAANHg+vNBxSTJrGbA
KzrBtgqS2ehz+VB9m4XvWpMM37pGCRr67ByQOCNgtbZx2DU8CVkTSmmI2F+y
1bLc3H0F0ykaSFm2/e/qcb4LeHSRVrDUm55rE8J7WNvqFxRc0hEUHp9dCItg
U3/o8H6Uo26N6+wageUPNrCuIL8NS/LUVAeHtE4Ue02S8mm3b8Mh/CZmpPs1
XXECec+m5lwV+Yyv0JW93aj8Wb7g6cT8FfOex3wECEiGyksbkNt67ejEY5UB
gPSqwy9v316vDLutO8QcsxN4MRjdXjIrznOlonKwoG3k1ByKwROs5rc2+PUu
VoqEAff5/MWNXQeHJ+l0d8hxTPjOBq4rRpyLqhIaxu49iTE+p3+PEM/zaDH2
etuuC1hymGv7rsuF3j4nfg1nzKtW3xC0O2PenX9nbn6w8hgVTDy+D0lAQUqb
D6CewhCEDjgNB5l0xxIfbNMNgbVI28esvrSJxwGhp+/Q+Ch6CfspqdSP2UZg
NMzHKJ959gAALy+4rItBxYRD9VZwYdWgSP4lgQenZoWLLgouH3VsllKEZgTA
DnKRHtHq4OIgvJ6vQBsb83CRoAvungIu7IDTXr0jrUBaifixHESKG5ucHgK4
Vzu9EDW1zPo1f2zH1U0UvSvgzWdPJ70u9JotOdfLcfv6LAtWWfnVZPyaTR4X
aDMQn8C+KJTBPvo6fowYOssteTijPN6CuKk2C2tgscGW+uVcIZx38KbKkyrS
EyJX+j3nuq8PWQjvtpil01lah2E4CzzmrOh5h/OROF2RgpMJBGLw3c5BtH/P
JYNLSnwo8bnSEbZjTot23xyDZwErmBwKmcBMI8LCeX31yc7Ap2Kj7tF8Ak9o
N+9yi9AL9hIn/B3TiXNUTejQQwi8PaXoFAw7zzjmb00PhA0QtZ7GqtjgpDel
er0qigIVz1bJeKzts15BGk/12eTfq6rPQUFYuiWtIYn/vs7u5AkSqaIYIECn
tnumO9AlwMoL1C5/qH/v+g2FNCLbzSgT6/4D/9kUTX+Zjnku3dT/fNOl7hzV
6pPi0vJBGqwhPXnqDHt9hKqTdSmikpxidppMzu8FMf5oCyX40FVdE5KJEuKx
TqVzdWrr8YBsqEyTMW360UhLjHDoiVUDoguPCGiauiYBspUW+w9+PDehea1A
C+33KGB9/q6SlO7SaLPRrFZo7IhZsTqUSWfMdAOJ4Nb+DR7Wf4lXGIc0zuKN
bBAJB7LFAeAy80N3CZw73wijHobFf2l7H3HJ0QGD0dJ0nCrwhzAz1P9pLjvt
SZbMb51TYUK01Y5rK7wodPeYBj27MjeFkwaBXbxi6vt1Z5/bum4ESaMCLLL4
J+fwsW64ga22aChhI2BA9s+pIC1y3zBn/FWP/g/2ftfS82pNGrHIinSy1Qdn
tCwh9o8a2zuMOgoRVOUtE+rjc2JaWtyxOCaP6Z6YCGjrknJeYzJ7a4kf+Ztf
TeUXZYqvm42427hcPEqpWWwPo1lodMsKmTBeOLpxuHscNApXoekwmYn4l7PT
HLi8Z868tSEu6umxiUdT8Mo2JP0WZ/a+Vmkg1a9BRFDHYFy3hVZ3DxuLoi4H
ZlLUt7XHO1llhdI/e1VMryeZ+IOPXSQG0ulticerXmFc///ubdEaC3iuUjLT
EIxDOlBlnAS+VTpi7viVAbl1J8INJmLDfwh1iNQ35AsT37T+HMHZczTO+KBN
0wsyT76CnJZAq0U++sDLiDZgmU3KuTby46Zpy0oELOP+Z7P7T3yoDoi1x5ij
dgh5kXsWdXvkuKVCOwhukrtFvMDEdBVc9hymMMuYBe55guseIPAUyjqwEftP
ZeBbQzTk6V1eQFZ1HXzJFX71bc8/3fj6oHY04g59DgfeOS3GjZVv43ySP+ey
TF1qzj5YfpxfJsYGdKx/e8HTgMtocsvHeoKSjbkZqDZ1bQOcp76LZS967IMx
wx8N0yhpDL5boSwA9E+iqtvNx47R42tuFTUktqy7eJFbPqjxZGh6WD9vVeBW
zXttzWq2unGHOYmS8L0eM6uuCePGltMS/pwFVATcF2H8otewlIsyiXMMFgXg
DTvtvQhITcJx9Qz/Q3c1NAEFQK9KBAgdZ7c6lvPhK91bGsLSM917wHnmdyIL
0qvFsdzbgsubwtxgL9xoO1g9/5mf+wCX0l8w1T+yHqRfX6aY8i634Oo6vYUn
eevUe6qTcfVVv9cw1u94SIM0D5EFKQ+ogcx6SX+d+I+2EVdQgSAic8yYmBzO
trPcFWfWAnBPCJfcrL21RCFG44AajtViQMFdo+hFguDgqe2e43wnV9rFQAY3
3FbnR4nq6wmr0fP0XJSMj1RdKF+/4M5xYz6z5lz+C7IgdIx1z/y+Qi0tzLo/
QA13YE7fzm7MR53lv/us+T+pXHVlwaGUX0mlxML6WoGlEbtMa9v7dliwvx4W
lQ08YTP5pLAX3awHsalzFbRgIs+K0+aS112TPUzH7CtYxmTyDz+KPFPTn3xI
8iEduGtMN3HSKFA2oFNxM3ZRg/2WC0uCrmNK+kK3TJwNvXynjE6dzlBv119p
6+LKhuqsJZcTuz4723nTM4q04Ssixb+k5PVCsyTX1F3/WBd3m+RBsekS0b/f
znPuRILCJig8S7GcpQLQiFuhLNzH80ITFh51pn+8f1P1+XxiaD3Yb9Iz/R5s
/rtM36JsjyXfrTQ7bPvTansEzOVaMZL/4MG5GvDEYLQZs4fXd3PEy5klrOuL
DQ5uwufguC1I7spJKjFJUHfQqR+TQHioABohj3QCz7///U6wsr3Tv/RwJYuh
bUm8nJfEbFSqORI0lAMTYG2rdeI00ZVsq7lzUXt3saAaXYuPlPHnZR4g1FVh
JSZGu8aWmqBqIsFx21TojWK/Y3hq0+l4D+E/PqaKqaBVxZ+45xie86eewL9K
SAYu3q0nhRHW4GOpVV+QXon7f7ggWgunqK7vzYkE1L8n1GSwIWpuiRk4mQmC
AI9PCUccETU9QsyllqVaUnq+1DFhSC1V99aVa1fYTMvl12N4328aEk/uIlQ7
puOvOQdIaF07O5XtIobXdgV11vwnSagnVy/uIY4je8E/k4ABBf0OLDqZcVrq
XHnpRqNLR/SYDLRwvE879AEz05dQp0RlEIvx84abhxPSlw9v3NNSnd2+RAKL
og9CivBsKABIkRLk5jzPDAtnZbVsGZzns3uJAfQ4zwqEhC5oHf3d6TlRkmXE
Mw8bK6Uc4C0skwFDaXyoTSpAofaoqVrc3wjZIyrSHt48BczwDNbK8g+7VPYz
OQicqqHxSZPOj8nDTrsGOExJ29Adt71U8a7qaB5NfvtPj1NSzun44btFJjHL
x9xMXK2bfZztvX3P+3CQTPJN8lIsBuYxT5vw9yRpwnTfRvrE7ZNRhs/Ykync
okGygxiZQG+jCYFgcO3MgXbdy+GPhG3WjyrpFGNvpgNsB77YnaW+XManY6PV
JfxFcfJcILv5xsoDaCaJqswzSWYqZVrxWbxEbbSRj6o0IDYoWJ6ag3gOBEO5
wxyIBGfbt8QUBuSSa6k0+lhEK72jB1KQadOG4zHYzkSZ5/RDqievETEDkWhN
yvrXkDWpA+KuUmy+gCiKrgGkoREF/O+dZFpE/lsqOtsewwFevgvsLWlMvhmU
qVDz85Dl/cvvVgFKHNxafHhph8rwAIx9Yn1+mUXkj14M51I7I+O7hjrJ2LVV
38E9j0vw3jprPja4dH+QSy3CyNlhtgKnzt6FJxJOCGvAM3ZKZ0tB1Jzo0rAU
QXq6o9pNRxpd9PsWlyvC1kGhQo9Nbi9PvBqmZfw8cV2+XEP9Y5SbCVw9DtfQ
epGskiUvJdbZG28kZARMWadCXIqd0hKT6gz55O5CCXdbCV0cB8iBmfltZ5xN
Umtl01uKjmvHpVRUsFkHLrwq49wu8BOs70ZDpwAkL1OJoQRfWc+baRSfOK7R
N+lkclOquMpSLm56trMPFpJJJTP57T6gohCW4q6Z/aOsFqIfg5zdPKo0keYu
xfFaY+tZDG9ZJVm2asO8BFRHbfpGRd2+roBzloGsoRH6V3cnUsHPkTW0Cv7L
HKv0iuqB+9vpqEojAHce23wUig7c7MM/UKHNBISAU9Aig0uCff8u5eaY975r
k0oQ6JsfIddkuuH74InLl+lsEi5xc3HWapQ7iD/vU1DzmhdTxD1qRS4ejG2K
6kT8icHqGaxPFWnPozNvPD39uPZuYWG/mX4VH5Mkj+Em8Wiy9ItJthK40UI1
qOHD9CVJPRvs/KIoJmEMQGud7a+QDZeXZBDdVAfcSoNp0FteYFnFpAXcR3Bv
5sy869FC2RFfCFv7YYz1oJ70QV3j54raSF2dRpjaRv+hUPmXc+3RjtbBCGII
CH132KDHdnUz/I4k58bFjhqNt1zJMbhXX2HasN3zb7XiScnvDD9vSETXSgVG
r9hmw1K+Y8cG+Z35oEFoxkaKNbiI/kgPlwDKU+IQlDBr6aBWEcJ2V1K+wDIn
XNrELB4Tz9D26/+H3mCvTKlb2myou8U24B8jL4QRWLLCQfAIWITZ7swxwJsr
Gs3CF6k5dUZdh0WcmLg1OzIbWOrUwOE9PGEB56ZNqo+X3dEfj3AusZFWhlQj
Dd/0dV9iHtxDTtgNu35uCCKZS0RRmi/43ar+LpFEqKfRDcmusS5gx1u+vhd9
I3ye9U9VMLLF5V6+KGyTVuIvTXORVoAli8HC7IGs3Li7eVkRJHOV5TMtaHMN
Px7GBTAUdrqqPBUPnsUiIMk1HBE3ij67VZE/mTRbY1HzBHIlbO3pPCux/tjh
H4V+zxhBV4J84wH2Fev480AapNkB1wMqLvwXffr6QacB+/fTL3WI9roXUg6n
Z+ZrOHOE8GBsuXsOORosPQhIMJpZKXu2yCk54VmpUY/Tz6tbe7M0CSZhGpDF
c+aGKE5mP9wlLTvyRagxMmIF/Bte8dqJbtQlWt/sxlI4ZGnjb06a7Mo6FImI
wgmusrjrq8pgIsaRgOBpKdM539NePr2GYRvuL1g9DxepGAUZGcHjItCJgMgh
66OwD21PQ14g4MTqXKIwKXYhCor2JI2RU0EMLuM/2iBdhZl+wmH+dMXFynCn
FGob4dES555TRHHm4zwXGN8T/tU6kKJmFgGvcpYHgZMcQkldJgllxGZb44HW
Gvvzvw00aqWrHWYl1TPTi3N/eJJM7Z2+CdpWQ+UbuqajTx6BrQu6qFgdVnbK
W48ikCO8wdzofq7SMF+KG7YRmzWgBDOeMS3dC3BPM32b/WxdtWYeT3TTeDQ9
Pb76w5i6sP27T5aOznkcCncYMkxYKUqRVH4dYLU74T+oRRFC1XOK8avepz2+
jS9FBLiy+5um6Hg71YuK8VXbSylo8OBgLsuuewBjO87diz7fw2LEXPC7EvsK
a5b98gng0vdjjChHnv0Cfjn/z+vUpQFRudya+qn0YE8WWP5S6MhoGix1Js+c
k4edeewk4/SeKjGxb4iNtEyROgjqYpBsgJ3jPw3PmS4iC+BPCYuWa8OBRVCW
/OvCoFIi4wNmEq27UkGcAefSkRkOpaSsSwbgP03XUDMbnk3W3iJzzAg4eimH
lA3jX3gWh841HsIMR5eJRTRZDEHVGTz35GMxHCx0IrPOvMXqg5MLa7laQdsK
QijGWTFyR9B/9GRfieZTbHlfbL87xWV5gj+2HqDv9xjjKCIFImHpxbGbkauS
NwQS11dOyM7bemeRkxpEn0OmJ+qLLZi4TD+M9X9n0REcEaAHHNSp58bfduwT
yYEh8N5eufpjjEnAEkIU+kapS3B2mODcmE6D+5TdfapgYmTANi2A5M2/6b2W
+VTeXGcnmx2NmlwzXWEEKpPH1AIFuzAhazMBmcNCO7HDqEDN74VSMTKDMJvO
Z1vHhvHYHo8WxmKAmeDvN8u/RarpT5YS4eoOwaZSEWcVmRHO6TzTNnqgsMLo
s7NWJSY7SYnIrvPqDuJnOnLH3UMm8aryUlJPzJgfa20RLuufD/DpQt4l/QCF
dbv/Iv19ZAGcrKIZIa7zNVRLIGaU+aVyCutgKR0aKl7dDkhXBqiKikG/YYlq
6r6LlVTZokuQ6zO3EUp3Rj/BcDziGuAj8tJoP8fjM09sYiv1bJk9zLfDZw+c
rPO1LYbFpCA+zkPu1RmAoPSqMaEJ9idm0Vv27AjjkjGchJ76jp+nrgoNXvsE
XEgs0kYB6FAS2KQQSB/npVGv4Su9sXNkBvqzup8oPfoMRcoZy0UD9odwzQt3
Erql4JtAYNvvP7JWTM+QMwrtQhAlCoUEKSOTEzOsT9M0W1H56T/Y3RB8KEwS
HoNAIp8P0T9YzfmY3jN0xMhd1bi5MWsZshHESnyaOKzSRGnzcqQzANiQ9XCt
DPOJnHTjPvFcE7AYYojp6pLopXrj88l2sPZj/GZcLG6fG+ddXRjnBpE/HGTX
G7Gdx/6OUhHUqFz1RVYKKhALv39l6e084z3Cg2YAF0XBc5fJty1cg89E3Egu
HlsLbyDPOSywR6sFqzFeHVCet3om9b0pxQWBELActvuy7thwqk0Klot/7CFX
2UpKqMvFc6tGmmBtROAZ96zwGBP3kfyxWBCF34NrdghQVKpqlz7h5LjfdFg8
1KuB49qSve26eNXCu1TJJ9qJTyCKzlyKGZQ3thUP2ntPoBV+5CXcBMLx8cEy
Xz6AT8ejxzuJ6/eu3vRyf4n6mbCs1lBpwpIZI6zv+h7prOrtNs2Ib2+AGErM
rPD0ia88zbKrGeodH27uNFmy+Who/OcVX5BdSMdOPmsM/puR2e0tfiu2yFsZ
d6ubT4ebi9ShjwLBX5uGVZFcmhjXiqqaZfQEkjreQSZ/vFwJPUEu3K915L7g
eMzo8XF/HZ1/rIP3Ebh06SfbsCjVaB534rnZoOmGZWP8p90n3+FAbyokK1pI
QhW0S9sTGDTd3a20Q3xPS8MbB+l6nuO1SPhUAfg5RXE6se57/7a42x4v8owe
dfXUTsyB0SCxiU1K/GmOb3/duMNjGTTPnC4/MTKeVw5i5hvWKdH2aXwGYPhZ
d9RuG9f5qN64WBvzc/FrnfnpvH03jLMsZ6g5auhd24Ift8jIubh08RkKm2+H
N8X8Daw3UaIUhXnbJa7Jnedc3pZ9QVRMkfJoMHcZSIPH64vOUqsj/W8Vp7Y8
ykVKTwbAwUnnxz4BMyyagSLL6U/uiymh3p/b4v8I6dBAGvy3abSq5ilEY2Ng
7sMwb3fYfxkH2oiqipgySaQk3U34MbUW8MhSfha/DBUD7JT+sM0qmrRoX93k
4FkJW10WzrXrJx3io3gecyhrvMSR/V3/p266fH+sib1KORzoKunFHF7r2EoN
6oNs1u5LD1NeOD6B0LnnXwZHMkWxr7xs+tlpTW3eDpQmfaxHOdVogdHZXZKg
CetfkWwQDC8ZvBQX4OXkcXv/VTjavGjTGEwjddo2I7AneNJtPp+P2pS8SV5P
E2BONhLcLDlH8gJ/xOggKPMIJMggWnm7H6dC44KPsYLmTeJ1fFbqOm23jKrH
BoMVfumx3efalO3Vl7ikQE7zqT2joIdwiHWCY1uvAjqb0O8OS/lCHJCT6W8o
xOPKF17h9GFNmNgQEZreKaq4B/PuzTWi9jq5cLxXqMQKSYO4u9pzfF2pjgTm
dzgzBBs1V4m/N207AMZKgFAsBm6lq3GaOTCQNkGd34YFQbHlI9Z3Ztuh4U8R
CRjUqvONI7Pd0H9aXXfwy6moVwToQD+o5RDiS/4ggOSHwECUN2uGi0jtteGQ
NPqqN9m8KIEPur9IR4YOPlE8gCATfn9UDWnLn3zHp4Na6k2QJiOfSMvQTR/m
cV1u+TEhbzu0cd/ipKp7+YTQ2QtWv5uQMlCjeRm2gK3qu6gTnnCMQuvqK4RN
Y33ImjSL2C+ji5hYNX/T725M909RZFqqRx8AT6WptTSDXT7uI652Ufk4CBFB
SSx1Mp0L7rXahjlOuqUX6aDlSYq+lv7UGZ2BSKTh3ByOAyODx7DUj8mtfHvv
3uIHGkSF4k2KuLak0lxip74muk+200I4bkXTEpzmmmpUQ4Cd3HfQG5zUDtRX
eyWmZFZFHZkTYEuAUDIOfCa0I4KvJWqqI74f4rvfEj6PVzr7MeTMfyBjgVdv
am1hUwU7I+sUTSvftQdyU1f6Z2zKgSTVZ5kNzFRAYRo6Y7j1EcmEzGdVIn9D
Hyi6GPvZMtDV88TU6M7IiSYsDT37FLbA92YX+WoSVsnTtGxXSGs/T4QZJcb0
2xcU1g0BqKgrRlCwP59oGok25MchrDFl8lr+m1aOHIn7jpN1PjiSpL14vrKv
0YbnCy/KkRy2fmg93aKGY6J3PRbZ1WSBf5X2MyPA7Qqpv6aYfQZT2i1GBkpU
HHd//VV4QHbErpfeFFJqoUBhMYpaFAZ5IhzAnwknWDh0XYPXVext6sNm4nEK
WHIwQ0AG/uXlszj3eW/rQaK8s3+UQvt44wKxVzcAHfzNijnXaGZ0PvE3ViwU
HEK7UgraaxbPzgxlZ0MBg2ljr4hOSxasLJcTz5a8gg0D4m/lgrsjsjBiL7Bg
rYrNtd8nY2yfgIvWc08SNJ9qt07lLJllk3kf8KpmGpXlluXeFY6vh/BVwJT+
tmNU9d6EW7+n5n4MDRV34akEvzbKP7Qterh4v6JbYGA21cBMAGOOwbZYQwUd
yJb2WfXAEbDYwbdiSBFofVudzEczzhxiw/nU4yM3mKEUqVZLkasKxrYsLhcV
unyIJE4QChADmUu9GpSy36BoKDHoSbbn4CcD9YP43LI/qpOwbMop8kZ3ERBH
4iHdq4sv1jP2lzTQWh23U4SUukeWfDUsotvdrJBWFXNKlz4hYhQ1e0bBQ3hG
y3/NZyLgcnvZhirx43fMOf0eYUaE4rRNavqwLvFDnZJ4CRRXvOQc8Lw7y5B4
r6tr+6r1euBR/9EiAuQMbI6U4fIWAH2tak6vMSLuecyQnlejHcpPwew/LGb4
LNwNtNohQ24TQLZjwZEPvHPShYfBY9pzUBd2WqOLOWKDR0OwsDA7cgZHvKqV
e/jEhT4PjftJthtOpnKgJKUX0HAOtR3j8jDLIK9BxENaNIZHRrylCw7IkGKS
Y2uBZF/1Y9mvLYnsRzMqJMSS54bI43UL8NwR1AUqRDu9IxpmSI7BeL1wrhWc
9aCyHUyYlWc+SkSgET2SjYHspOjaNZjsWe33IsuF7FhqcvjLMG4JqC8EPCui
TCdMIdCN6Kpa38Pu19bWXe22482GU7wiGfBWe7wOA4zOcYHUTeW82AUDQgvC
aDfQ4jIXwkJvAnbpKHAgRyzxdLelafvV1is/5TMMC770cXlLMiaWcr5++12y
+3xcZTEHySO9DLs9Gd3WdU0HULI9TrMedM4p4Eay1oA0gThIEW4AR78N5qbk
ajlUFte4tVr1jEVIiYdhgvis6M9jPDIBB7AlrOAv2hF0IfI6rh7jcDPc5FGC
j2WL/C8ZZFG+S3K0POQXQZ6+AgMtaNLnsBgEUytJX6bKTbE1AfBV4pLosPjQ
/gg2+lLfhTNjLmo8A3RhdKmXWIrKjT67iKORAVgDNnPLoab8813FGMf7jQ07
A/i9l45r8CxSXHqSp/+TgwQoce5nOQ6uaJba9MJQ7jI8z5IGxMfkwBBE14OY
d5No5vNAPVu1EmiGWPpWs7Fzff3alGSGrVHq1mypCWCTycI5lA5ntJgl0+9A
GhrUW67HFSeiL9M/0vEN9S3z6CJCyPZGvSeuRKvjkxOs0lgr4leQJTlgCElX
Y8mysRzqRPEtCmafjdr2U/woQUDhnI3Wp1dcdjunsLLZXqW0q5U7QSsr65At
FzvOfQqMDdapDvrNUNpN8m9Ur87xvrnPjP+5nMJZcgaJ0lPj9a+8mjVsL0m7
z5MYP4SdIZGeoyEpC5vpuA64qQ/iGXjXXdLEfZyEuO/W2O9RxuhTo6/xUO4S
+RoD0wn74p+TQvWnMBvCo06pRNEpBdmPhF26BzlW7CT27LZEsI2f5bh9VcL7
V8b8dSqCnPT6eFBShKVfMHzkb5/2OALeYZkqJ39kib5pBzrgTaCNNVRzA6Ns
ZcV1lqF3kwuvZQB8idcKuHvLzXY+yP8CJM2uYPgDQRNDOCJHbfObcGgYbc22
9CE7LXe8g0+GsePG6ncJm13DTCypsgf7Qi+fEfIBJbG5SLYjutZxzKGT0dda
tOWeCWZV23SKkdhppGFWnGpfuG3lDmM+xz1uqvjPIn5QAp5h0x5Nj+ClW6ei
SFdq+0Y0e0QDl+M3sKGXgY0LQhlHyV0qv6nPs767UkRJMWlKmCbaGL3Uemov
fj2kxMtjyrAan6WSmuiBr0ZmwggV/nQ/DZ9XZPjsZqxfJmBm+seD3wjO2v2F
DPvIQaeaKqb0p3Ccf6avJiWMmjC0+PImemBZkPnTKVJGnlx6psVhx6HZF3IA
EwIlD7qOXj2niq8MgJJQLCz8UhwyQHOm/ztbX3nPTXc2ket5vwVjGkYGH3A4
B4iCSGyKvAi7qzAbb9Td5cYvdPsg6LITxs4KmhW8hZGl3IVQv6jPwG2uJaiw
37k5DhtzOlRbfLMbc40qP/qBeNfA6mAvx1gklCJqbkaSyySNKE5dEVhsy/34
I/XkQw1ClRl5mi0GGTX5zXgZ9Kg2ogPcVpQTJWscjNFDBaqEX27UCwLwWJAO
C7QrlKiC1tJU3Vk+34jUgKz58uW+4KjSR7dIPAVEAmELm4wLSFfcy4AZMMWH
CXX+NV1tyiy8CrFdJv4o1o3yjfPKGuF+VHNgBxt3/l3oGcYFw9Wu6gEMrqmL
t7s23i0lndMs8b5MBt9dVq0Vx5Q2C97+WjXbxsXJ1trsJ71/p1jWY27SAu5L
xZErP9ZgaDCY2uPDCwWbx47EX955iuSCcTaGl0AbQRXFVnlf/wU7kFzljILF
5d+F8cQ7wFFqVHKq6HfIgORf3ODOofpdpJnv9iyVB/dkkN2fzoy1uyRHo9lK
luF4Ro0BHx0po3Tb1nf2BlXLRNd5zC+eeUH+q1lEJIy7OGTRRcNFvaHlQH6u
C75Jf8qW9qT9+22P6ynAhUTJLolVrVWS2HIi9lfzDHKD+San0iWR5y/g0udG
YVU/JPZuP5XFuwN7RUBTb6CvPQrEaXK8nX2oAbcNTho3A6FHzmEP4id4xucr
jt999ivx00cGBrd1/E9Jt+8zf+1jyBPhT2M03nCXrbH2qZ8aX0Cy6e+pqYCj
er6YRjig5iFyCUVfjXjlg2CSQORhf1PG+L9KifVPjgclHv55raZwmixrDSRK
JmRKDlsXQsiEjKsGWXE7PgHrhWD18f+CePPTcnzUXigEeipRT7SpTjHNQj0I
gKHj+kP7Rj2TmAu0886uVabxzX6aK32bWy+MlwNGCZQhfZ/w2qMz1HlpS6GW
ei7AFBPbv5b44PiNxZwpwxRhG3m8oWC/NimrEqzewXsT+CZOc+NB1uZHDJ1j
CPWGWs8XonI0Vo065O9VRvrXhAnV4z5vyBdZ10HArPkCNv6Lb8c+uJx5dadE
ljieh2fybq/xPGaNE/lkv7aeEUw2+RLdsQYb5gpTkhAUnDRCwk+QFZIt4Lgn
YPaNsqIFLA7QFSEMyKnwH5fx7HFHRQLJj665v6B8g7QCPEKpsd19PVjBhXn2
g41Nuanfr2fPLQ/HjMZ3H6wpr5mFJQcyFcjtgkK4J6tqDcBeZRDNG40Tv25q
p/loa641R2TUmJy2yN18Qi6G5uRCRuOSuLHIazFxsv84u9ZyWFot4qLCemvM
XEtorvs5oX9HdGgFd55fOtIa45N1i8aj30MA2exqfnKfGpWEgkXaWLqhXCbi
9bkHOxHDHJcEyhW+EC0mqWvngUhO6Y3Gt+0VpCMsl5nP7iF7Knpp+FjZVuFl
2zKIJ4EzQ3e/s5mqN20fKAgW5HwVxBQ4i2vvgvYaBCEhjiltjl/kzWVrnlwr
J5W3wLsjtX7Ycn9CSNMd0B/5AYLTFlBwFRmBUOImNrzDpbhiS/sngOUFK3qT
HNSstLVbM/jSv2iUXfDsPam1zOqXNSisFlc37ZxhVkNkCo/6/xAW4PdLbjoq
phpeh4XmLuYa1F92Ac06o5AfBqSIL6jOcCzdThT1EXIaHBsO/HvfuA5g19wx
UPfuddfYzJteNJID0vYYjzTfxsFpIKh6MK2SQjaR14Hmdrm04vAYK/DZqt3v
NGitul84cn7sh/o99YL9VbNwbfqK1pKMa+zh5aKpCVjIkdfHKScDWF6yCSmz
iltHUoEO5NsYb2zbizYFuh22Ny7rdJ4bnV31xvquSNtZOI+sYB40PuKO00pe
GVokC9nfMjvF2pjqHOJAvM9jE7wmJUGHMZqnWbg1v8xYbzBtOcZjinp4bH9m
Ez9Vxx3nqO3l5adrSm7YJB+CdffIkVFVEMZ5iC5LkmgwTD9ZjFEbUFeHRmDS
MVcnb6+r5so2dQhtCh5UVaC50i2k2InARaFOJNgX4IGgkFoshmS4349PN8o4
oW2tm5qLQGIxx+xZF70TmIIVA3gGHiGCBfsQx9fuIIE1UiaqT7TZKSMhxgF+
fg6UC87aUZ4mMkj0ldI4tnHZIEPTtIVWgAZr+gj3wfaTth8VzO09HjVKLurm
1RYXBGIBWmxXwu8ECnWwAgDLCRcimR+fRR73WzONIzaZ8an369mVElQqObZP
2nSAGtdUnfTwXxFU6ZyH/5gH96saHKtQlrpw7/CEmQhIchtMovCMbzeGFKwn
9OvWD/2+LHpsV4ImJVg6Vy54WDJ1h1vYOTJH9X5AZc32YORcIwBXSqsA6laW
MyL8SLYhV9Ric18URJ5oJXKBgoACnthmtLV8c2LlIUBOCBcCDax7yRIt/tNO
BjqxUPhHKEfv314XHwYLKxnORne1uRovJkZBItCo4fI5u7RulK1UP9h7FAYr
e+IfpX0LCl15dFpEKNOYgjrCYeeXyzcTdVkCT8g2Gzq1N0Gl9rgElpn1Rror
uPuw0NMsJVMAHcBE0jeb618KuTnfStpezLGkr24Mb/vBItKfeym3kNuDZtHT
1GVGZvrc0UNjXsk2cWcA2pDdrCHGMNzrSM9RMo0W1Y0HwIXUZ7mk6NCnyWob
olA+VxkTmwFsJ20i/xeFKCG6P4+/S9ADEzlrLFUKQfxpwu1bEuD4O0VMz9f+
CeUOwYlA4idHUQlwtDSl2OenGzNTEaSsvG2/ndOpvS5+YsU8yE+5udRH/pbm
S9Hgv4Wb6Bt4m2E3+DLvOiMrZ3UmgEnPaDN8SHzlbRM4q8lsKaWQZAu0gz9O
dxYoinWHNVqU80JGC9XPgwYx4Sf3sMVujpynQiomtXhYXF+KDUnFnCoZSj0R
WeXq2uC+WDGgpVv4NFqqj7hlmJLE6sKBWkIWsp0h0ZeHGTSQYY8wD0Dtjuhv
9S7GLWgUMjGIl12h5BiGBJyMLFb8PW6WbyuiUk0q2UwOH3uKtKqaFUzANSaw
+3SLtBBlttA/rMGPHEEpM0cX7Ah2O/tYu0QU1noYpcVcCZGE96o2+wzb483Z
P/aK/hJZcrsFIZTY+OMR83Ph9fhyKsy/ygasK1dz9zYexZ3CPVb2iCyYIbnK
3LlsWtv7R4BUuCWbNk/cK/wKBbjTUIUwacQdIKuIGwSnSTaVo5ifv+2c06A8
gAe+lc5rNxxL0AneIElyooh3NeV3KD1Olrizbiib9wKwk9BEL9WAqeTbgiSO
q6cSFroVeEA9xPTG7rR8dOq6+Wnmxiv9tkzKaFYz0/KEEZYtaOa+jBADxgjj
RaPSgpCGf7b0m13AQTdh0JdaMdnUzsN9TcXydT1LlVKREGMbKLWKuFQlNrkv
cG5kevrmpad2ROoJ2+lDuyIZ3ZB+g+JhVuAK2xxE4dhYfyPZteLhrr/fX19D
VHPY4Lxy2Qf/BUj9ToEqkbRvJL6RGPGYZv3vFJSY5se8ejoESU+mFu8bCwau
pAlIA42Ws+DY1uiczJeqc6PfxG3TDbhWEqWbiiQX9hiytSFMnb+OgeyPXUKQ
gXJ/SFZrqW2C5N3YOwQ151oLlG8erGd0VEMGsMWA2QN5WqrLqqaj9PpTVm71
Y0LIRZFAhI9kvQWVDj83Q436OUy/2fFaqpDbRe27EJGIsZbmTWFvHQx/dwCw
ZFN5xJo4uz2MWArrcHTUK/plnLps/Dk07tSplyx9rLEpA62XDF4Ly5A/h0Bp
/8X6ZN5irn/VPVhPflW6exY450itmfKyvAdGIKNuFytojpU2T8Y7jj3QXJR5
N4BZnVSfShNHCodWAwCPAkD2/KMK+g+GxXHYdQhSZ6eyS/eqfCYaN9XRhHtg
yD0OE2aj10D0tiwMC3nYyvSJ7JNLBRfAWRJ8OEIIdRQl6IXg9fw4HZCN5FfU
Y+a/DJs5RTlNed9HH8/XpcAJjSVsC5jQfISdvxO4akD/8/ZsBsIT8AWSPf0L
FgmrHhy1LnL+No0IgdE96M3oqdNeEMnjRqvuxX/XsPxK2fnLzhPuNVXJGgsq
S3M7EcMbUM3rxTDvDrdiHtVjP7AZs4Jg903LKn7bJmg28JT6fcnUrDMZFSUt
cZqBLq6EPV7OaKXCb12RT+tgjzxuX6FhSXleavwB4u5dPFB5HmZz9SX5WkaG
KkER925OtIXc2lOrTQ6CkFMpAoEm9rDhf7aGpI5Vem33QEF2SItbrtDbcdPV
zb+SLDS2K03Tu0jXEUUDTrcJpMBGmHpBu1mDUB2qusUl4v/TWLwPvvAoqR2B
ozCzRp6VEB1f+wgZ2IYfDIRzuNxZA3sPokVFLKadFmvM8zkBJeBmgbPEioyc
WcWoTI/4tOAfP6T6T6ZCXgd1UrIWkl0oD8jpoDPA0m5q8qCDhnIqlnV4kc88
ssLdjieHpPLn9z/tfStbiPKg+NH2gLdbDiOo0n13hAMheBRq+wANGNmngEeE
9zxd5dEdavWm9P3ZQdx1Avkc1jDv9EUcFvXL/t6ZYCoM4q/IPCr+qgUS7/tL
fZNLpOazGHZZFRt2Ev3AyMLlFc6sTQtSzcwtD2hkZQjDvbCubez6ILINBs8Y
nbdHEOB9ukSyTC5fks+1Z4iD8TkEwsrNAN/DlQGb9Nkw0SZra7Fxk2QQxn18
Yw8I+swoCPHbQuTxzJ3uci7ZxLFbwhu6RCr+PI94BqhzmWyhlpvIvitDlr/E
54nfH1XZRv3DnzhtmUj3O+ALtm5cw3x+u8dL2gCO84C9nYtze1idUrqMTjcd
lVOzvftJYjqqTwsZxRstWmjKWXMpGBlP1tXam6xPZp1dG9wSl+UqT/SMfcmz
9rc/WsoMAHxZmMPreA2hRalRgCV8YVg8MVbsbWG4OmO4ndBm+3R6mXNgSK/n
cNXrAaojTT5YB1oF+Z8TmENvb4/JC5Op2pRRidEk1BqKrZWOf+2Icbz0LLRp
0NmKSrLhZV3XFZNe02cbvJIZ/xrIxYjS86p1/0NHJte9jqW735R5t6f/wCjf
quKWkOgXW2JpcCQm9AEpT+SI8yDximUyvI4LkvHFZAk7gyCEQXZN+dzxDAwB
Y2oFu8l9ADOEsZVAWEHeJfh2z4Y5lwhScMYzgV3nlwPRDDukMKsUPOy6Bl9c
89g9N6NAP0TQ52a0quU2WpIc46KGu0633zWdvRNiURu4uW4AfHiX3EVKFZEC
V7t4/36G62muObmk/IfIg9szjvy+C7KN5qXrqJvVEYYgeBaBwb12/Sn0dfc9
SnwctR4CDEQHdIZ8vD6DY6LVLlHYLJxffmXUqfeNcCoMHNlkpVNZZjfGFAiD
4aUlhkf+bH77MwbbX9kZUOrsbTIHWu22RhnabstTrVbi0uFmZksE+ADAhmJC
oXNeJS/IViQTxtYiXo7gJBaUC/NJFPi9Ot8u9azigvNmK+lKZjnSH4sW1OGn
pQ3eL2rTG4KpNBBST9ZBnFquwNhMXXKTBPreILCv1iQBIoucDIL+0u+OVUdm
sZCN5KUxUwGfOe5fYOU1nwYC7fe/p0TLzXUyazNUnr7h9kZFRZd+QJyU3EPg
OjkVkkKSxcNLH67n4AU9EZBnlEtg7s8wMSY/WRCS7SCBXI2LBAxk9joa7IbW
ZAMewFnPAf4DtETvrDxOZeNVKwfFK+VoLDDI4cw1HXkKe/S+mVFcKZovOLFD
va25PajgiFidgVmkCAjhch+N1JQTrFsGF6bByV6GC7kxjBkuTTIfrDeAd6Ut
7V7gLQ95t/H9xZBrDojAdeCIvdLRkN8zhhOnm/EeK3j43IcaPVEWUyCesABF
SyVQZm3sUy/4L/IQQuLcowE4rjmz2RL7gdUv6XyJ4fvqaglnZDFYWM3eKBtE
Fm+rcGyvfx2NGG0OLBMtfGxszwTbeLRANBA+PHbJOAQVtI+rcT2ovhdLMe5l
RFYr6sSKFq7n5u61LrtzsWIjFVwZ2RvV9zn67QYUcOJQC9UEGIdBP1Jdq0OO
n2iJpXl6IjmMysca5792d1WO65zYqImy544dNLoibhywdw6P2e4im7swKXDE
NcMyrK6s3jDuYina74zD5LTt4BmRRHV+Bma/LQUeCCTDhNoZy5r7p/v9RVk1
2sYQlH0+tbqV6FdesM1M4wiQ+oHHZz112S7BpF4fikJrV8oIPazMQMx6p2z/
Gwr1f0PJCBzZHuLiqjCetOypoqvtCnTWLonNqg8nSEgQwEVHEcJA5gUGW0TC
A60pQyNZSC2zB5UZh4PNw3i519i2WFXDJGfT+qdOHdqM/3AGOpEZElsdBsiY
v4PN4iC6niVxDjuAGOZ1sKCDibsIouxvCfReP9rYYpSX1owpQFZbUmqYSwUh
IYN/VrXSfx7iu8AckxMAXgsdjU2uiy6P5wrG152DW7YmdHKKZtYvrPC5N+Lf
SGw37Xhg+GqcD1CTRew7XdXajPP6KyG0VvUNCOrOQdi2+RYyFbRv2AdVWNxi
WX2txKuweJNJMcvptkXAnsZlgrLPmzVNbzoFJhnJXS41eFEdV7r9C1QlvmIr
2J2SSmREFbSphbj4aqb5iGN9UoHfgGd5LcJxh6Hgf1xwn4DvS68cddSsE2Wi
pWIo3P2/emAQnUOx/ZaaiViO8WnCq2eMhZOmJTFgN2bVctlaiv40Gbz2bDov
uovLpQJCVgi0PyGJuR1u/iO9U/T+UW7uqe7XlZwnXGzMEjNlqtc7Z8+ed6If
oyQBlK+GX9yCeY9gz7AdrJY9TkvC/tt9h3othzvYnw+nWnamv27zqqKJZ6YO
6q4ym8dKyzMpEn3GXZDyGls17sNFqT3doLYj/p3KjVT60dd0yLEnW30n+mMP
nOX8xGlJJwePWAc2FO0fymd/E6HhCt8ScINVRxAprGWMyx36hWgl3VgJ9pfI
WSV/Q1I0KyQQPuxyYUPlXP449AZBdRMDd9Gubur+2hLAg9sTC5GiDjp/uME9
7XHGjgRHLEbUmpNGOGlynBwNKWoWmw4DJzkaqdGbxfNAi/5TYmDRqnRJ8G0s
nyOLyDBE5NoUy6tE+Cyd/LxCHdbO0u3x4KPk8BsIyHT6dPj/TiECyhoPwrm0
8puAbhhwsn11WVHN3s8wFWtE08oWAdYO0Wn1zNupR6DwsjLjqmPU+Y/lWNaK
ixKz7UhIf6DI8Ev37GbLKtpgIvufOm80Ouj/Y1AjfJR1Q5dKHvJ3oKC3QOXG
mZCR1lADbdV3RbVPrBdn6Dvqcg/mPfJrT+vNGljodLpiOpGRLDZY8ofeTjub
SiaTTiacu4O0xrfSWahJ8Wol+MDG5WpB8J4srSaJZrHPfU4iPh2Yde+qhYAl
b2x9us9wRiaPkeXRVR2QvOHe9Od9SHQ3cM8avQ0sNbuQymfoFcgu9kwnKQHu
TE21MlDmudg5/0ieJfF5W28YLUAasuOIgoA5QoSE5a1o8A+WbbSxO6HjnY7k
T447mGWxJLoRj4oCOQSsqwImWOiVuHYgAnb6TyYjGyBbfSyBx/5WBUKvvtxO
ftPYoH70DdOjpVrP+wshpbsWb/rJjq872DlSMIH68kCec8YTBJpSAbzf6vWD
e6PzJvEpcxvZk7t5svBtf6J6hDw3rZ6FVrBOsKlZ0uzQ3RcfApio/RfcjasU
e2rugQ8qASdIpFtFX/GaPjzPSdlonK9QFzV1LstevsG8mun4c0MrxvFeS96a
XL+1Orism+oqLY+ejpAvlkuDOpftQA2ds8greqrQiP57Zyl2PF66lhxW33uW
uKHKdpL7OzepDun42E66+yj5ogIYIIQWNxMnlCpHiuwiFYyoo+VjcPZ7imRL
M7EPHEbewhHwMUHjmX9XQcLAurOmWfsXIALkBHB/KfnhfR30YBNdrIz/SEBN
zs48ZegjbzsRqRRR2j3dkm2umRbyk+aGN6HOML5iM05h43fBPAq7DufXEKu9
k+9RvEiLuhpJoURZgLMq9CXa7I0ltvTE95liAiobydPVIKodk+xYvqPS0WUW
BHvNwH4oJp6b5VJ5ZKLy9FVg+9/5RENMguoZ+EDlJ6LT/UZ/5p0u2UtrpXue
WG36koc0JwRGhfR+lnAXmI/8tM/8OA9V3/vma9Rmf/SRTBU8pL7zZ5PU3ghC
F76olC9I9txozx8IEZETxO5fKE65kpEUOBwGDoOvRYqcun7uriC4I6PDW46p
Q22IdeWALz+wxug+PT0AlqejTqg7b8qZdfg2qfMK0axAjnLjsLHfMtnRsRDb
vrg0FWjS22WsOkuOgoEm9Y2tKeYhpWJ+DbWedW4iUjwU7y+DY380DqbeufNx
BpHqu1MRpQfmqLQmmAl4rUoDvqNJ0Bv/NI+mxQZSclrY0quhGOlr538G2dwQ
Bo+4QR5qIVxYD5n7TXPq8Q/U5T7MqT7kScZQux2qW90zZixlRoP9s/8/IWKi
9SJVhjznbxfnlW4Dg2yneIpJ80AFeaESD3iJpev4IGcppkZnQ6KBYZPJ63hE
as6ewVFZdZJ6A0LfaX+GFnM5Ba3fk2jeoRd8bUgHFxk0d+QpOMeILGbVtDaD
FkMfhEIje1QTp+3AEI20eVYkTbxi9YzfcI3NeHcQbgP63M8nckTLG9/jcfe0
aA7V26/wo8oSjbS9vtDb/HHs1JWUhEz1SgiHtqr+fbtzbv+Lc6SjqJyBZueA
8ygzlKHbckTqX3oUN5uzTPazeOr639Oy8jqM2rJ+TxcomHfB+O8K6fl+nYu8
gDk+mPMdx8+pmb0EIZL5WIfKjwsL5JS0fa6kk76R5aVxX3L8XxkAZ8MwAhBd
ASQhvl72dQZviItGvVmkE8RB2+6XP9fNJwZA0ZyWxEN8uF1V+MW3wHjGGVfg
oDmzrJWjJJpv8AyUi/rupUwtgLdjfyC/suq1uIFuAVWG28c/iziWMXWawcZ0
yQSryCmdLnpQ/LUKcLg8DJkaKI0dQk+Wea2S7SiYFXhRWGZ5ty7C90M0ygh+
jLthH4KdGcUiYifJSDhyIQF1OnA6wCp91l6MewP2UhkwFknCNhRPlp4Cml70
AqBnV5tVO9fk+ohUJNKjXuDEKSMsKm2BsZVm8UeY+lW9FelB6YvOCafj8B0+
MHPCd++aJKmI/cs4sa9tj3y5LSmcDR8S7F5B7kM9b6gHdgGKVv1s5GHWvin+
Ns97Xi3Ybss0+d7B4IxJ6R6Go/AYuLhsZFDpnx6I6LZqIPEv9IzppvzZNpii
iaBYS6xJCGEFvmH0PGSuFNobEAiTO4HB9H/crhax2RiG72XbBPNZgTqmK6VE
zJxnVJUG2ivQr/IxVngN0Q20kZD/VZSWFFrj1z+q3JhW0yCrWiLi1PcZ/2/r
Bsfhbqjg3Z3zxJPMC2hFVxPBwYg13Tde+f6+Knqh7WN6JpQawd7ZS6iNRgzq
+0v/k4E03NzJcPQRuu9D+hFCCSNz7RCF+aqX2mgBEy9d/lsUr2L3uws6VC8d
2MH+Eut9ND/dyvs75cN3eo22vYQQq9PGaGmkIGpZNYgv6ITcqRLFloFgh7iV
J46t0uE6l34YvhbgKoOvwvybsXkudA9w3tUy+fbHDZyP7eVva9vZcKJ1vRZl
2C8H7aOI95w91uFIiHQ5cCLRorh8b5tdq/6JxFIb4rH1pd/SeQWPVktpGSLj
MX3Tm9wvpixRGFXIAZs2B72p1BTbjn4umdq/r1YcoqdpEvNBWCNNjSG901kJ
EfBnpLV/sAHlBGkfmuv5MVceMEOsOohKBq/4iF6KsgyJFwk70cCQE+x+KwDl
ca1GXpK7zFsbZ8cu0Aslij9/WBiQhLus7Z2wETQrDWR6l1BCjjWuogQnlqVv
WxXoZPK19J7PdMC4vlIA+bZg8COXvXcawI6iXaA/WWk5oFRdS/wTcd8lfGam
+pw9IrNkcX/6STPFMzs+67dFGJy62IhM1pB1efRYZox8AHC/UeeGmaxXCCYx
MK5pS5Es6M3AYCEl2XEAu/BRq+kfVGjQ7GY9NKAavEuCptojSEhwMLh2LKnx
957d4ihBT5DtG16vtFhNQa0Yw2qQrZ+V0STwYD6rcZkOTKV/tQo5eMbq7eCE
WHwP3g9G8NkcPiBQLsMNjSWU4/3Q+cOjdxId2//bqZmjJtW8cNIgeBRn+0aB
tJiGuNqHyia+9OmmVaguH9jblfzErj1mzqaGoJ8givkiTvMvP4Ad59/LRM2n
6Tk1dBJEOmy3rMjlEivqYJVXxMT/+rnedpeqRkun5j0OkxtC964seruYRcwq
W4bazt0/ywNMVkrW9emzGApXF/aFh8lYnPDqtpSMJo8UtXG0xs0P7prUodWh
XmbMeQDSBdf6D2IuId/PCIGcmJTrbhFnBwGW21rYVHYlkDzSx2zNW2hpRdv3
JkZkH9c4usOzWR0UIGBJjmpuBynWnWEuP3LCBn++Nq75iFVqG0T9431+P2sH
DysUV2zzxXsXQk7wA/gUzCIJhDj6EDE9aPgrPg78cpO5c3uF+4uLUfNBFDBy
LhOoAqWYzvTyO4ZU7RHAjsaIf9zTbIXaT3DYH1ALSxOSQG+YwoSEfggtanlH
iFMSdajkHVT9y2g/9iflckoMlQU4Ws+CvA8PJLhPAXtoaloTZc/X9RYM7sJW
osUcjrr2+bU4MCj6YufXiG6DLJIVCLMPJRm2NLncFrVYHsV9P1TtNhROMi9k
3qC/8+u54mIy/cWJ8jCyc/azV5nk/0Gqyh8qt/l/epbW1Gg2XMrLJFrMIx+g
tzTY8fiLhc2f4fpKIFmiBoeubEh++bvc7N639MgTF5Y0pT66VzRQmMaxoSd1
fOfrkYv8XWaQH1bCA06VQNwcJLK205vGH/iStTqBS1ExOM2vWBSjJBdMnLhP
hzgb+nTSF/jIE/v8nP+WV4AjpBqjB+khAFso4OadltJ5MQcHbhfZNcEz/beO
Rg072psSnAFpHfyTwNfVjvmjMHO1k3W1bpHuAg/uDhPnTbHibjYRoOUNgkX3
33JauVsxwS3CfaFybfJ4Co1VobLH2Cf1aPL5dVAUipbF+nanclVG4DGdUObD
MMII3TZP008k3/tXSwYhtyG/RmakGGzOLV4sBkzaCg/FVyJs+e9D/62SIdyy
/Vd7B649/P3Qz45I6HH4T2lCC20z5uQoGPlKyfkndCSAXjJtTyZpKXv5g13U
e7dq9bVjGDQLYX9ODk86jrITGwm1VV7GT8UJzov5PehhhB4b9rEcccXC14XS
VCouX4lDTl59EOeqc209ivg13V24wB6xrKynGjMd9Valwg8lHUtqvgGORKl5
+EMQEIcmw3JBOVgZM0cCkSP9IL1S/cgqH8Yv/R4RWKV6KsrNsvqxmOS37yu5
D1a29I2hOOE5JvJnFJIRBRPIjgXiWnU7mj7rk2F79UrEGnjjWAS5KsMOcOJY
tCtMBJ/qqL9b3JfWedDKjB2/Jl9rA2mlxPb1DwIdrBScdip/X+wF+bR0dy/N
NrwENjfyG+TmytoC18zF0c1zjBE6/oX8x5+BWPUh3qZeyJkze37A5zHRDtKx
MtesKucwookb9K+bCvOH+IUi56cAzG2WK1K3WzmCmKTaPrX/91K1WzMZ4D4S
IcJtLhp/wVo9QwhVx26HIvnUw8nUHcthkcvlSGxJPZ677cJi37dAs7BMUIXr
3m6UWwIC+/Dt6DR5RvMCkgHAoRFpCopYjhjlONMaroyqrov9m3Hhgb/hcueg
4vOIdCR3RjduzTT6kBK8nJi01UDy0GniIdKFTc4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG1akfpi3jIN3UjXvG6B2TvF1Yi2jRexRYI2vGTcXAC7E98BChMvGKUQn58pSGPhV1uNpeGohP17B9DKNw+JbwvtFK/1gk1Sq4Vzo3dwePp3sX+xkbGkkHgqqSDTTVWvJToUGYG2GXxdluruP0dkXw33t13H1xsQbOLA5PU0LyoRFK099GiK4a0PyzAbnE7Y90kpK3V/6nrmXhad397YFSiliCtYmEpaGiqG/6Av00IriZcE0gFH15QAS+hFcLspTliIm3Sd7Y091RHYwQF3ws5FPg2arPMBcQSDdHfvw9j1n7SMHL2zbfJcUHK5PtfF6b6+yUHXb2UjiJJdsLNoGMmb+NceFv2mD9itYyv2YQigppdB9H9e+kiE96nrxR/4UYmsTqTTQutIB+SLOhvV6YMTlhlbeOYF7hAFmRZxoolsQpVA0hl23mpKhuwyAQIrtzBWYsFRyDIavLd+U1Flo2snabnxzEr3Rlkmauor1byJtiEXDOKwsmsLlNnTNfFibu8xTCkCdFry9a7r5MAxKR3VEJIM6bpgpp6zCy20Bvz65LyFAX4QuDsQg5W+3BrH+qdLrrj4U47L+XFjARMH3nRp7kfnZwnnAiW0YZbARRq/zDje1I9EQ4ymiKa+l3pw77jmpRezmkit4Pfm1iVC9UMsYXOeK1WniDinOSC7xi+PKXRWHM9LQSe6o04QKigXc7BHAAMGQk76GD2OoATAXoEc7ZexX4sUS0iJEe0cMzkqoUdG+7YdNt0nJ0Py8Ul1uRujnXAX1XSmvBb7p3fAVCLE"
`endif