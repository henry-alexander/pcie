// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q0tTvZYzcP87bWaIuH4+LLJZlzrzO62WW/cU4OZOQ94c4xei3bWYg9Tp22ek
lZJJaNimnykYdGe/DCQO2FPThJyW8RMo8z9v3+jXgpfI1CVhQ3NGTEcr7jrA
O2zC11ywfU6tHvQ7y9QOBxF4ILqTX3tG9JpDzuqDuvgWMtfibN4sKItanu+X
ipXc4X9zM5JzAxFgPVULlWFVFHvgmWg/YDp6Lu5NLjxDmNepVsDjO9IJDFvy
hwVCDGjq/Zn+STyoeT9L4oK2HcuhpoBQCd62se0w6psyRxV5o+7C6jBGkFnX
xymG5TvNQ4SWnecNIsDBclJyj54rabh7PtRqiBHdcA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E1hqFQR+7EC3AFVqsmYeu0WZUrF2+xogY+XmGwu8MWNFd/cDsnBXgbob//fh
SXBg5KoKKAOTwnCIXqaJbdMW6871IlcpxkIHVMPMPg/uGcuWAu+dz0Ip4Fru
Sy2c80QjEyXgN4eDYjE+w+Aucbo1Ia5ZLhfYG9STiTHh/Y0tmc2TDirkZUoV
7YYnTcd3CF+7Wr01YxoR6zRd5ULZxEFGSOS8hCBASmc85js7vCn5agDumc2V
eVPbzPdWrGF1SSiGd8haO1DYXmYsJZokdgo97RHZ3Erfke2KH093dBJsKEY2
uTJWEVxPwL/p0khidZSzzxTZbGy7AHB26GTz/XB/OQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gUED9NpCE4DkQk4PrXaSVcC4Fl+LpF0SgmXf7WSI/H3q+GCDJ5Ko8Rm6wfww
eLhuYTu02JII5jI4rp1Ch68QgcTU7NHhfBdwvmLCaD1+b0OL8GR7HQRHN2uw
xVGthwn9d68yQ3hxssCiWd3spMOR9C6AQyiA5s6T6+6S/VblhvXknGBrDbcL
eiZw6IKq/dpX1dV1gaEBIKsV6rdNBOYHOeFrOEOQvyJL/MpUpwkYFI1+0jns
if5xxa1SzLiQsBkob4k6TJPe40u4Hi8SWd4bGFh+WxA7hciSOXh9T/lw68ee
eEfkN6D+59Xb/obIChOGxxTy7ELHNnj4WUBqYa2U3g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jrPCMc1uD48j+zZ2sJzFjgnMjBkxfnpyb3DyMvdg7dd11oAsdbXSxn9koK3z
c3Y+pKfHTsfMBFrqMuGaHhityU8Rvq8Einh+mNFsfxysBBf6a4EBF0UIasPW
O+Moqf5iPVpzhhyEM8iikTsZ/EWFKI+53iw8d4RcO2cJ+fsdJT4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
jfrYWLTBY58lIjDLm4Wnx6WRDnIL1VKh1MToFmmAoa1Tp2igNgJx/n3Ne25i
8NXYvJ47+54mFn3bxZ3ZBa8W9NQvljgkl7tZemu73SgzZBNLmAOWZZ9I6L9Z
S9E5K3DcjyMOl3Ctpjx0Cd7Kwn71kZ+hV8gzV+pguNHqDmGk2ysyVZ/Ts9x9
JZfKQjtrfzOSv5ubsRrQLYeMPBcwzcX8pLHnPsHre15pVYVG8I8Fpcxbthup
TU9aqrJcWAQkYCT1Bd1wsZKu3HNqI/ayBJM4cWWE97sSW/rg5B0cs5hzyv4n
P8vplsN5Y2ACloOvdjlal2M5nxvhCe7Ubk9R5GZZTmzba+xvD+NT/B5x3gS6
9rdjSI28AuZJ9VpkzEv45xCM6K5lbL0NldKXc8hV2B3eMVzB7G7QmLvkhpuC
YB3Q73UCpPSt3IkIgxB6Rj2bZB33WixVswHMj7Y2qT0OvCj1hPB3JWaDL3Os
AOo+bajIBnnB6VnMyy0KhxaHwPpN0zjP


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
t3g2VDVU7d+Hyfu6yhaTMmxfj9UVjCiEN7ZoUFQ6mggIzDeA1de5yAv856OL
Enre4l7GEUMSvDXYFY2JeaB4SoXnKwOVJ9MV/DAulSJoqVZ29rpRha0v5R1b
fCHazbFkSWUaFnw0+7sW4C8JfzXgfW+oH25G24BMyd0hQMY1mdk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WsdiEPLfkfJsFr3LTPJJRlGqKRaWKStNqhVqK5d6t2qckPH+1aFHqbXUt4GB
D53axerOSQYiNbA25RLkYCj/aHLhia1exsmnTTkbM42dKzXsbQrh0ZQT84DR
A0ZlU5mBcBMUvgnb0ichKYskIKrAYaV5oFhD09g+YyNV2gT643c=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4064)
`pragma protect data_block
/3k5J7tMNr0eqgvUhZ2mMdmMeysld5wlLk/hx0UgACFpOGARIkmuRWbxWpW2
yv0dkoiEKl64vPr3CMmlFppGvbKB5PVF1i0q3outXvTUacXNZAShsQPcUEpj
sRHfTntXCne/RfTX64uRfCw3+4yxwyorEbVQqK9fglZ4YH+iELp4BEb3pTES
yzAYg8kk/u+bB97HlncffJxjb9A7Ae18gufp+1pi04JFq7S6NJojE2/mHC2q
vmCBy0e/W+CKJ+8CdC16dZ13R/DAVWP5UR1/7EpYFSHBzFg6i41vFQu22aJh
QUSzyPuGCs67kSd2rsPxqW6ph0aRrlTOEAOTKhvbeHcO4wnC7yeQx5nGd4sX
riXCLrU/+oy1QSzGZJhCzvuIQ1i9vfzQnpTubNPatF0qgWP7QrJaOLO+46FS
JfcpqRBn1IFivxcW7TW25ID9QX5w7GhZc6/m8tjOR5n49ao9HXtRx2aFPUPU
X5mPlBwU5vZLfMXszwdCKxkQrOruOyV17TfhKI1UTecnwhLt97y3+LvWmxDM
3GKIe0xh7J3akL9cphxo7R4ZWXK0Tr48WuuwZI4JwJxb9UiHA2krQT2A545+
euYQc1Qd2P/dCCBWaRNk5CsO+gdViFskdQpfCfh50/YCExsdAf+0q3OSHxIy
Qpg6hhncYedNFgGWvjRSOGETqdfADvLCoVkb/nXc7SkP6Sm6Uh4XW9Jlky21
WpX68g0kuvKC9NibFlKloHgfe/yzuI6Qc3MEM7RkI74EVNtuXBt9AvqmRxPg
qTxfG5BD5zvBk78pE6T6/p1F3ArgHKXNuMBHbUi/Ii4h1wJm5DsKmXfqSgEM
AzMyr2vZh/63J9u5xtsp2QFnzVIJlb2ObbOMhfzVExIdQbfTpID4qGbLdDU9
hACrTq4o1ec0DbC28TBJRezQ5oSUtXTfBIClzG7Qt93AKfv2xVG8oG3wAYEO
+zFNmtPl5K54ECoXDDoB1lVs7tMoV1TlTjOe6DwsvmXjvszR4TRXy9DcsohU
6cZNltq95ja+KShOjWQIGA57dd8CpdkxGOI/0hV5o45iG7Fq+1+rMYOruwkz
vU+/tD8nbuspbQb4/l/mfJtKdyXsk9lmjZjeqjfp5OJSwAcxJjRSLL/ZJkMD
y4skOfVwv4FEB9y7oCEQgPNBYHEv9W6Ljo4Z9nadUXReM/hQb9rBnRrDaF/2
qc4S4BgU0o9zztkDBtNha2GcPMuGUUKI351a3MTLRmCL+rtDq9mvsOBKHCGr
OwU6SRei2p2Xb1XVmF8AciK2qhDLMO2BIXXXcsa8aEdxF5LFzP3XS1X3+241
YelXmrhLBLPDjou/aTJB6LNpH/WBpxyqx1B5RxiVI5HPfEgm3TC0Rkf9Ui6h
8VIJaMnd/ttb0WVtK8QLIIIAsjanXnqYecMTiTI4SSDxP+5NgaIfFRBiAeQN
9TmYkYnkvzMb1Sh4h8h4AiODNLyq8EIWu6p8vhbLTsP7xqzoFdtt7nQAW3b/
4hf74+jzdD5jMfSl6+pqFiD6y4oIlbdB2jHobEgjrAvsKki2smjoIHICiBKi
QE1PPrqD7Wq/xdk1zGbvxcu27+3GuTkoHVkqPXf0o1ot4Et127eLb5pE2+ak
+bSdxDm64c58bfy9TpMM7nHPmzAcNEPQVqKanGFdvFVJNkJvIA5Bie+BJZxV
rmX9NTf/XmtfWawPNN6XnTqHbBI+B2kBNVczd0ev6Wanru1mNdQ+phLrfe++
xAdY/S4cgLKPX3WO7INX63BMO2f+zf13cfxneiwaZ9tGsaoOYha90MW1Tq+Z
L9ehh10mtfwODxESjOuI0fztALDZMvXhLUtRwIQ5ofqeK5N75yMblU+MlCCE
vS17ykAGiL50TrPHzROkadOLt+Kpt1iXbu3X+jpZXxIHPOLBZ7pzc62l/HqN
IfFiTFnF1PDlCA/MX+/S96kEdxFvYeLxjYR87ywNJXbKpHANrEIGuQRAiBZD
ZiC5d15//wjiYz0HFIih4MrwzIgYMhyXMwu3LzuWVT4G715810HXjv5fKrcJ
FTWrsDaMFqM+C2oVXG/tTsZjdgfAvdFJpchtz7WYbJbxdd6yG5b3rjFbDFw2
8nHhMcAOT64x0GhfxVSBzdwc/8MRVEA3V3xPzQzoEe6g8ndXhJmPlKctjhYb
B1+Vh/zyUoTvxxqWn8JtQ8N+TutejqcbGxqZ/i+uwfxy8FUdD0kpkZ2N+6o+
ny5isgtu5ozFtZ49ahN3WHpNISiOmGL5SaBJGJFOvZ7ZeNm04qyz4hppUOok
e2CXO6e3NuN48dY7PnAmYcqzLznSzx1X+6S7vcGtIQS8dtSUyy/5ArVcEFI0
8fZGasgIAyWearSx9v5HYEUvy/4eeLmROj+cPPr99yxODpg7SM7VKb9SlY95
f+ev//SplPhK3k9YCwgSEPAwN/7nXDCpsuLGGFidMBVM8a8eiohj57QP96Gj
+M7k6O1oh2WkCXwcbBTVMowuh/DX5LA6KHjJiVBwOu6QX03crdYVZ9lqXz4M
BhQeOO4oQbLvrhztzQPmdW+QhvReqqq8CxtSe11RtbiTwjdBgeUJrxZLMv1w
qiqE/vFuN/XrgRDxkZbRg2zuzZaZbJVhqzJ03slzYsYDrq30CKBNWg3xcxU2
GY6n15xixBleWFt8ZmA9sce6lEKa8jV2OTUE93VFloWedg19WpQccMV9sCIy
1NhOKRAVqxfpTCRMwsew2fdSCvDdJuid0czWyMZ9f4mxJ1+rnNcPGvVk/CaM
9g6/8faDKdhFHnSkJOMNajpDAOCEQc6dDAYtQkcuAJ2L1sgVefP54YLp13dj
upWosAuInEYR/Qe+ai1MJ+0UKANrJDGw8TREg4l/NQfSP6/ehNHY5mAUXCCA
IwRLPExgXuq9I/HYuQKyQct+X+ZZBcal7PYwFyKww9zIYN+fEvVHajQQWaix
ielReBlk1smhmtv99WxQg1u8p9QS5mAZx94Enc8YKZJdDTHxqvg1G/lDXxEE
R9UzF35Che3b6+a2zKS6vwqVgl+Ft1V/GQhzRG6CmyDvPsqpMsIrvknCq+0p
Gj+53FZDlUn97HHPbUPu6YqfzH4cvyyNA8a4zIe7ylTjhTgqpBhyuIX5i75O
NJGJSy8Iw0ToWA3n7Hrdv/giUbc/w0l2xe+WYahOvnQqqwxWc2rq4HkmQUaS
Mi9CI7UiHHuQCdVclTHCcpWtXrZDwEXpov2bLdS1Q0L4WDXVsWjS1NjBrHKr
VykFLpRNvk7elR468q9TKAXnuqkGsOplg6KI8g+ZkGgdhwAPAPSYLyZ1wMQS
2i1f4vXPU8wgHHyV1Jet4XxVe5CpoJcshaVnfl0PXcReUMjGtr4siG5WmmnB
or5XDrml/CKjX3D7sWg5q33irA8Z35iydvenPZqhsREuds9THqK0PDTZTPmC
OTa4OwYxj5jQGXwY9AJtilQuhh/iCPB8/l04dOXHq/6YRcIFUFG95Nqwk8mF
hgbS83leB4FEwZVH+yaUDjt4/g9b/CGIcHunipMUtmhY/5dXkWHHgFhTuq97
pTKQx3n82KcFzFA+NdugxAW6SWbEMIKEpLRRZ4perUwUxy2lofbt7QjVB6jy
ZiAMsg7Y97Kz7c9Q4lA5gp2YR+holV/ztXPPEfFK49Zrl+9JWUA9L0RYZPYe
iFOFxobPYdd4r5dN87xhd8Tva6uiGZRnejbuFDUI7zmo6sRM0Gqa1Cu4t1NY
egphQ+MPnyz4zc6cvM3G4oTLNXb5BjvC8DmQHydMd+sm3jNUypFUkT50rPoZ
CA5ZBwHFmP6MKMxPZgZ18zisevhju7jGOUP49ofr+UB5pkrPrES4w8CXKwCM
ck/JSXtQne3ONyvpp/N68TW2y9m5EeeHDFNjvvQGj0T9kjYXhV7AeZVdXMVM
YJsXDqQ0IJ65vyA4tNWICDKm8TqoqkBZRF95NOxY5X9qfuizuUEmxxicSeOU
SYU+BpDlaaG2tEKLMaUAs2yCGpglVKTCcyJG5EF1FtSMrjLaOZMHUoir1dY0
NPekZuUoWNe7EsNWQIdNbD5zUwLq2XzmKt5+v/n8H0eBhvX7PSSn9f54BF2P
WCfzNJimYGO5n7KHfQaub7bSB7hV2VCFKijvNm6/zbKpgJz94+lbbskpKLNL
IqujhJoUfIrrJPpaIp/nNBtryu2E3TbhnBFS5DrocbwD3cH4R/VmOGbfxRtg
5fsqHTVMv/y1dT0q6dPq/znhsBIE93qRspuMwTfrW5HWdgMs/LDDybkXr2Ww
fYQL07NNfgUuRNbCJUQjJrPeYYDlQAucm6FoEfLqpC8f5aMimcC0VGgDHQyO
4BKqo6LoVqZUEPAfELpM8UUpp2O2CTXYZEFpaKwJBaHozks2T6MI5RMjNjMs
oS1LXEzBn7lBMXHdYHD8PvW85JDI4gailVT1Mr0G7aXUxxD7Cgr1RfoSDb/n
a5iWh3RmsD/u15l5mI792b9728+cihGczeiXygaTqo/n/M601hHi3IH0gpa2
c4swFffcpf+VHIdCe0YbmCmv0FQYSjibDSFkVQVvaNQB4o5YNFPYjZY60/i+
NXYUST23vn3fnhvVjaAVu08C/6FarHU+k5SO/clCgkukgZGwGShLDi7TGLsL
FOrgtIQyooNJJu4KvI6rBx3EA4m+/JrTyTCCBaZ0sQD1npXXcJ+Ioyi7W+z9
5H+q7YOZGOAVfRVXOzSLCcqxfkbUl6FYnL7zpWBU9ggPwODNq7/gD8Sj1slx
xjWqmerDAnz+9YrEjUSP4rSEt8RCuJlLzCIlh3UJPdl9yl38I/xYZlTpDjAa
IIzg30JF353JIhGl1+9lkCfGt6uaAzm06qDsEm2Hom7Y3k1JwGdbmESfkhVj
byKFnlQVOrqXNZheKR3+/9amvkeCR0eUx1HIHaZaiX+zKUoTyTepanO1q7o9
SXfiR4uojfuQ7ZeR/DCOVAmKu2+8z/LM+w93W9edlYbKzDhgrEn+lNV4h8jt
e8i6M/NlP+LWcKI7nT2/LwCtzT/A1QWx99M6Ui4Zj2S0MXuLBl0AWLzVy7Ix
lxMU5Rqcsf/SEj43bfhU3TctUWI6JOkZW+3B6on1Kg8kkgZ0A5X8JdksOV6N
n+qXvq+wc89s+Exk6Se0QZoOCiTYFLuoOJRoFHbWPuBWj8kudyQQVZKapFhq
c5Auxqq+X77lrNRGFmkWv1adEeZlSy/OK0/y4gb3w3bCWW5ErNEUqd96HpQ9
R/1pGY6vuW/JW65552um8+vLOWONA/qZpbce1sdvBXyDCmSgmT3zLApZDqAU
dVUxaIko9prao++HstWygrVPvh1ja9+l1DNbUAYUwpUz+qMDAnUZJ7sDXMG0
1/rSKbn/GDHhlUFDETruphUjlkHliMcEAasDsndGqRy/BPdgAoj/0Mb+/Pos
LQA0Shb1FKRpThfKdOE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfSiY76SUVoesnBkCLLTal50kGafTUzBCkckSunwTBwc+r4MOQ6848dX1qVwkoTDZSLGBYtad1vjiuYYUW5SBtdzvW1ZHfM6Vs0OoQTzM/LCRc66LXkhKfNRLAr+qZ8F/LeSINcXG1ncRVkUVW1opdo+N12jU6LFntveP7oCLEpgBYLJF+YJErRlZaHf4urDDhiy6gUT95AkTdy+kEZQapg9f9BNeOX9jUxyMzVghjBPs63WuA5AhhhIXN/DDM3Fq3hPmoaau03+OL1phFH7Y+01maXUXp4Fi2f/Thm3UUbS5LB/9Z96F5gKu6/AvpnK1o+fL3HS8fpJGDmMA82RarJROfiX/Ls7xVhDmBgssbqmCe8cqD8zgzF7LdKnnSMc6fiQdR4EVQ8bxpfyy2hVQCTi/gDZfeSUBO8YSDI10ORJsZJBs4EgM6W+e3gaBGRxHQkC+xMCczqwuqNNwYfmyPwxjELjQXSIgIgrkbEly8BhSII9h9Jt+xyhb8qGY25g9JKNq6WOOTfZNZlFPJG/bGQzHmkIqeWMDKD7bljFOFZwsmtFlSTO11jyyLK3d1+dSxCLfsHxwpsuE1LiHtFF+TP91127CqksIqbs3zqNxgykGNBrmYwoMKOGw/ZuesvvPNwjem1u2gbHHatg8JMSUJxsdkG8Gr1ZGSkbaW9sf+ooib5WdHaylm3m4O8teBdorV+KWF5YzURH98r98q8N8xNysAI1ni9bilkIznWck8QFpAOdQiw4Uzu0R+4MheGYoBeeIcxJUsyZeLjLq3O5LsxC"
`endif