// system_intel_pcie_gts_0_pcie_hal_top_pipe_hal_2100_e6uglya.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_intel_pcie_gts_0_pcie_hal_top_pipe_hal_2100_e6uglya #(
		parameter       sris_enable   = "SRIS_ENABLE_DISABLED",
		parameter       pcie_pcs_mode = "PCIE_PCS_MODE_PCIE",
		parameter[31:0] pclk_clk_hz   = 32'b00111011100110101100101000000000,
		parameter       num_of_lanes  = 4
	) (
		input  wire [16:0] i_ch0_lavmm_pcie_addr,                          // pipe_hal.i_ch0_lavmm_pcie_addr,                          Check User Guide for details
		input  wire [3:0]  i_ch0_lavmm_pcie_be,                            //         .i_ch0_lavmm_pcie_be,                            Check User Guide for details
		input  wire        i_ch0_lavmm_pcie_clk,                           //         .i_ch0_lavmm_pcie_clk,                           Check User Guide for details
		input  wire        i_ch0_lavmm_pcie_read,                          //         .i_ch0_lavmm_pcie_read,                          Check User Guide for details
		input  wire        i_ch0_lavmm_pcie_rstn,                          //         .i_ch0_lavmm_pcie_rstn,                          Check User Guide for details
		input  wire [31:0] i_ch0_lavmm_pcie_wdata,                         //         .i_ch0_lavmm_pcie_wdata,                         Check User Guide for details
		input  wire        i_ch0_lavmm_pcie_write,                         //         .i_ch0_lavmm_pcie_write,                         Check User Guide for details
		input  wire        i_ch0_pcie_rxword_clk,                          //         .i_ch0_pcie_rxword_clk,                          Check User Guide for details
		input  wire        i_ch0_pcie_txword_clk,                          //         .i_ch0_pcie_txword_clk,                          Check User Guide for details
		input  wire        i_ch0_pcs_pclk,                                 //         .i_ch0_pcs_pclk,                                 Check User Guide for details
		input  wire        i_ch0_pcs_pipe_rstn,                            //         .i_ch0_pcs_pipe_rstn,                            Check User Guide for details
		input  wire        i_ch0_txpipe_asyncpowerchangeack,               //         .i_ch0_txpipe_asyncpowerchangeack,               Check User Guide for details
		input  wire        i_ch0_txpipe_blockaligncontrol,                 //         .i_ch0_txpipe_blockaligncontrol,                 Check User Guide for details
		input  wire        i_ch0_txpipe_cfg_hw_auto_sp_dis,                //         .i_ch0_txpipe_cfg_hw_auto_sp_dis,                Check User Guide for details
		input  wire        i_ch0_txpipe_dirchange,                         //         .i_ch0_txpipe_dirchange,                         Check User Guide for details
		input  wire        i_ch0_txpipe_ebuf_mode,                         //         .i_ch0_txpipe_ebuf_mode,                         Check User Guide for details
		input  wire        i_ch0_txpipe_encodedecodebypass,                //         .i_ch0_txpipe_encodedecodebypass,                Check User Guide for details
		input  wire [5:0]  i_ch0_txpipe_fs,                                //         .i_ch0_txpipe_fs,                                Check User Guide for details
		input  wire        i_ch0_txpipe_getlocalpresetcoefficients,        //         .i_ch0_txpipe_getlocalpresetcoefficients,        Check User Guide for details
		input  wire        i_ch0_txpipe_invalidrequest,                    //         .i_ch0_txpipe_invalidrequest,                    Check User Guide for details
		input  wire [5:0]  i_ch0_txpipe_lf,                                //         .i_ch0_txpipe_lf,                                Check User Guide for details
		input  wire [4:0]  i_ch0_txpipe_localpresetindex,                  //         .i_ch0_txpipe_localpresetindex,                  Check User Guide for details
		input  wire        i_ch0_txpipe_lowpin_nt,                         //         .i_ch0_txpipe_lowpin_nt,                         Check User Guide for details
		input  wire [7:0]  i_ch0_txpipe_m2p_bus,                           //         .i_ch0_txpipe_m2p_bus,                           Check User Guide for details
		input  wire [2:0]  i_ch0_txpipe_pclk_rate,                         //         .i_ch0_txpipe_pclk_rate,                         Check User Guide for details
		input  wire        i_ch0_txpipe_pclkchangeack,                     //         .i_ch0_txpipe_pclkchangeack,                     Check User Guide for details
		input  wire [3:0]  i_ch0_txpipe_phy_mode_nt,                       //         .i_ch0_txpipe_phy_mode_nt,                       Check User Guide for details
		input  wire [3:0]  i_ch0_txpipe_powerdown,                         //         .i_ch0_txpipe_powerdown,                         Check User Guide for details
		input  wire [2:0]  i_ch0_txpipe_rate,                              //         .i_ch0_txpipe_rate,                              Check User Guide for details
		input  wire        i_ch0_txpipe_rxelecidle_disable_a,              //         .i_ch0_txpipe_rxelecidle_disable_a,              Check User Guide for details
		input  wire        i_ch0_txpipe_rxeqclr,                           //         .i_ch0_txpipe_rxeqclr,                           Check User Guide for details
		input  wire        i_ch0_txpipe_rxeqeval,                          //         .i_ch0_txpipe_rxeqeval,                          Check User Guide for details
		input  wire        i_ch0_txpipe_rxeqinprogress,                    //         .i_ch0_txpipe_rxeqinprogress,                    Check User Guide for details
		input  wire        i_ch0_txpipe_rxeqtraining,                      //         .i_ch0_txpipe_rxeqtraining,                      Check User Guide for details
		input  wire        i_ch0_txpipe_rxpolarity,                        //         .i_ch0_txpipe_rxpolarity,                        Check User Guide for details
		input  wire [2:0]  i_ch0_txpipe_rxpresethint,                      //         .i_ch0_txpipe_rxpresethint,                      Check User Guide for details
		input  wire        i_ch0_txpipe_rxstandby,                         //         .i_ch0_txpipe_rxstandby,                         Check User Guide for details
		input  wire        i_ch0_txpipe_rxtermination,                     //         .i_ch0_txpipe_rxtermination,                     Check User Guide for details
		input  wire        i_ch0_txpipe_srisenable,                        //         .i_ch0_txpipe_srisenable,                        Check User Guide for details
		input  wire        i_ch0_txpipe_txcmnmode_disable_a,               //         .i_ch0_txpipe_txcmnmode_disable_a,               Check User Guide for details
		input  wire        i_ch0_txpipe_txcompliance,                      //         .i_ch0_txpipe_txcompliance,                      Check User Guide for details
		input  wire [39:0] i_ch0_txpipe_txdata,                            //         .i_ch0_txpipe_txdata,                            Check User Guide for details
		input  wire [3:0]  i_ch0_txpipe_txdatak,                           //         .i_ch0_txpipe_txdatak,                           Check User Guide for details
		input  wire        i_ch0_txpipe_txdatavalid,                       //         .i_ch0_txpipe_txdatavalid,                       Check User Guide for details
		input  wire [17:0] i_ch0_txpipe_txdeemph,                          //         .i_ch0_txpipe_txdeemph,                          Check User Guide for details
		input  wire        i_ch0_txpipe_txdtctrx_lb,                       //         .i_ch0_txpipe_txdtctrx_lb,                       Check User Guide for details
		input  wire        i_ch0_txpipe_txelecidle,                        //         .i_ch0_txpipe_txelecidle,                        Check User Guide for details
		input  wire [2:0]  i_ch0_txpipe_txmargin,                          //         .i_ch0_txpipe_txmargin,                          Check User Guide for details
		input  wire        i_ch0_txpipe_txoneszeros,                       //         .i_ch0_txpipe_txoneszeros,                       Check User Guide for details
		input  wire        i_ch0_txpipe_txstartblock,                      //         .i_ch0_txpipe_txstartblock,                      Check User Guide for details
		input  wire        i_ch0_txpipe_txswing,                           //         .i_ch0_txpipe_txswing,                           Check User Guide for details
		input  wire [3:0]  i_ch0_txpipe_txsyncheader,                      //         .i_ch0_txpipe_txsyncheader,                      Check User Guide for details
		input  wire [2:0]  i_ch0_txpipe_width,                             //         .i_ch0_txpipe_width,                             Check User Guide for details
		input  wire        i_ch0_uxq_rxcdrlock2dataa,                      //         .i_ch0_uxq_rxcdrlock2dataa,                      Check User Guide for details
		input  wire [13:0] i_ch0_uxq_rxeq_best_eye_vala,                   //         .i_ch0_uxq_rxeq_best_eye_vala,                   Check User Guide for details
		input  wire        i_ch0_uxq_rxeq_donea,                           //         .i_ch0_uxq_rxeq_donea,                           Check User Guide for details
		input  wire        i_ch0_uxq_rxmargin_nacka,                       //         .i_ch0_uxq_rxmargin_nacka,                       Check User Guide for details
		input  wire [1:0]  i_ch0_uxq_rxmargin_status_gray_a,               //         .i_ch0_uxq_rxmargin_status_gray_a,               Check User Guide for details
		input  wire        i_ch0_uxq_rxmargin_statusa,                     //         .i_ch0_uxq_rxmargin_statusa,                     Check User Guide for details
		input  wire        i_ch0_uxq_rxsignaldetect_lfpsa,                 //         .i_ch0_uxq_rxsignaldetect_lfpsa,                 Check User Guide for details
		input  wire        i_ch0_uxq_rxsignaldetecta,                      //         .i_ch0_uxq_rxsignaldetecta,                      Check User Guide for details
		input  wire        i_ch0_uxq_rxstatusa,                            //         .i_ch0_uxq_rxstatusa,                            Check User Guide for details
		input  wire [39:0] i_ch0_uxq_rxword,                               //         .i_ch0_uxq_rxword,                               Check User Guide for details
		input  wire        i_ch0_uxq_synthlcfast_postdiv,                  //         .i_ch0_uxq_synthlcfast_postdiv,                  Check User Guide for details
		input  wire        i_ch0_uxq_synthlcmed_postdiv,                   //         .i_ch0_uxq_synthlcmed_postdiv,                   Check User Guide for details
		input  wire        i_ch0_uxq_synthlcslow_postdiv,                  //         .i_ch0_uxq_synthlcslow_postdiv,                  Check User Guide for details
		input  wire        i_ch0_uxq_txdetectrx_acka,                      //         .i_ch0_uxq_txdetectrx_acka,                      Check User Guide for details
		input  wire        i_ch0_uxq_txdetectrx_statct,                    //         .i_ch0_uxq_txdetectrx_statct,                    Check User Guide for details
		input  wire        i_ch0_uxq_txstatusa,                            //         .i_ch0_uxq_txstatusa,                            Check User Guide for details
		output wire [31:0] o_ch0_lavmm_pcie_rdata,                         //         .o_ch0_lavmm_pcie_rdata,                         Check User Guide for details
		output wire        o_ch0_lavmm_pcie_rdata_valid,                   //         .o_ch0_lavmm_pcie_rdata_valid,                   Check User Guide for details
		output wire        o_ch0_lavmm_pcie_waitreq,                       //         .o_ch0_lavmm_pcie_waitreq,                       Check User Guide for details
		output wire        o_ch0_pcs_pclk,                                 //         .o_ch0_pcs_pclk,                                 Check User Guide for details
		output wire        o_ch0_pcs_pipe_rstn,                            //         .o_ch0_pcs_pipe_rstn,                            Check User Guide for details
		output wire [5:0]  o_ch0_rxpipe_dirfeedback,                       //         .o_ch0_rxpipe_dirfeedback,                       Check User Guide for details
		output wire [7:0]  o_ch0_rxpipe_linkevaluationfeedbackfiguremerit, //         .o_ch0_rxpipe_linkevaluationfeedbackfiguremerit, Check User Guide for details
		output wire [5:0]  o_ch0_rxpipe_localfs,                           //         .o_ch0_rxpipe_localfs,                           Check User Guide for details
		output wire [5:0]  o_ch0_rxpipe_locallf,                           //         .o_ch0_rxpipe_locallf,                           Check User Guide for details
		output wire        o_ch0_rxpipe_localtxcoefficientsvalid,          //         .o_ch0_rxpipe_localtxcoefficientsvalid,          Check User Guide for details
		output wire [17:0] o_ch0_rxpipe_localtxpresetcoefficients,         //         .o_ch0_rxpipe_localtxpresetcoefficients,         Check User Guide for details
		output wire [7:0]  o_ch0_rxpipe_p2m_bus,                           //         .o_ch0_rxpipe_p2m_bus,                           Check User Guide for details
		output wire        o_ch0_rxpipe_pclkchangeok,                      //         .o_ch0_rxpipe_pclkchangeok,                      Check User Guide for details
		output wire        o_ch0_rxpipe_phystatus,                         //         .o_ch0_rxpipe_phystatus,                         Check User Guide for details
		output wire [39:0] o_ch0_rxpipe_rxdata,                            //         .o_ch0_rxpipe_rxdata,                            Check User Guide for details
		output wire [3:0]  o_ch0_rxpipe_rxdatak,                           //         .o_ch0_rxpipe_rxdatak,                           Check User Guide for details
		output wire        o_ch0_rxpipe_rxdatavalid,                       //         .o_ch0_rxpipe_rxdatavalid,                       Check User Guide for details
		output wire        o_ch0_rxpipe_rxelecidlea,                       //         .o_ch0_rxpipe_rxelecidlea,                       Check User Guide for details
		output wire        o_ch0_rxpipe_rxstandbystatus,                   //         .o_ch0_rxpipe_rxstandbystatus,                   Check User Guide for details
		output wire        o_ch0_rxpipe_rxstartblock,                      //         .o_ch0_rxpipe_rxstartblock,                      Check User Guide for details
		output wire [2:0]  o_ch0_rxpipe_rxstatus,                          //         .o_ch0_rxpipe_rxstatus,                          Check User Guide for details
		output wire [3:0]  o_ch0_rxpipe_rxsyncheader,                      //         .o_ch0_rxpipe_rxsyncheader,                      Check User Guide for details
		output wire        o_ch0_rxpipe_rxvalid,                           //         .o_ch0_rxpipe_rxvalid,                           Check User Guide for details
		output wire        o_ch0_ux_ock_pma_clk,                           //         .o_ch0_ux_ock_pma_clk,                           Check User Guide for details
		output wire        o_ch0_uxq_lfps_ennt,                            //         .o_ch0_uxq_lfps_ennt,                            Check User Guide for details
		output wire [1:0]  o_ch0_uxq_pcie_l1ctrla,                         //         .o_ch0_uxq_pcie_l1ctrla,                         Check User Guide for details
		output wire        o_ch0_uxq_pma_cmn_ctrl,                         //         .o_ch0_uxq_pma_cmn_ctrl,                         Check User Guide for details
		output wire        o_ch0_uxq_pma_ctrl,                             //         .o_ch0_uxq_pma_ctrl,                             Check User Guide for details
		output wire        o_ch0_uxq_rst_pcs_rx_b_a,                       //         .o_ch0_uxq_rst_pcs_rx_b_a,                       Check User Guide for details
		output wire        o_ch0_uxq_rst_pcs_tx_b_a,                       //         .o_ch0_uxq_rst_pcs_tx_b_a,                       Check User Guide for details
		output wire        o_ch0_uxq_rxeiosdetectstata,                    //         .o_ch0_uxq_rxeiosdetectstata,                    Check User Guide for details
		output wire [2:0]  o_ch0_uxq_rxeq_precal_code_selnt,               //         .o_ch0_uxq_rxeq_precal_code_selnt,               Check User Guide for details
		output wire        o_ch0_uxq_rxeq_starta,                          //         .o_ch0_uxq_rxeq_starta,                          Check User Guide for details
		output wire        o_ch0_uxq_rxeq_static_ena,                      //         .o_ch0_uxq_rxeq_static_ena,                      Check User Guide for details
		output wire        o_ch0_uxq_rxmargin_direction_nt,                //         .o_ch0_uxq_rxmargin_direction_nt,                Check User Guide for details
		output wire        o_ch0_uxq_rxmargin_mode_nt,                     //         .o_ch0_uxq_rxmargin_mode_nt,                     Check User Guide for details
		output wire        o_ch0_uxq_rxmargin_offset_change_a,             //         .o_ch0_uxq_rxmargin_offset_change_a,             Check User Guide for details
		output wire [6:0]  o_ch0_uxq_rxmargin_offset_nt,                   //         .o_ch0_uxq_rxmargin_offset_nt,                   Check User Guide for details
		output wire        o_ch0_uxq_rxmargin_start_a,                     //         .o_ch0_uxq_rxmargin_start_a,                     Check User Guide for details
		output wire [2:0]  o_ch0_uxq_rxpstate,                             //         .o_ch0_uxq_rxpstate,                             Check User Guide for details
		output wire [3:0]  o_ch0_uxq_rxrate,                               //         .o_ch0_uxq_rxrate,                               Check User Guide for details
		output wire        o_ch0_uxq_rxterm_hiz_ena,                       //         .o_ch0_uxq_rxterm_hiz_ena,                       Check User Guide for details
		output wire [2:0]  o_ch0_uxq_rxwidth,                              //         .o_ch0_uxq_rxwidth,                              Check User Guide for details
		output wire        o_ch0_uxq_tstbus_lane,                          //         .o_ch0_uxq_tstbus_lane,                          Check User Guide for details
		output wire        o_ch0_uxq_txbeacona,                            //         .o_ch0_uxq_txbeacona,                            Check User Guide for details
		output wire [2:0]  o_ch0_uxq_txclkdivrate,                         //         .o_ch0_uxq_txclkdivrate,                         Check User Guide for details
		output wire        o_ch0_uxq_txdetectrx_reqa,                      //         .o_ch0_uxq_txdetectrx_reqa,                      Check User Guide for details
		output wire [5:0]  o_ch0_uxq_txdrv_levn,                           //         .o_ch0_uxq_txdrv_levn,                           Check User Guide for details
		output wire [4:0]  o_ch0_uxq_txdrv_levnm1,                         //         .o_ch0_uxq_txdrv_levnm1,                         Check User Guide for details
		output wire [2:0]  o_ch0_uxq_txdrv_levnm2,                         //         .o_ch0_uxq_txdrv_levnm2,                         Check User Guide for details
		output wire [4:0]  o_ch0_uxq_txdrv_levnp1,                         //         .o_ch0_uxq_txdrv_levnp1,                         Check User Guide for details
		output wire [3:0]  o_ch0_uxq_txdrv_slew,                           //         .o_ch0_uxq_txdrv_slew,                           Check User Guide for details
		output wire [3:0]  o_ch0_uxq_txelecidle,                           //         .o_ch0_uxq_txelecidle,                           Check User Guide for details
		output wire [2:0]  o_ch0_uxq_txpstate,                             //         .o_ch0_uxq_txpstate,                             Check User Guide for details
		output wire [3:0]  o_ch0_uxq_txrate,                               //         .o_ch0_uxq_txrate,                               Check User Guide for details
		output wire [2:0]  o_ch0_uxq_txwidth,                              //         .o_ch0_uxq_txwidth,                              Check User Guide for details
		output wire [39:0] o_ch0_uxq_txword,                               //         .o_ch0_uxq_txword,                               Check User Guide for details
		input  wire [16:0] i_ch1_lavmm_pcie_addr,                          //         .i_ch1_lavmm_pcie_addr,                          Check User Guide for details
		input  wire [3:0]  i_ch1_lavmm_pcie_be,                            //         .i_ch1_lavmm_pcie_be,                            Check User Guide for details
		input  wire        i_ch1_lavmm_pcie_clk,                           //         .i_ch1_lavmm_pcie_clk,                           Check User Guide for details
		input  wire        i_ch1_lavmm_pcie_read,                          //         .i_ch1_lavmm_pcie_read,                          Check User Guide for details
		input  wire        i_ch1_lavmm_pcie_rstn,                          //         .i_ch1_lavmm_pcie_rstn,                          Check User Guide for details
		input  wire [31:0] i_ch1_lavmm_pcie_wdata,                         //         .i_ch1_lavmm_pcie_wdata,                         Check User Guide for details
		input  wire        i_ch1_lavmm_pcie_write,                         //         .i_ch1_lavmm_pcie_write,                         Check User Guide for details
		input  wire        i_ch1_pcie_rxword_clk,                          //         .i_ch1_pcie_rxword_clk,                          Check User Guide for details
		input  wire        i_ch1_pcie_txword_clk,                          //         .i_ch1_pcie_txword_clk,                          Check User Guide for details
		input  wire        i_ch1_pcs_pclk,                                 //         .i_ch1_pcs_pclk,                                 Check User Guide for details
		input  wire        i_ch1_pcs_pipe_rstn,                            //         .i_ch1_pcs_pipe_rstn,                            Check User Guide for details
		input  wire        i_ch1_txpipe_asyncpowerchangeack,               //         .i_ch1_txpipe_asyncpowerchangeack,               Check User Guide for details
		input  wire        i_ch1_txpipe_blockaligncontrol,                 //         .i_ch1_txpipe_blockaligncontrol,                 Check User Guide for details
		input  wire        i_ch1_txpipe_cfg_hw_auto_sp_dis,                //         .i_ch1_txpipe_cfg_hw_auto_sp_dis,                Check User Guide for details
		input  wire        i_ch1_txpipe_dirchange,                         //         .i_ch1_txpipe_dirchange,                         Check User Guide for details
		input  wire        i_ch1_txpipe_ebuf_mode,                         //         .i_ch1_txpipe_ebuf_mode,                         Check User Guide for details
		input  wire        i_ch1_txpipe_encodedecodebypass,                //         .i_ch1_txpipe_encodedecodebypass,                Check User Guide for details
		input  wire [5:0]  i_ch1_txpipe_fs,                                //         .i_ch1_txpipe_fs,                                Check User Guide for details
		input  wire        i_ch1_txpipe_getlocalpresetcoefficients,        //         .i_ch1_txpipe_getlocalpresetcoefficients,        Check User Guide for details
		input  wire        i_ch1_txpipe_invalidrequest,                    //         .i_ch1_txpipe_invalidrequest,                    Check User Guide for details
		input  wire [5:0]  i_ch1_txpipe_lf,                                //         .i_ch1_txpipe_lf,                                Check User Guide for details
		input  wire [4:0]  i_ch1_txpipe_localpresetindex,                  //         .i_ch1_txpipe_localpresetindex,                  Check User Guide for details
		input  wire        i_ch1_txpipe_lowpin_nt,                         //         .i_ch1_txpipe_lowpin_nt,                         Check User Guide for details
		input  wire [7:0]  i_ch1_txpipe_m2p_bus,                           //         .i_ch1_txpipe_m2p_bus,                           Check User Guide for details
		input  wire [2:0]  i_ch1_txpipe_pclk_rate,                         //         .i_ch1_txpipe_pclk_rate,                         Check User Guide for details
		input  wire        i_ch1_txpipe_pclkchangeack,                     //         .i_ch1_txpipe_pclkchangeack,                     Check User Guide for details
		input  wire [3:0]  i_ch1_txpipe_phy_mode_nt,                       //         .i_ch1_txpipe_phy_mode_nt,                       Check User Guide for details
		input  wire [3:0]  i_ch1_txpipe_powerdown,                         //         .i_ch1_txpipe_powerdown,                         Check User Guide for details
		input  wire [2:0]  i_ch1_txpipe_rate,                              //         .i_ch1_txpipe_rate,                              Check User Guide for details
		input  wire        i_ch1_txpipe_rxelecidle_disable_a,              //         .i_ch1_txpipe_rxelecidle_disable_a,              Check User Guide for details
		input  wire        i_ch1_txpipe_rxeqclr,                           //         .i_ch1_txpipe_rxeqclr,                           Check User Guide for details
		input  wire        i_ch1_txpipe_rxeqeval,                          //         .i_ch1_txpipe_rxeqeval,                          Check User Guide for details
		input  wire        i_ch1_txpipe_rxeqinprogress,                    //         .i_ch1_txpipe_rxeqinprogress,                    Check User Guide for details
		input  wire        i_ch1_txpipe_rxeqtraining,                      //         .i_ch1_txpipe_rxeqtraining,                      Check User Guide for details
		input  wire        i_ch1_txpipe_rxpolarity,                        //         .i_ch1_txpipe_rxpolarity,                        Check User Guide for details
		input  wire [2:0]  i_ch1_txpipe_rxpresethint,                      //         .i_ch1_txpipe_rxpresethint,                      Check User Guide for details
		input  wire        i_ch1_txpipe_rxstandby,                         //         .i_ch1_txpipe_rxstandby,                         Check User Guide for details
		input  wire        i_ch1_txpipe_rxtermination,                     //         .i_ch1_txpipe_rxtermination,                     Check User Guide for details
		input  wire        i_ch1_txpipe_srisenable,                        //         .i_ch1_txpipe_srisenable,                        Check User Guide for details
		input  wire        i_ch1_txpipe_txcmnmode_disable_a,               //         .i_ch1_txpipe_txcmnmode_disable_a,               Check User Guide for details
		input  wire        i_ch1_txpipe_txcompliance,                      //         .i_ch1_txpipe_txcompliance,                      Check User Guide for details
		input  wire [39:0] i_ch1_txpipe_txdata,                            //         .i_ch1_txpipe_txdata,                            Check User Guide for details
		input  wire [3:0]  i_ch1_txpipe_txdatak,                           //         .i_ch1_txpipe_txdatak,                           Check User Guide for details
		input  wire        i_ch1_txpipe_txdatavalid,                       //         .i_ch1_txpipe_txdatavalid,                       Check User Guide for details
		input  wire [17:0] i_ch1_txpipe_txdeemph,                          //         .i_ch1_txpipe_txdeemph,                          Check User Guide for details
		input  wire        i_ch1_txpipe_txdtctrx_lb,                       //         .i_ch1_txpipe_txdtctrx_lb,                       Check User Guide for details
		input  wire        i_ch1_txpipe_txelecidle,                        //         .i_ch1_txpipe_txelecidle,                        Check User Guide for details
		input  wire [2:0]  i_ch1_txpipe_txmargin,                          //         .i_ch1_txpipe_txmargin,                          Check User Guide for details
		input  wire        i_ch1_txpipe_txoneszeros,                       //         .i_ch1_txpipe_txoneszeros,                       Check User Guide for details
		input  wire        i_ch1_txpipe_txstartblock,                      //         .i_ch1_txpipe_txstartblock,                      Check User Guide for details
		input  wire        i_ch1_txpipe_txswing,                           //         .i_ch1_txpipe_txswing,                           Check User Guide for details
		input  wire [3:0]  i_ch1_txpipe_txsyncheader,                      //         .i_ch1_txpipe_txsyncheader,                      Check User Guide for details
		input  wire [2:0]  i_ch1_txpipe_width,                             //         .i_ch1_txpipe_width,                             Check User Guide for details
		input  wire        i_ch1_uxq_rxcdrlock2dataa,                      //         .i_ch1_uxq_rxcdrlock2dataa,                      Check User Guide for details
		input  wire [13:0] i_ch1_uxq_rxeq_best_eye_vala,                   //         .i_ch1_uxq_rxeq_best_eye_vala,                   Check User Guide for details
		input  wire        i_ch1_uxq_rxeq_donea,                           //         .i_ch1_uxq_rxeq_donea,                           Check User Guide for details
		input  wire        i_ch1_uxq_rxmargin_nacka,                       //         .i_ch1_uxq_rxmargin_nacka,                       Check User Guide for details
		input  wire [1:0]  i_ch1_uxq_rxmargin_status_gray_a,               //         .i_ch1_uxq_rxmargin_status_gray_a,               Check User Guide for details
		input  wire        i_ch1_uxq_rxmargin_statusa,                     //         .i_ch1_uxq_rxmargin_statusa,                     Check User Guide for details
		input  wire        i_ch1_uxq_rxsignaldetect_lfpsa,                 //         .i_ch1_uxq_rxsignaldetect_lfpsa,                 Check User Guide for details
		input  wire        i_ch1_uxq_rxsignaldetecta,                      //         .i_ch1_uxq_rxsignaldetecta,                      Check User Guide for details
		input  wire        i_ch1_uxq_rxstatusa,                            //         .i_ch1_uxq_rxstatusa,                            Check User Guide for details
		input  wire [39:0] i_ch1_uxq_rxword,                               //         .i_ch1_uxq_rxword,                               Check User Guide for details
		input  wire        i_ch1_uxq_synthlcfast_postdiv,                  //         .i_ch1_uxq_synthlcfast_postdiv,                  Check User Guide for details
		input  wire        i_ch1_uxq_synthlcmed_postdiv,                   //         .i_ch1_uxq_synthlcmed_postdiv,                   Check User Guide for details
		input  wire        i_ch1_uxq_synthlcslow_postdiv,                  //         .i_ch1_uxq_synthlcslow_postdiv,                  Check User Guide for details
		input  wire        i_ch1_uxq_txdetectrx_acka,                      //         .i_ch1_uxq_txdetectrx_acka,                      Check User Guide for details
		input  wire        i_ch1_uxq_txdetectrx_statct,                    //         .i_ch1_uxq_txdetectrx_statct,                    Check User Guide for details
		input  wire        i_ch1_uxq_txstatusa,                            //         .i_ch1_uxq_txstatusa,                            Check User Guide for details
		output wire [31:0] o_ch1_lavmm_pcie_rdata,                         //         .o_ch1_lavmm_pcie_rdata,                         Check User Guide for details
		output wire        o_ch1_lavmm_pcie_rdata_valid,                   //         .o_ch1_lavmm_pcie_rdata_valid,                   Check User Guide for details
		output wire        o_ch1_lavmm_pcie_waitreq,                       //         .o_ch1_lavmm_pcie_waitreq,                       Check User Guide for details
		output wire        o_ch1_pcs_pclk,                                 //         .o_ch1_pcs_pclk,                                 Check User Guide for details
		output wire        o_ch1_pcs_pipe_rstn,                            //         .o_ch1_pcs_pipe_rstn,                            Check User Guide for details
		output wire [5:0]  o_ch1_rxpipe_dirfeedback,                       //         .o_ch1_rxpipe_dirfeedback,                       Check User Guide for details
		output wire [7:0]  o_ch1_rxpipe_linkevaluationfeedbackfiguremerit, //         .o_ch1_rxpipe_linkevaluationfeedbackfiguremerit, Check User Guide for details
		output wire [5:0]  o_ch1_rxpipe_localfs,                           //         .o_ch1_rxpipe_localfs,                           Check User Guide for details
		output wire [5:0]  o_ch1_rxpipe_locallf,                           //         .o_ch1_rxpipe_locallf,                           Check User Guide for details
		output wire        o_ch1_rxpipe_localtxcoefficientsvalid,          //         .o_ch1_rxpipe_localtxcoefficientsvalid,          Check User Guide for details
		output wire [17:0] o_ch1_rxpipe_localtxpresetcoefficients,         //         .o_ch1_rxpipe_localtxpresetcoefficients,         Check User Guide for details
		output wire [7:0]  o_ch1_rxpipe_p2m_bus,                           //         .o_ch1_rxpipe_p2m_bus,                           Check User Guide for details
		output wire        o_ch1_rxpipe_pclkchangeok,                      //         .o_ch1_rxpipe_pclkchangeok,                      Check User Guide for details
		output wire        o_ch1_rxpipe_phystatus,                         //         .o_ch1_rxpipe_phystatus,                         Check User Guide for details
		output wire [39:0] o_ch1_rxpipe_rxdata,                            //         .o_ch1_rxpipe_rxdata,                            Check User Guide for details
		output wire [3:0]  o_ch1_rxpipe_rxdatak,                           //         .o_ch1_rxpipe_rxdatak,                           Check User Guide for details
		output wire        o_ch1_rxpipe_rxdatavalid,                       //         .o_ch1_rxpipe_rxdatavalid,                       Check User Guide for details
		output wire        o_ch1_rxpipe_rxelecidlea,                       //         .o_ch1_rxpipe_rxelecidlea,                       Check User Guide for details
		output wire        o_ch1_rxpipe_rxstandbystatus,                   //         .o_ch1_rxpipe_rxstandbystatus,                   Check User Guide for details
		output wire        o_ch1_rxpipe_rxstartblock,                      //         .o_ch1_rxpipe_rxstartblock,                      Check User Guide for details
		output wire [2:0]  o_ch1_rxpipe_rxstatus,                          //         .o_ch1_rxpipe_rxstatus,                          Check User Guide for details
		output wire [3:0]  o_ch1_rxpipe_rxsyncheader,                      //         .o_ch1_rxpipe_rxsyncheader,                      Check User Guide for details
		output wire        o_ch1_rxpipe_rxvalid,                           //         .o_ch1_rxpipe_rxvalid,                           Check User Guide for details
		output wire        o_ch1_ux_ock_pma_clk,                           //         .o_ch1_ux_ock_pma_clk,                           Check User Guide for details
		output wire        o_ch1_uxq_lfps_ennt,                            //         .o_ch1_uxq_lfps_ennt,                            Check User Guide for details
		output wire [1:0]  o_ch1_uxq_pcie_l1ctrla,                         //         .o_ch1_uxq_pcie_l1ctrla,                         Check User Guide for details
		output wire        o_ch1_uxq_pma_cmn_ctrl,                         //         .o_ch1_uxq_pma_cmn_ctrl,                         Check User Guide for details
		output wire        o_ch1_uxq_pma_ctrl,                             //         .o_ch1_uxq_pma_ctrl,                             Check User Guide for details
		output wire        o_ch1_uxq_rst_pcs_rx_b_a,                       //         .o_ch1_uxq_rst_pcs_rx_b_a,                       Check User Guide for details
		output wire        o_ch1_uxq_rst_pcs_tx_b_a,                       //         .o_ch1_uxq_rst_pcs_tx_b_a,                       Check User Guide for details
		output wire        o_ch1_uxq_rxeiosdetectstata,                    //         .o_ch1_uxq_rxeiosdetectstata,                    Check User Guide for details
		output wire [2:0]  o_ch1_uxq_rxeq_precal_code_selnt,               //         .o_ch1_uxq_rxeq_precal_code_selnt,               Check User Guide for details
		output wire        o_ch1_uxq_rxeq_starta,                          //         .o_ch1_uxq_rxeq_starta,                          Check User Guide for details
		output wire        o_ch1_uxq_rxeq_static_ena,                      //         .o_ch1_uxq_rxeq_static_ena,                      Check User Guide for details
		output wire        o_ch1_uxq_rxmargin_direction_nt,                //         .o_ch1_uxq_rxmargin_direction_nt,                Check User Guide for details
		output wire        o_ch1_uxq_rxmargin_mode_nt,                     //         .o_ch1_uxq_rxmargin_mode_nt,                     Check User Guide for details
		output wire        o_ch1_uxq_rxmargin_offset_change_a,             //         .o_ch1_uxq_rxmargin_offset_change_a,             Check User Guide for details
		output wire [6:0]  o_ch1_uxq_rxmargin_offset_nt,                   //         .o_ch1_uxq_rxmargin_offset_nt,                   Check User Guide for details
		output wire        o_ch1_uxq_rxmargin_start_a,                     //         .o_ch1_uxq_rxmargin_start_a,                     Check User Guide for details
		output wire [2:0]  o_ch1_uxq_rxpstate,                             //         .o_ch1_uxq_rxpstate,                             Check User Guide for details
		output wire [3:0]  o_ch1_uxq_rxrate,                               //         .o_ch1_uxq_rxrate,                               Check User Guide for details
		output wire        o_ch1_uxq_rxterm_hiz_ena,                       //         .o_ch1_uxq_rxterm_hiz_ena,                       Check User Guide for details
		output wire [2:0]  o_ch1_uxq_rxwidth,                              //         .o_ch1_uxq_rxwidth,                              Check User Guide for details
		output wire        o_ch1_uxq_tstbus_lane,                          //         .o_ch1_uxq_tstbus_lane,                          Check User Guide for details
		output wire        o_ch1_uxq_txbeacona,                            //         .o_ch1_uxq_txbeacona,                            Check User Guide for details
		output wire [2:0]  o_ch1_uxq_txclkdivrate,                         //         .o_ch1_uxq_txclkdivrate,                         Check User Guide for details
		output wire        o_ch1_uxq_txdetectrx_reqa,                      //         .o_ch1_uxq_txdetectrx_reqa,                      Check User Guide for details
		output wire [5:0]  o_ch1_uxq_txdrv_levn,                           //         .o_ch1_uxq_txdrv_levn,                           Check User Guide for details
		output wire [4:0]  o_ch1_uxq_txdrv_levnm1,                         //         .o_ch1_uxq_txdrv_levnm1,                         Check User Guide for details
		output wire [2:0]  o_ch1_uxq_txdrv_levnm2,                         //         .o_ch1_uxq_txdrv_levnm2,                         Check User Guide for details
		output wire [4:0]  o_ch1_uxq_txdrv_levnp1,                         //         .o_ch1_uxq_txdrv_levnp1,                         Check User Guide for details
		output wire [3:0]  o_ch1_uxq_txdrv_slew,                           //         .o_ch1_uxq_txdrv_slew,                           Check User Guide for details
		output wire [3:0]  o_ch1_uxq_txelecidle,                           //         .o_ch1_uxq_txelecidle,                           Check User Guide for details
		output wire [2:0]  o_ch1_uxq_txpstate,                             //         .o_ch1_uxq_txpstate,                             Check User Guide for details
		output wire [3:0]  o_ch1_uxq_txrate,                               //         .o_ch1_uxq_txrate,                               Check User Guide for details
		output wire [2:0]  o_ch1_uxq_txwidth,                              //         .o_ch1_uxq_txwidth,                              Check User Guide for details
		output wire [39:0] o_ch1_uxq_txword,                               //         .o_ch1_uxq_txword,                               Check User Guide for details
		input  wire [16:0] i_ch2_lavmm_pcie_addr,                          //         .i_ch2_lavmm_pcie_addr,                          Check User Guide for details
		input  wire [3:0]  i_ch2_lavmm_pcie_be,                            //         .i_ch2_lavmm_pcie_be,                            Check User Guide for details
		input  wire        i_ch2_lavmm_pcie_clk,                           //         .i_ch2_lavmm_pcie_clk,                           Check User Guide for details
		input  wire        i_ch2_lavmm_pcie_read,                          //         .i_ch2_lavmm_pcie_read,                          Check User Guide for details
		input  wire        i_ch2_lavmm_pcie_rstn,                          //         .i_ch2_lavmm_pcie_rstn,                          Check User Guide for details
		input  wire [31:0] i_ch2_lavmm_pcie_wdata,                         //         .i_ch2_lavmm_pcie_wdata,                         Check User Guide for details
		input  wire        i_ch2_lavmm_pcie_write,                         //         .i_ch2_lavmm_pcie_write,                         Check User Guide for details
		input  wire        i_ch2_pcie_rxword_clk,                          //         .i_ch2_pcie_rxword_clk,                          Check User Guide for details
		input  wire        i_ch2_pcie_txword_clk,                          //         .i_ch2_pcie_txword_clk,                          Check User Guide for details
		input  wire        i_ch2_pcs_pclk,                                 //         .i_ch2_pcs_pclk,                                 Check User Guide for details
		input  wire        i_ch2_pcs_pipe_rstn,                            //         .i_ch2_pcs_pipe_rstn,                            Check User Guide for details
		input  wire        i_ch2_txpipe_asyncpowerchangeack,               //         .i_ch2_txpipe_asyncpowerchangeack,               Check User Guide for details
		input  wire        i_ch2_txpipe_blockaligncontrol,                 //         .i_ch2_txpipe_blockaligncontrol,                 Check User Guide for details
		input  wire        i_ch2_txpipe_cfg_hw_auto_sp_dis,                //         .i_ch2_txpipe_cfg_hw_auto_sp_dis,                Check User Guide for details
		input  wire        i_ch2_txpipe_dirchange,                         //         .i_ch2_txpipe_dirchange,                         Check User Guide for details
		input  wire        i_ch2_txpipe_ebuf_mode,                         //         .i_ch2_txpipe_ebuf_mode,                         Check User Guide for details
		input  wire        i_ch2_txpipe_encodedecodebypass,                //         .i_ch2_txpipe_encodedecodebypass,                Check User Guide for details
		input  wire [5:0]  i_ch2_txpipe_fs,                                //         .i_ch2_txpipe_fs,                                Check User Guide for details
		input  wire        i_ch2_txpipe_getlocalpresetcoefficients,        //         .i_ch2_txpipe_getlocalpresetcoefficients,        Check User Guide for details
		input  wire        i_ch2_txpipe_invalidrequest,                    //         .i_ch2_txpipe_invalidrequest,                    Check User Guide for details
		input  wire [5:0]  i_ch2_txpipe_lf,                                //         .i_ch2_txpipe_lf,                                Check User Guide for details
		input  wire [4:0]  i_ch2_txpipe_localpresetindex,                  //         .i_ch2_txpipe_localpresetindex,                  Check User Guide for details
		input  wire        i_ch2_txpipe_lowpin_nt,                         //         .i_ch2_txpipe_lowpin_nt,                         Check User Guide for details
		input  wire [7:0]  i_ch2_txpipe_m2p_bus,                           //         .i_ch2_txpipe_m2p_bus,                           Check User Guide for details
		input  wire [2:0]  i_ch2_txpipe_pclk_rate,                         //         .i_ch2_txpipe_pclk_rate,                         Check User Guide for details
		input  wire        i_ch2_txpipe_pclkchangeack,                     //         .i_ch2_txpipe_pclkchangeack,                     Check User Guide for details
		input  wire [3:0]  i_ch2_txpipe_phy_mode_nt,                       //         .i_ch2_txpipe_phy_mode_nt,                       Check User Guide for details
		input  wire [3:0]  i_ch2_txpipe_powerdown,                         //         .i_ch2_txpipe_powerdown,                         Check User Guide for details
		input  wire [2:0]  i_ch2_txpipe_rate,                              //         .i_ch2_txpipe_rate,                              Check User Guide for details
		input  wire        i_ch2_txpipe_rxelecidle_disable_a,              //         .i_ch2_txpipe_rxelecidle_disable_a,              Check User Guide for details
		input  wire        i_ch2_txpipe_rxeqclr,                           //         .i_ch2_txpipe_rxeqclr,                           Check User Guide for details
		input  wire        i_ch2_txpipe_rxeqeval,                          //         .i_ch2_txpipe_rxeqeval,                          Check User Guide for details
		input  wire        i_ch2_txpipe_rxeqinprogress,                    //         .i_ch2_txpipe_rxeqinprogress,                    Check User Guide for details
		input  wire        i_ch2_txpipe_rxeqtraining,                      //         .i_ch2_txpipe_rxeqtraining,                      Check User Guide for details
		input  wire        i_ch2_txpipe_rxpolarity,                        //         .i_ch2_txpipe_rxpolarity,                        Check User Guide for details
		input  wire [2:0]  i_ch2_txpipe_rxpresethint,                      //         .i_ch2_txpipe_rxpresethint,                      Check User Guide for details
		input  wire        i_ch2_txpipe_rxstandby,                         //         .i_ch2_txpipe_rxstandby,                         Check User Guide for details
		input  wire        i_ch2_txpipe_rxtermination,                     //         .i_ch2_txpipe_rxtermination,                     Check User Guide for details
		input  wire        i_ch2_txpipe_srisenable,                        //         .i_ch2_txpipe_srisenable,                        Check User Guide for details
		input  wire        i_ch2_txpipe_txcmnmode_disable_a,               //         .i_ch2_txpipe_txcmnmode_disable_a,               Check User Guide for details
		input  wire        i_ch2_txpipe_txcompliance,                      //         .i_ch2_txpipe_txcompliance,                      Check User Guide for details
		input  wire [39:0] i_ch2_txpipe_txdata,                            //         .i_ch2_txpipe_txdata,                            Check User Guide for details
		input  wire [3:0]  i_ch2_txpipe_txdatak,                           //         .i_ch2_txpipe_txdatak,                           Check User Guide for details
		input  wire        i_ch2_txpipe_txdatavalid,                       //         .i_ch2_txpipe_txdatavalid,                       Check User Guide for details
		input  wire [17:0] i_ch2_txpipe_txdeemph,                          //         .i_ch2_txpipe_txdeemph,                          Check User Guide for details
		input  wire        i_ch2_txpipe_txdtctrx_lb,                       //         .i_ch2_txpipe_txdtctrx_lb,                       Check User Guide for details
		input  wire        i_ch2_txpipe_txelecidle,                        //         .i_ch2_txpipe_txelecidle,                        Check User Guide for details
		input  wire [2:0]  i_ch2_txpipe_txmargin,                          //         .i_ch2_txpipe_txmargin,                          Check User Guide for details
		input  wire        i_ch2_txpipe_txoneszeros,                       //         .i_ch2_txpipe_txoneszeros,                       Check User Guide for details
		input  wire        i_ch2_txpipe_txstartblock,                      //         .i_ch2_txpipe_txstartblock,                      Check User Guide for details
		input  wire        i_ch2_txpipe_txswing,                           //         .i_ch2_txpipe_txswing,                           Check User Guide for details
		input  wire [3:0]  i_ch2_txpipe_txsyncheader,                      //         .i_ch2_txpipe_txsyncheader,                      Check User Guide for details
		input  wire [2:0]  i_ch2_txpipe_width,                             //         .i_ch2_txpipe_width,                             Check User Guide for details
		input  wire        i_ch2_uxq_rxcdrlock2dataa,                      //         .i_ch2_uxq_rxcdrlock2dataa,                      Check User Guide for details
		input  wire [13:0] i_ch2_uxq_rxeq_best_eye_vala,                   //         .i_ch2_uxq_rxeq_best_eye_vala,                   Check User Guide for details
		input  wire        i_ch2_uxq_rxeq_donea,                           //         .i_ch2_uxq_rxeq_donea,                           Check User Guide for details
		input  wire        i_ch2_uxq_rxmargin_nacka,                       //         .i_ch2_uxq_rxmargin_nacka,                       Check User Guide for details
		input  wire [1:0]  i_ch2_uxq_rxmargin_status_gray_a,               //         .i_ch2_uxq_rxmargin_status_gray_a,               Check User Guide for details
		input  wire        i_ch2_uxq_rxmargin_statusa,                     //         .i_ch2_uxq_rxmargin_statusa,                     Check User Guide for details
		input  wire        i_ch2_uxq_rxsignaldetect_lfpsa,                 //         .i_ch2_uxq_rxsignaldetect_lfpsa,                 Check User Guide for details
		input  wire        i_ch2_uxq_rxsignaldetecta,                      //         .i_ch2_uxq_rxsignaldetecta,                      Check User Guide for details
		input  wire        i_ch2_uxq_rxstatusa,                            //         .i_ch2_uxq_rxstatusa,                            Check User Guide for details
		input  wire [39:0] i_ch2_uxq_rxword,                               //         .i_ch2_uxq_rxword,                               Check User Guide for details
		input  wire        i_ch2_uxq_synthlcfast_postdiv,                  //         .i_ch2_uxq_synthlcfast_postdiv,                  Check User Guide for details
		input  wire        i_ch2_uxq_synthlcmed_postdiv,                   //         .i_ch2_uxq_synthlcmed_postdiv,                   Check User Guide for details
		input  wire        i_ch2_uxq_synthlcslow_postdiv,                  //         .i_ch2_uxq_synthlcslow_postdiv,                  Check User Guide for details
		input  wire        i_ch2_uxq_txdetectrx_acka,                      //         .i_ch2_uxq_txdetectrx_acka,                      Check User Guide for details
		input  wire        i_ch2_uxq_txdetectrx_statct,                    //         .i_ch2_uxq_txdetectrx_statct,                    Check User Guide for details
		input  wire        i_ch2_uxq_txstatusa,                            //         .i_ch2_uxq_txstatusa,                            Check User Guide for details
		output wire [31:0] o_ch2_lavmm_pcie_rdata,                         //         .o_ch2_lavmm_pcie_rdata,                         Check User Guide for details
		output wire        o_ch2_lavmm_pcie_rdata_valid,                   //         .o_ch2_lavmm_pcie_rdata_valid,                   Check User Guide for details
		output wire        o_ch2_lavmm_pcie_waitreq,                       //         .o_ch2_lavmm_pcie_waitreq,                       Check User Guide for details
		output wire        o_ch2_pcs_pclk,                                 //         .o_ch2_pcs_pclk,                                 Check User Guide for details
		output wire        o_ch2_pcs_pipe_rstn,                            //         .o_ch2_pcs_pipe_rstn,                            Check User Guide for details
		output wire [5:0]  o_ch2_rxpipe_dirfeedback,                       //         .o_ch2_rxpipe_dirfeedback,                       Check User Guide for details
		output wire [7:0]  o_ch2_rxpipe_linkevaluationfeedbackfiguremerit, //         .o_ch2_rxpipe_linkevaluationfeedbackfiguremerit, Check User Guide for details
		output wire [5:0]  o_ch2_rxpipe_localfs,                           //         .o_ch2_rxpipe_localfs,                           Check User Guide for details
		output wire [5:0]  o_ch2_rxpipe_locallf,                           //         .o_ch2_rxpipe_locallf,                           Check User Guide for details
		output wire        o_ch2_rxpipe_localtxcoefficientsvalid,          //         .o_ch2_rxpipe_localtxcoefficientsvalid,          Check User Guide for details
		output wire [17:0] o_ch2_rxpipe_localtxpresetcoefficients,         //         .o_ch2_rxpipe_localtxpresetcoefficients,         Check User Guide for details
		output wire [7:0]  o_ch2_rxpipe_p2m_bus,                           //         .o_ch2_rxpipe_p2m_bus,                           Check User Guide for details
		output wire        o_ch2_rxpipe_pclkchangeok,                      //         .o_ch2_rxpipe_pclkchangeok,                      Check User Guide for details
		output wire        o_ch2_rxpipe_phystatus,                         //         .o_ch2_rxpipe_phystatus,                         Check User Guide for details
		output wire [39:0] o_ch2_rxpipe_rxdata,                            //         .o_ch2_rxpipe_rxdata,                            Check User Guide for details
		output wire [3:0]  o_ch2_rxpipe_rxdatak,                           //         .o_ch2_rxpipe_rxdatak,                           Check User Guide for details
		output wire        o_ch2_rxpipe_rxdatavalid,                       //         .o_ch2_rxpipe_rxdatavalid,                       Check User Guide for details
		output wire        o_ch2_rxpipe_rxelecidlea,                       //         .o_ch2_rxpipe_rxelecidlea,                       Check User Guide for details
		output wire        o_ch2_rxpipe_rxstandbystatus,                   //         .o_ch2_rxpipe_rxstandbystatus,                   Check User Guide for details
		output wire        o_ch2_rxpipe_rxstartblock,                      //         .o_ch2_rxpipe_rxstartblock,                      Check User Guide for details
		output wire [2:0]  o_ch2_rxpipe_rxstatus,                          //         .o_ch2_rxpipe_rxstatus,                          Check User Guide for details
		output wire [3:0]  o_ch2_rxpipe_rxsyncheader,                      //         .o_ch2_rxpipe_rxsyncheader,                      Check User Guide for details
		output wire        o_ch2_rxpipe_rxvalid,                           //         .o_ch2_rxpipe_rxvalid,                           Check User Guide for details
		output wire        o_ch2_ux_ock_pma_clk,                           //         .o_ch2_ux_ock_pma_clk,                           Check User Guide for details
		output wire        o_ch2_uxq_lfps_ennt,                            //         .o_ch2_uxq_lfps_ennt,                            Check User Guide for details
		output wire [1:0]  o_ch2_uxq_pcie_l1ctrla,                         //         .o_ch2_uxq_pcie_l1ctrla,                         Check User Guide for details
		output wire        o_ch2_uxq_pma_cmn_ctrl,                         //         .o_ch2_uxq_pma_cmn_ctrl,                         Check User Guide for details
		output wire        o_ch2_uxq_pma_ctrl,                             //         .o_ch2_uxq_pma_ctrl,                             Check User Guide for details
		output wire        o_ch2_uxq_rst_pcs_rx_b_a,                       //         .o_ch2_uxq_rst_pcs_rx_b_a,                       Check User Guide for details
		output wire        o_ch2_uxq_rst_pcs_tx_b_a,                       //         .o_ch2_uxq_rst_pcs_tx_b_a,                       Check User Guide for details
		output wire        o_ch2_uxq_rxeiosdetectstata,                    //         .o_ch2_uxq_rxeiosdetectstata,                    Check User Guide for details
		output wire [2:0]  o_ch2_uxq_rxeq_precal_code_selnt,               //         .o_ch2_uxq_rxeq_precal_code_selnt,               Check User Guide for details
		output wire        o_ch2_uxq_rxeq_starta,                          //         .o_ch2_uxq_rxeq_starta,                          Check User Guide for details
		output wire        o_ch2_uxq_rxeq_static_ena,                      //         .o_ch2_uxq_rxeq_static_ena,                      Check User Guide for details
		output wire        o_ch2_uxq_rxmargin_direction_nt,                //         .o_ch2_uxq_rxmargin_direction_nt,                Check User Guide for details
		output wire        o_ch2_uxq_rxmargin_mode_nt,                     //         .o_ch2_uxq_rxmargin_mode_nt,                     Check User Guide for details
		output wire        o_ch2_uxq_rxmargin_offset_change_a,             //         .o_ch2_uxq_rxmargin_offset_change_a,             Check User Guide for details
		output wire [6:0]  o_ch2_uxq_rxmargin_offset_nt,                   //         .o_ch2_uxq_rxmargin_offset_nt,                   Check User Guide for details
		output wire        o_ch2_uxq_rxmargin_start_a,                     //         .o_ch2_uxq_rxmargin_start_a,                     Check User Guide for details
		output wire [2:0]  o_ch2_uxq_rxpstate,                             //         .o_ch2_uxq_rxpstate,                             Check User Guide for details
		output wire [3:0]  o_ch2_uxq_rxrate,                               //         .o_ch2_uxq_rxrate,                               Check User Guide for details
		output wire        o_ch2_uxq_rxterm_hiz_ena,                       //         .o_ch2_uxq_rxterm_hiz_ena,                       Check User Guide for details
		output wire [2:0]  o_ch2_uxq_rxwidth,                              //         .o_ch2_uxq_rxwidth,                              Check User Guide for details
		output wire        o_ch2_uxq_tstbus_lane,                          //         .o_ch2_uxq_tstbus_lane,                          Check User Guide for details
		output wire        o_ch2_uxq_txbeacona,                            //         .o_ch2_uxq_txbeacona,                            Check User Guide for details
		output wire [2:0]  o_ch2_uxq_txclkdivrate,                         //         .o_ch2_uxq_txclkdivrate,                         Check User Guide for details
		output wire        o_ch2_uxq_txdetectrx_reqa,                      //         .o_ch2_uxq_txdetectrx_reqa,                      Check User Guide for details
		output wire [5:0]  o_ch2_uxq_txdrv_levn,                           //         .o_ch2_uxq_txdrv_levn,                           Check User Guide for details
		output wire [4:0]  o_ch2_uxq_txdrv_levnm1,                         //         .o_ch2_uxq_txdrv_levnm1,                         Check User Guide for details
		output wire [2:0]  o_ch2_uxq_txdrv_levnm2,                         //         .o_ch2_uxq_txdrv_levnm2,                         Check User Guide for details
		output wire [4:0]  o_ch2_uxq_txdrv_levnp1,                         //         .o_ch2_uxq_txdrv_levnp1,                         Check User Guide for details
		output wire [3:0]  o_ch2_uxq_txdrv_slew,                           //         .o_ch2_uxq_txdrv_slew,                           Check User Guide for details
		output wire [3:0]  o_ch2_uxq_txelecidle,                           //         .o_ch2_uxq_txelecidle,                           Check User Guide for details
		output wire [2:0]  o_ch2_uxq_txpstate,                             //         .o_ch2_uxq_txpstate,                             Check User Guide for details
		output wire [3:0]  o_ch2_uxq_txrate,                               //         .o_ch2_uxq_txrate,                               Check User Guide for details
		output wire [2:0]  o_ch2_uxq_txwidth,                              //         .o_ch2_uxq_txwidth,                              Check User Guide for details
		output wire [39:0] o_ch2_uxq_txword,                               //         .o_ch2_uxq_txword,                               Check User Guide for details
		input  wire [16:0] i_ch3_lavmm_pcie_addr,                          //         .i_ch3_lavmm_pcie_addr,                          Check User Guide for details
		input  wire [3:0]  i_ch3_lavmm_pcie_be,                            //         .i_ch3_lavmm_pcie_be,                            Check User Guide for details
		input  wire        i_ch3_lavmm_pcie_clk,                           //         .i_ch3_lavmm_pcie_clk,                           Check User Guide for details
		input  wire        i_ch3_lavmm_pcie_read,                          //         .i_ch3_lavmm_pcie_read,                          Check User Guide for details
		input  wire        i_ch3_lavmm_pcie_rstn,                          //         .i_ch3_lavmm_pcie_rstn,                          Check User Guide for details
		input  wire [31:0] i_ch3_lavmm_pcie_wdata,                         //         .i_ch3_lavmm_pcie_wdata,                         Check User Guide for details
		input  wire        i_ch3_lavmm_pcie_write,                         //         .i_ch3_lavmm_pcie_write,                         Check User Guide for details
		input  wire        i_ch3_pcie_rxword_clk,                          //         .i_ch3_pcie_rxword_clk,                          Check User Guide for details
		input  wire        i_ch3_pcie_txword_clk,                          //         .i_ch3_pcie_txword_clk,                          Check User Guide for details
		input  wire        i_ch3_pcs_pclk,                                 //         .i_ch3_pcs_pclk,                                 Check User Guide for details
		input  wire        i_ch3_pcs_pipe_rstn,                            //         .i_ch3_pcs_pipe_rstn,                            Check User Guide for details
		input  wire        i_ch3_txpipe_asyncpowerchangeack,               //         .i_ch3_txpipe_asyncpowerchangeack,               Check User Guide for details
		input  wire        i_ch3_txpipe_blockaligncontrol,                 //         .i_ch3_txpipe_blockaligncontrol,                 Check User Guide for details
		input  wire        i_ch3_txpipe_cfg_hw_auto_sp_dis,                //         .i_ch3_txpipe_cfg_hw_auto_sp_dis,                Check User Guide for details
		input  wire        i_ch3_txpipe_dirchange,                         //         .i_ch3_txpipe_dirchange,                         Check User Guide for details
		input  wire        i_ch3_txpipe_ebuf_mode,                         //         .i_ch3_txpipe_ebuf_mode,                         Check User Guide for details
		input  wire        i_ch3_txpipe_encodedecodebypass,                //         .i_ch3_txpipe_encodedecodebypass,                Check User Guide for details
		input  wire [5:0]  i_ch3_txpipe_fs,                                //         .i_ch3_txpipe_fs,                                Check User Guide for details
		input  wire        i_ch3_txpipe_getlocalpresetcoefficients,        //         .i_ch3_txpipe_getlocalpresetcoefficients,        Check User Guide for details
		input  wire        i_ch3_txpipe_invalidrequest,                    //         .i_ch3_txpipe_invalidrequest,                    Check User Guide for details
		input  wire [5:0]  i_ch3_txpipe_lf,                                //         .i_ch3_txpipe_lf,                                Check User Guide for details
		input  wire [4:0]  i_ch3_txpipe_localpresetindex,                  //         .i_ch3_txpipe_localpresetindex,                  Check User Guide for details
		input  wire        i_ch3_txpipe_lowpin_nt,                         //         .i_ch3_txpipe_lowpin_nt,                         Check User Guide for details
		input  wire [7:0]  i_ch3_txpipe_m2p_bus,                           //         .i_ch3_txpipe_m2p_bus,                           Check User Guide for details
		input  wire [2:0]  i_ch3_txpipe_pclk_rate,                         //         .i_ch3_txpipe_pclk_rate,                         Check User Guide for details
		input  wire        i_ch3_txpipe_pclkchangeack,                     //         .i_ch3_txpipe_pclkchangeack,                     Check User Guide for details
		input  wire [3:0]  i_ch3_txpipe_phy_mode_nt,                       //         .i_ch3_txpipe_phy_mode_nt,                       Check User Guide for details
		input  wire [3:0]  i_ch3_txpipe_powerdown,                         //         .i_ch3_txpipe_powerdown,                         Check User Guide for details
		input  wire [2:0]  i_ch3_txpipe_rate,                              //         .i_ch3_txpipe_rate,                              Check User Guide for details
		input  wire        i_ch3_txpipe_rxelecidle_disable_a,              //         .i_ch3_txpipe_rxelecidle_disable_a,              Check User Guide for details
		input  wire        i_ch3_txpipe_rxeqclr,                           //         .i_ch3_txpipe_rxeqclr,                           Check User Guide for details
		input  wire        i_ch3_txpipe_rxeqeval,                          //         .i_ch3_txpipe_rxeqeval,                          Check User Guide for details
		input  wire        i_ch3_txpipe_rxeqinprogress,                    //         .i_ch3_txpipe_rxeqinprogress,                    Check User Guide for details
		input  wire        i_ch3_txpipe_rxeqtraining,                      //         .i_ch3_txpipe_rxeqtraining,                      Check User Guide for details
		input  wire        i_ch3_txpipe_rxpolarity,                        //         .i_ch3_txpipe_rxpolarity,                        Check User Guide for details
		input  wire [2:0]  i_ch3_txpipe_rxpresethint,                      //         .i_ch3_txpipe_rxpresethint,                      Check User Guide for details
		input  wire        i_ch3_txpipe_rxstandby,                         //         .i_ch3_txpipe_rxstandby,                         Check User Guide for details
		input  wire        i_ch3_txpipe_rxtermination,                     //         .i_ch3_txpipe_rxtermination,                     Check User Guide for details
		input  wire        i_ch3_txpipe_srisenable,                        //         .i_ch3_txpipe_srisenable,                        Check User Guide for details
		input  wire        i_ch3_txpipe_txcmnmode_disable_a,               //         .i_ch3_txpipe_txcmnmode_disable_a,               Check User Guide for details
		input  wire        i_ch3_txpipe_txcompliance,                      //         .i_ch3_txpipe_txcompliance,                      Check User Guide for details
		input  wire [39:0] i_ch3_txpipe_txdata,                            //         .i_ch3_txpipe_txdata,                            Check User Guide for details
		input  wire [3:0]  i_ch3_txpipe_txdatak,                           //         .i_ch3_txpipe_txdatak,                           Check User Guide for details
		input  wire        i_ch3_txpipe_txdatavalid,                       //         .i_ch3_txpipe_txdatavalid,                       Check User Guide for details
		input  wire [17:0] i_ch3_txpipe_txdeemph,                          //         .i_ch3_txpipe_txdeemph,                          Check User Guide for details
		input  wire        i_ch3_txpipe_txdtctrx_lb,                       //         .i_ch3_txpipe_txdtctrx_lb,                       Check User Guide for details
		input  wire        i_ch3_txpipe_txelecidle,                        //         .i_ch3_txpipe_txelecidle,                        Check User Guide for details
		input  wire [2:0]  i_ch3_txpipe_txmargin,                          //         .i_ch3_txpipe_txmargin,                          Check User Guide for details
		input  wire        i_ch3_txpipe_txoneszeros,                       //         .i_ch3_txpipe_txoneszeros,                       Check User Guide for details
		input  wire        i_ch3_txpipe_txstartblock,                      //         .i_ch3_txpipe_txstartblock,                      Check User Guide for details
		input  wire        i_ch3_txpipe_txswing,                           //         .i_ch3_txpipe_txswing,                           Check User Guide for details
		input  wire [3:0]  i_ch3_txpipe_txsyncheader,                      //         .i_ch3_txpipe_txsyncheader,                      Check User Guide for details
		input  wire [2:0]  i_ch3_txpipe_width,                             //         .i_ch3_txpipe_width,                             Check User Guide for details
		input  wire        i_ch3_uxq_rxcdrlock2dataa,                      //         .i_ch3_uxq_rxcdrlock2dataa,                      Check User Guide for details
		input  wire [13:0] i_ch3_uxq_rxeq_best_eye_vala,                   //         .i_ch3_uxq_rxeq_best_eye_vala,                   Check User Guide for details
		input  wire        i_ch3_uxq_rxeq_donea,                           //         .i_ch3_uxq_rxeq_donea,                           Check User Guide for details
		input  wire        i_ch3_uxq_rxmargin_nacka,                       //         .i_ch3_uxq_rxmargin_nacka,                       Check User Guide for details
		input  wire [1:0]  i_ch3_uxq_rxmargin_status_gray_a,               //         .i_ch3_uxq_rxmargin_status_gray_a,               Check User Guide for details
		input  wire        i_ch3_uxq_rxmargin_statusa,                     //         .i_ch3_uxq_rxmargin_statusa,                     Check User Guide for details
		input  wire        i_ch3_uxq_rxsignaldetect_lfpsa,                 //         .i_ch3_uxq_rxsignaldetect_lfpsa,                 Check User Guide for details
		input  wire        i_ch3_uxq_rxsignaldetecta,                      //         .i_ch3_uxq_rxsignaldetecta,                      Check User Guide for details
		input  wire        i_ch3_uxq_rxstatusa,                            //         .i_ch3_uxq_rxstatusa,                            Check User Guide for details
		input  wire [39:0] i_ch3_uxq_rxword,                               //         .i_ch3_uxq_rxword,                               Check User Guide for details
		input  wire        i_ch3_uxq_synthlcfast_postdiv,                  //         .i_ch3_uxq_synthlcfast_postdiv,                  Check User Guide for details
		input  wire        i_ch3_uxq_synthlcmed_postdiv,                   //         .i_ch3_uxq_synthlcmed_postdiv,                   Check User Guide for details
		input  wire        i_ch3_uxq_synthlcslow_postdiv,                  //         .i_ch3_uxq_synthlcslow_postdiv,                  Check User Guide for details
		input  wire        i_ch3_uxq_txdetectrx_acka,                      //         .i_ch3_uxq_txdetectrx_acka,                      Check User Guide for details
		input  wire        i_ch3_uxq_txdetectrx_statct,                    //         .i_ch3_uxq_txdetectrx_statct,                    Check User Guide for details
		input  wire        i_ch3_uxq_txstatusa,                            //         .i_ch3_uxq_txstatusa,                            Check User Guide for details
		output wire [31:0] o_ch3_lavmm_pcie_rdata,                         //         .o_ch3_lavmm_pcie_rdata,                         Check User Guide for details
		output wire        o_ch3_lavmm_pcie_rdata_valid,                   //         .o_ch3_lavmm_pcie_rdata_valid,                   Check User Guide for details
		output wire        o_ch3_lavmm_pcie_waitreq,                       //         .o_ch3_lavmm_pcie_waitreq,                       Check User Guide for details
		output wire        o_ch3_pcs_pclk,                                 //         .o_ch3_pcs_pclk,                                 Check User Guide for details
		output wire        o_ch3_pcs_pipe_rstn,                            //         .o_ch3_pcs_pipe_rstn,                            Check User Guide for details
		output wire [5:0]  o_ch3_rxpipe_dirfeedback,                       //         .o_ch3_rxpipe_dirfeedback,                       Check User Guide for details
		output wire [7:0]  o_ch3_rxpipe_linkevaluationfeedbackfiguremerit, //         .o_ch3_rxpipe_linkevaluationfeedbackfiguremerit, Check User Guide for details
		output wire [5:0]  o_ch3_rxpipe_localfs,                           //         .o_ch3_rxpipe_localfs,                           Check User Guide for details
		output wire [5:0]  o_ch3_rxpipe_locallf,                           //         .o_ch3_rxpipe_locallf,                           Check User Guide for details
		output wire        o_ch3_rxpipe_localtxcoefficientsvalid,          //         .o_ch3_rxpipe_localtxcoefficientsvalid,          Check User Guide for details
		output wire [17:0] o_ch3_rxpipe_localtxpresetcoefficients,         //         .o_ch3_rxpipe_localtxpresetcoefficients,         Check User Guide for details
		output wire [7:0]  o_ch3_rxpipe_p2m_bus,                           //         .o_ch3_rxpipe_p2m_bus,                           Check User Guide for details
		output wire        o_ch3_rxpipe_pclkchangeok,                      //         .o_ch3_rxpipe_pclkchangeok,                      Check User Guide for details
		output wire        o_ch3_rxpipe_phystatus,                         //         .o_ch3_rxpipe_phystatus,                         Check User Guide for details
		output wire [39:0] o_ch3_rxpipe_rxdata,                            //         .o_ch3_rxpipe_rxdata,                            Check User Guide for details
		output wire [3:0]  o_ch3_rxpipe_rxdatak,                           //         .o_ch3_rxpipe_rxdatak,                           Check User Guide for details
		output wire        o_ch3_rxpipe_rxdatavalid,                       //         .o_ch3_rxpipe_rxdatavalid,                       Check User Guide for details
		output wire        o_ch3_rxpipe_rxelecidlea,                       //         .o_ch3_rxpipe_rxelecidlea,                       Check User Guide for details
		output wire        o_ch3_rxpipe_rxstandbystatus,                   //         .o_ch3_rxpipe_rxstandbystatus,                   Check User Guide for details
		output wire        o_ch3_rxpipe_rxstartblock,                      //         .o_ch3_rxpipe_rxstartblock,                      Check User Guide for details
		output wire [2:0]  o_ch3_rxpipe_rxstatus,                          //         .o_ch3_rxpipe_rxstatus,                          Check User Guide for details
		output wire [3:0]  o_ch3_rxpipe_rxsyncheader,                      //         .o_ch3_rxpipe_rxsyncheader,                      Check User Guide for details
		output wire        o_ch3_rxpipe_rxvalid,                           //         .o_ch3_rxpipe_rxvalid,                           Check User Guide for details
		output wire        o_ch3_ux_ock_pma_clk,                           //         .o_ch3_ux_ock_pma_clk,                           Check User Guide for details
		output wire        o_ch3_uxq_lfps_ennt,                            //         .o_ch3_uxq_lfps_ennt,                            Check User Guide for details
		output wire [1:0]  o_ch3_uxq_pcie_l1ctrla,                         //         .o_ch3_uxq_pcie_l1ctrla,                         Check User Guide for details
		output wire        o_ch3_uxq_pma_cmn_ctrl,                         //         .o_ch3_uxq_pma_cmn_ctrl,                         Check User Guide for details
		output wire        o_ch3_uxq_pma_ctrl,                             //         .o_ch3_uxq_pma_ctrl,                             Check User Guide for details
		output wire        o_ch3_uxq_rst_pcs_rx_b_a,                       //         .o_ch3_uxq_rst_pcs_rx_b_a,                       Check User Guide for details
		output wire        o_ch3_uxq_rst_pcs_tx_b_a,                       //         .o_ch3_uxq_rst_pcs_tx_b_a,                       Check User Guide for details
		output wire        o_ch3_uxq_rxeiosdetectstata,                    //         .o_ch3_uxq_rxeiosdetectstata,                    Check User Guide for details
		output wire [2:0]  o_ch3_uxq_rxeq_precal_code_selnt,               //         .o_ch3_uxq_rxeq_precal_code_selnt,               Check User Guide for details
		output wire        o_ch3_uxq_rxeq_starta,                          //         .o_ch3_uxq_rxeq_starta,                          Check User Guide for details
		output wire        o_ch3_uxq_rxeq_static_ena,                      //         .o_ch3_uxq_rxeq_static_ena,                      Check User Guide for details
		output wire        o_ch3_uxq_rxmargin_direction_nt,                //         .o_ch3_uxq_rxmargin_direction_nt,                Check User Guide for details
		output wire        o_ch3_uxq_rxmargin_mode_nt,                     //         .o_ch3_uxq_rxmargin_mode_nt,                     Check User Guide for details
		output wire        o_ch3_uxq_rxmargin_offset_change_a,             //         .o_ch3_uxq_rxmargin_offset_change_a,             Check User Guide for details
		output wire [6:0]  o_ch3_uxq_rxmargin_offset_nt,                   //         .o_ch3_uxq_rxmargin_offset_nt,                   Check User Guide for details
		output wire        o_ch3_uxq_rxmargin_start_a,                     //         .o_ch3_uxq_rxmargin_start_a,                     Check User Guide for details
		output wire [2:0]  o_ch3_uxq_rxpstate,                             //         .o_ch3_uxq_rxpstate,                             Check User Guide for details
		output wire [3:0]  o_ch3_uxq_rxrate,                               //         .o_ch3_uxq_rxrate,                               Check User Guide for details
		output wire        o_ch3_uxq_rxterm_hiz_ena,                       //         .o_ch3_uxq_rxterm_hiz_ena,                       Check User Guide for details
		output wire [2:0]  o_ch3_uxq_rxwidth,                              //         .o_ch3_uxq_rxwidth,                              Check User Guide for details
		output wire        o_ch3_uxq_tstbus_lane,                          //         .o_ch3_uxq_tstbus_lane,                          Check User Guide for details
		output wire        o_ch3_uxq_txbeacona,                            //         .o_ch3_uxq_txbeacona,                            Check User Guide for details
		output wire [2:0]  o_ch3_uxq_txclkdivrate,                         //         .o_ch3_uxq_txclkdivrate,                         Check User Guide for details
		output wire        o_ch3_uxq_txdetectrx_reqa,                      //         .o_ch3_uxq_txdetectrx_reqa,                      Check User Guide for details
		output wire [5:0]  o_ch3_uxq_txdrv_levn,                           //         .o_ch3_uxq_txdrv_levn,                           Check User Guide for details
		output wire [4:0]  o_ch3_uxq_txdrv_levnm1,                         //         .o_ch3_uxq_txdrv_levnm1,                         Check User Guide for details
		output wire [2:0]  o_ch3_uxq_txdrv_levnm2,                         //         .o_ch3_uxq_txdrv_levnm2,                         Check User Guide for details
		output wire [4:0]  o_ch3_uxq_txdrv_levnp1,                         //         .o_ch3_uxq_txdrv_levnp1,                         Check User Guide for details
		output wire [3:0]  o_ch3_uxq_txdrv_slew,                           //         .o_ch3_uxq_txdrv_slew,                           Check User Guide for details
		output wire [3:0]  o_ch3_uxq_txelecidle,                           //         .o_ch3_uxq_txelecidle,                           Check User Guide for details
		output wire [2:0]  o_ch3_uxq_txpstate,                             //         .o_ch3_uxq_txpstate,                             Check User Guide for details
		output wire [3:0]  o_ch3_uxq_txrate,                               //         .o_ch3_uxq_txrate,                               Check User Guide for details
		output wire [2:0]  o_ch3_uxq_txwidth,                              //         .o_ch3_uxq_txwidth,                              Check User Guide for details
		output wire [39:0] o_ch3_uxq_txword                                //         .o_ch3_uxq_txword,                               Check User Guide for details
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (sris_enable != "SRIS_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sris_enable_check ( .error(1'b1) );
		end
		if (pcie_pcs_mode != "PCIE_PCS_MODE_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pcie_pcs_mode_check ( .error(1'b1) );
		end
		if (pclk_clk_hz != 32'b00111011100110101100101000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pclk_clk_hz_check ( .error(1'b1) );
		end
		if (num_of_lanes != 4)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					num_of_lanes_check ( .error(1'b1) );
		end
	endgenerate

	system_intel_pcie_gts_0_pipe_hal_2100_g57zsoa #(
		.sris_enable   ("SRIS_ENABLE_DISABLED"),
		.pcie_pcs_mode ("PCIE_PCS_MODE_PCIE"),
		.pclk_clk_hz   (32'b00111011100110101100101000000000),
		.num_of_lanes  (4)
	) pcie_pipe_hal_top (
		.i_ch0_lavmm_pcie_addr                          (i_ch0_lavmm_pcie_addr),                          //   input,  width = 17, pipe_hal.i_ch0_lavmm_pcie_addr
		.i_ch0_lavmm_pcie_be                            (i_ch0_lavmm_pcie_be),                            //   input,   width = 4,         .i_ch0_lavmm_pcie_be
		.i_ch0_lavmm_pcie_clk                           (i_ch0_lavmm_pcie_clk),                           //   input,   width = 1,         .i_ch0_lavmm_pcie_clk
		.i_ch0_lavmm_pcie_read                          (i_ch0_lavmm_pcie_read),                          //   input,   width = 1,         .i_ch0_lavmm_pcie_read
		.i_ch0_lavmm_pcie_rstn                          (i_ch0_lavmm_pcie_rstn),                          //   input,   width = 1,         .i_ch0_lavmm_pcie_rstn
		.i_ch0_lavmm_pcie_wdata                         (i_ch0_lavmm_pcie_wdata),                         //   input,  width = 32,         .i_ch0_lavmm_pcie_wdata
		.i_ch0_lavmm_pcie_write                         (i_ch0_lavmm_pcie_write),                         //   input,   width = 1,         .i_ch0_lavmm_pcie_write
		.i_ch0_pcie_rxword_clk                          (i_ch0_pcie_rxword_clk),                          //   input,   width = 1,         .i_ch0_pcie_rxword_clk
		.i_ch0_pcie_txword_clk                          (i_ch0_pcie_txword_clk),                          //   input,   width = 1,         .i_ch0_pcie_txword_clk
		.i_ch0_pcs_pclk                                 (i_ch0_pcs_pclk),                                 //   input,   width = 1,         .i_ch0_pcs_pclk
		.i_ch0_pcs_pipe_rstn                            (i_ch0_pcs_pipe_rstn),                            //   input,   width = 1,         .i_ch0_pcs_pipe_rstn
		.i_ch0_txpipe_asyncpowerchangeack               (i_ch0_txpipe_asyncpowerchangeack),               //   input,   width = 1,         .i_ch0_txpipe_asyncpowerchangeack
		.i_ch0_txpipe_blockaligncontrol                 (i_ch0_txpipe_blockaligncontrol),                 //   input,   width = 1,         .i_ch0_txpipe_blockaligncontrol
		.i_ch0_txpipe_cfg_hw_auto_sp_dis                (i_ch0_txpipe_cfg_hw_auto_sp_dis),                //   input,   width = 1,         .i_ch0_txpipe_cfg_hw_auto_sp_dis
		.i_ch0_txpipe_dirchange                         (i_ch0_txpipe_dirchange),                         //   input,   width = 1,         .i_ch0_txpipe_dirchange
		.i_ch0_txpipe_ebuf_mode                         (i_ch0_txpipe_ebuf_mode),                         //   input,   width = 1,         .i_ch0_txpipe_ebuf_mode
		.i_ch0_txpipe_encodedecodebypass                (i_ch0_txpipe_encodedecodebypass),                //   input,   width = 1,         .i_ch0_txpipe_encodedecodebypass
		.i_ch0_txpipe_fs                                (i_ch0_txpipe_fs),                                //   input,   width = 6,         .i_ch0_txpipe_fs
		.i_ch0_txpipe_getlocalpresetcoefficients        (i_ch0_txpipe_getlocalpresetcoefficients),        //   input,   width = 1,         .i_ch0_txpipe_getlocalpresetcoefficients
		.i_ch0_txpipe_invalidrequest                    (i_ch0_txpipe_invalidrequest),                    //   input,   width = 1,         .i_ch0_txpipe_invalidrequest
		.i_ch0_txpipe_lf                                (i_ch0_txpipe_lf),                                //   input,   width = 6,         .i_ch0_txpipe_lf
		.i_ch0_txpipe_localpresetindex                  (i_ch0_txpipe_localpresetindex),                  //   input,   width = 5,         .i_ch0_txpipe_localpresetindex
		.i_ch0_txpipe_lowpin_nt                         (i_ch0_txpipe_lowpin_nt),                         //   input,   width = 1,         .i_ch0_txpipe_lowpin_nt
		.i_ch0_txpipe_m2p_bus                           (i_ch0_txpipe_m2p_bus),                           //   input,   width = 8,         .i_ch0_txpipe_m2p_bus
		.i_ch0_txpipe_pclk_rate                         (i_ch0_txpipe_pclk_rate),                         //   input,   width = 3,         .i_ch0_txpipe_pclk_rate
		.i_ch0_txpipe_pclkchangeack                     (i_ch0_txpipe_pclkchangeack),                     //   input,   width = 1,         .i_ch0_txpipe_pclkchangeack
		.i_ch0_txpipe_phy_mode_nt                       (i_ch0_txpipe_phy_mode_nt),                       //   input,   width = 4,         .i_ch0_txpipe_phy_mode_nt
		.i_ch0_txpipe_powerdown                         (i_ch0_txpipe_powerdown),                         //   input,   width = 4,         .i_ch0_txpipe_powerdown
		.i_ch0_txpipe_rate                              (i_ch0_txpipe_rate),                              //   input,   width = 3,         .i_ch0_txpipe_rate
		.i_ch0_txpipe_rxelecidle_disable_a              (i_ch0_txpipe_rxelecidle_disable_a),              //   input,   width = 1,         .i_ch0_txpipe_rxelecidle_disable_a
		.i_ch0_txpipe_rxeqclr                           (i_ch0_txpipe_rxeqclr),                           //   input,   width = 1,         .i_ch0_txpipe_rxeqclr
		.i_ch0_txpipe_rxeqeval                          (i_ch0_txpipe_rxeqeval),                          //   input,   width = 1,         .i_ch0_txpipe_rxeqeval
		.i_ch0_txpipe_rxeqinprogress                    (i_ch0_txpipe_rxeqinprogress),                    //   input,   width = 1,         .i_ch0_txpipe_rxeqinprogress
		.i_ch0_txpipe_rxeqtraining                      (i_ch0_txpipe_rxeqtraining),                      //   input,   width = 1,         .i_ch0_txpipe_rxeqtraining
		.i_ch0_txpipe_rxpolarity                        (i_ch0_txpipe_rxpolarity),                        //   input,   width = 1,         .i_ch0_txpipe_rxpolarity
		.i_ch0_txpipe_rxpresethint                      (i_ch0_txpipe_rxpresethint),                      //   input,   width = 3,         .i_ch0_txpipe_rxpresethint
		.i_ch0_txpipe_rxstandby                         (i_ch0_txpipe_rxstandby),                         //   input,   width = 1,         .i_ch0_txpipe_rxstandby
		.i_ch0_txpipe_rxtermination                     (i_ch0_txpipe_rxtermination),                     //   input,   width = 1,         .i_ch0_txpipe_rxtermination
		.i_ch0_txpipe_srisenable                        (i_ch0_txpipe_srisenable),                        //   input,   width = 1,         .i_ch0_txpipe_srisenable
		.i_ch0_txpipe_txcmnmode_disable_a               (i_ch0_txpipe_txcmnmode_disable_a),               //   input,   width = 1,         .i_ch0_txpipe_txcmnmode_disable_a
		.i_ch0_txpipe_txcompliance                      (i_ch0_txpipe_txcompliance),                      //   input,   width = 1,         .i_ch0_txpipe_txcompliance
		.i_ch0_txpipe_txdata                            (i_ch0_txpipe_txdata),                            //   input,  width = 40,         .i_ch0_txpipe_txdata
		.i_ch0_txpipe_txdatak                           (i_ch0_txpipe_txdatak),                           //   input,   width = 4,         .i_ch0_txpipe_txdatak
		.i_ch0_txpipe_txdatavalid                       (i_ch0_txpipe_txdatavalid),                       //   input,   width = 1,         .i_ch0_txpipe_txdatavalid
		.i_ch0_txpipe_txdeemph                          (i_ch0_txpipe_txdeemph),                          //   input,  width = 18,         .i_ch0_txpipe_txdeemph
		.i_ch0_txpipe_txdtctrx_lb                       (i_ch0_txpipe_txdtctrx_lb),                       //   input,   width = 1,         .i_ch0_txpipe_txdtctrx_lb
		.i_ch0_txpipe_txelecidle                        (i_ch0_txpipe_txelecidle),                        //   input,   width = 1,         .i_ch0_txpipe_txelecidle
		.i_ch0_txpipe_txmargin                          (i_ch0_txpipe_txmargin),                          //   input,   width = 3,         .i_ch0_txpipe_txmargin
		.i_ch0_txpipe_txoneszeros                       (i_ch0_txpipe_txoneszeros),                       //   input,   width = 1,         .i_ch0_txpipe_txoneszeros
		.i_ch0_txpipe_txstartblock                      (i_ch0_txpipe_txstartblock),                      //   input,   width = 1,         .i_ch0_txpipe_txstartblock
		.i_ch0_txpipe_txswing                           (i_ch0_txpipe_txswing),                           //   input,   width = 1,         .i_ch0_txpipe_txswing
		.i_ch0_txpipe_txsyncheader                      (i_ch0_txpipe_txsyncheader),                      //   input,   width = 4,         .i_ch0_txpipe_txsyncheader
		.i_ch0_txpipe_width                             (i_ch0_txpipe_width),                             //   input,   width = 3,         .i_ch0_txpipe_width
		.i_ch0_uxq_rxcdrlock2dataa                      (i_ch0_uxq_rxcdrlock2dataa),                      //   input,   width = 1,         .i_ch0_uxq_rxcdrlock2dataa
		.i_ch0_uxq_rxeq_best_eye_vala                   (i_ch0_uxq_rxeq_best_eye_vala),                   //   input,  width = 14,         .i_ch0_uxq_rxeq_best_eye_vala
		.i_ch0_uxq_rxeq_donea                           (i_ch0_uxq_rxeq_donea),                           //   input,   width = 1,         .i_ch0_uxq_rxeq_donea
		.i_ch0_uxq_rxmargin_nacka                       (i_ch0_uxq_rxmargin_nacka),                       //   input,   width = 1,         .i_ch0_uxq_rxmargin_nacka
		.i_ch0_uxq_rxmargin_status_gray_a               (i_ch0_uxq_rxmargin_status_gray_a),               //   input,   width = 2,         .i_ch0_uxq_rxmargin_status_gray_a
		.i_ch0_uxq_rxmargin_statusa                     (i_ch0_uxq_rxmargin_statusa),                     //   input,   width = 1,         .i_ch0_uxq_rxmargin_statusa
		.i_ch0_uxq_rxsignaldetect_lfpsa                 (i_ch0_uxq_rxsignaldetect_lfpsa),                 //   input,   width = 1,         .i_ch0_uxq_rxsignaldetect_lfpsa
		.i_ch0_uxq_rxsignaldetecta                      (i_ch0_uxq_rxsignaldetecta),                      //   input,   width = 1,         .i_ch0_uxq_rxsignaldetecta
		.i_ch0_uxq_rxstatusa                            (i_ch0_uxq_rxstatusa),                            //   input,   width = 1,         .i_ch0_uxq_rxstatusa
		.i_ch0_uxq_rxword                               (i_ch0_uxq_rxword),                               //   input,  width = 40,         .i_ch0_uxq_rxword
		.i_ch0_uxq_synthlcfast_postdiv                  (i_ch0_uxq_synthlcfast_postdiv),                  //   input,   width = 1,         .i_ch0_uxq_synthlcfast_postdiv
		.i_ch0_uxq_synthlcmed_postdiv                   (i_ch0_uxq_synthlcmed_postdiv),                   //   input,   width = 1,         .i_ch0_uxq_synthlcmed_postdiv
		.i_ch0_uxq_synthlcslow_postdiv                  (i_ch0_uxq_synthlcslow_postdiv),                  //   input,   width = 1,         .i_ch0_uxq_synthlcslow_postdiv
		.i_ch0_uxq_txdetectrx_acka                      (i_ch0_uxq_txdetectrx_acka),                      //   input,   width = 1,         .i_ch0_uxq_txdetectrx_acka
		.i_ch0_uxq_txdetectrx_statct                    (i_ch0_uxq_txdetectrx_statct),                    //   input,   width = 1,         .i_ch0_uxq_txdetectrx_statct
		.i_ch0_uxq_txstatusa                            (i_ch0_uxq_txstatusa),                            //   input,   width = 1,         .i_ch0_uxq_txstatusa
		.o_ch0_lavmm_pcie_rdata                         (o_ch0_lavmm_pcie_rdata),                         //  output,  width = 32,         .o_ch0_lavmm_pcie_rdata
		.o_ch0_lavmm_pcie_rdata_valid                   (o_ch0_lavmm_pcie_rdata_valid),                   //  output,   width = 1,         .o_ch0_lavmm_pcie_rdata_valid
		.o_ch0_lavmm_pcie_waitreq                       (o_ch0_lavmm_pcie_waitreq),                       //  output,   width = 1,         .o_ch0_lavmm_pcie_waitreq
		.o_ch0_pcs_pclk                                 (o_ch0_pcs_pclk),                                 //  output,   width = 1,         .o_ch0_pcs_pclk
		.o_ch0_pcs_pipe_rstn                            (o_ch0_pcs_pipe_rstn),                            //  output,   width = 1,         .o_ch0_pcs_pipe_rstn
		.o_ch0_rxpipe_dirfeedback                       (o_ch0_rxpipe_dirfeedback),                       //  output,   width = 6,         .o_ch0_rxpipe_dirfeedback
		.o_ch0_rxpipe_linkevaluationfeedbackfiguremerit (o_ch0_rxpipe_linkevaluationfeedbackfiguremerit), //  output,   width = 8,         .o_ch0_rxpipe_linkevaluationfeedbackfiguremerit
		.o_ch0_rxpipe_localfs                           (o_ch0_rxpipe_localfs),                           //  output,   width = 6,         .o_ch0_rxpipe_localfs
		.o_ch0_rxpipe_locallf                           (o_ch0_rxpipe_locallf),                           //  output,   width = 6,         .o_ch0_rxpipe_locallf
		.o_ch0_rxpipe_localtxcoefficientsvalid          (o_ch0_rxpipe_localtxcoefficientsvalid),          //  output,   width = 1,         .o_ch0_rxpipe_localtxcoefficientsvalid
		.o_ch0_rxpipe_localtxpresetcoefficients         (o_ch0_rxpipe_localtxpresetcoefficients),         //  output,  width = 18,         .o_ch0_rxpipe_localtxpresetcoefficients
		.o_ch0_rxpipe_p2m_bus                           (o_ch0_rxpipe_p2m_bus),                           //  output,   width = 8,         .o_ch0_rxpipe_p2m_bus
		.o_ch0_rxpipe_pclkchangeok                      (o_ch0_rxpipe_pclkchangeok),                      //  output,   width = 1,         .o_ch0_rxpipe_pclkchangeok
		.o_ch0_rxpipe_phystatus                         (o_ch0_rxpipe_phystatus),                         //  output,   width = 1,         .o_ch0_rxpipe_phystatus
		.o_ch0_rxpipe_rxdata                            (o_ch0_rxpipe_rxdata),                            //  output,  width = 40,         .o_ch0_rxpipe_rxdata
		.o_ch0_rxpipe_rxdatak                           (o_ch0_rxpipe_rxdatak),                           //  output,   width = 4,         .o_ch0_rxpipe_rxdatak
		.o_ch0_rxpipe_rxdatavalid                       (o_ch0_rxpipe_rxdatavalid),                       //  output,   width = 1,         .o_ch0_rxpipe_rxdatavalid
		.o_ch0_rxpipe_rxelecidlea                       (o_ch0_rxpipe_rxelecidlea),                       //  output,   width = 1,         .o_ch0_rxpipe_rxelecidlea
		.o_ch0_rxpipe_rxstandbystatus                   (o_ch0_rxpipe_rxstandbystatus),                   //  output,   width = 1,         .o_ch0_rxpipe_rxstandbystatus
		.o_ch0_rxpipe_rxstartblock                      (o_ch0_rxpipe_rxstartblock),                      //  output,   width = 1,         .o_ch0_rxpipe_rxstartblock
		.o_ch0_rxpipe_rxstatus                          (o_ch0_rxpipe_rxstatus),                          //  output,   width = 3,         .o_ch0_rxpipe_rxstatus
		.o_ch0_rxpipe_rxsyncheader                      (o_ch0_rxpipe_rxsyncheader),                      //  output,   width = 4,         .o_ch0_rxpipe_rxsyncheader
		.o_ch0_rxpipe_rxvalid                           (o_ch0_rxpipe_rxvalid),                           //  output,   width = 1,         .o_ch0_rxpipe_rxvalid
		.o_ch0_ux_ock_pma_clk                           (o_ch0_ux_ock_pma_clk),                           //  output,   width = 1,         .o_ch0_ux_ock_pma_clk
		.o_ch0_uxq_lfps_ennt                            (o_ch0_uxq_lfps_ennt),                            //  output,   width = 1,         .o_ch0_uxq_lfps_ennt
		.o_ch0_uxq_pcie_l1ctrla                         (o_ch0_uxq_pcie_l1ctrla),                         //  output,   width = 2,         .o_ch0_uxq_pcie_l1ctrla
		.o_ch0_uxq_pma_cmn_ctrl                         (o_ch0_uxq_pma_cmn_ctrl),                         //  output,   width = 1,         .o_ch0_uxq_pma_cmn_ctrl
		.o_ch0_uxq_pma_ctrl                             (o_ch0_uxq_pma_ctrl),                             //  output,   width = 1,         .o_ch0_uxq_pma_ctrl
		.o_ch0_uxq_rst_pcs_rx_b_a                       (o_ch0_uxq_rst_pcs_rx_b_a),                       //  output,   width = 1,         .o_ch0_uxq_rst_pcs_rx_b_a
		.o_ch0_uxq_rst_pcs_tx_b_a                       (o_ch0_uxq_rst_pcs_tx_b_a),                       //  output,   width = 1,         .o_ch0_uxq_rst_pcs_tx_b_a
		.o_ch0_uxq_rxeiosdetectstata                    (o_ch0_uxq_rxeiosdetectstata),                    //  output,   width = 1,         .o_ch0_uxq_rxeiosdetectstata
		.o_ch0_uxq_rxeq_precal_code_selnt               (o_ch0_uxq_rxeq_precal_code_selnt),               //  output,   width = 3,         .o_ch0_uxq_rxeq_precal_code_selnt
		.o_ch0_uxq_rxeq_starta                          (o_ch0_uxq_rxeq_starta),                          //  output,   width = 1,         .o_ch0_uxq_rxeq_starta
		.o_ch0_uxq_rxeq_static_ena                      (o_ch0_uxq_rxeq_static_ena),                      //  output,   width = 1,         .o_ch0_uxq_rxeq_static_ena
		.o_ch0_uxq_rxmargin_direction_nt                (o_ch0_uxq_rxmargin_direction_nt),                //  output,   width = 1,         .o_ch0_uxq_rxmargin_direction_nt
		.o_ch0_uxq_rxmargin_mode_nt                     (o_ch0_uxq_rxmargin_mode_nt),                     //  output,   width = 1,         .o_ch0_uxq_rxmargin_mode_nt
		.o_ch0_uxq_rxmargin_offset_change_a             (o_ch0_uxq_rxmargin_offset_change_a),             //  output,   width = 1,         .o_ch0_uxq_rxmargin_offset_change_a
		.o_ch0_uxq_rxmargin_offset_nt                   (o_ch0_uxq_rxmargin_offset_nt),                   //  output,   width = 7,         .o_ch0_uxq_rxmargin_offset_nt
		.o_ch0_uxq_rxmargin_start_a                     (o_ch0_uxq_rxmargin_start_a),                     //  output,   width = 1,         .o_ch0_uxq_rxmargin_start_a
		.o_ch0_uxq_rxpstate                             (o_ch0_uxq_rxpstate),                             //  output,   width = 3,         .o_ch0_uxq_rxpstate
		.o_ch0_uxq_rxrate                               (o_ch0_uxq_rxrate),                               //  output,   width = 4,         .o_ch0_uxq_rxrate
		.o_ch0_uxq_rxterm_hiz_ena                       (o_ch0_uxq_rxterm_hiz_ena),                       //  output,   width = 1,         .o_ch0_uxq_rxterm_hiz_ena
		.o_ch0_uxq_rxwidth                              (o_ch0_uxq_rxwidth),                              //  output,   width = 3,         .o_ch0_uxq_rxwidth
		.o_ch0_uxq_tstbus_lane                          (o_ch0_uxq_tstbus_lane),                          //  output,   width = 1,         .o_ch0_uxq_tstbus_lane
		.o_ch0_uxq_txbeacona                            (o_ch0_uxq_txbeacona),                            //  output,   width = 1,         .o_ch0_uxq_txbeacona
		.o_ch0_uxq_txclkdivrate                         (o_ch0_uxq_txclkdivrate),                         //  output,   width = 3,         .o_ch0_uxq_txclkdivrate
		.o_ch0_uxq_txdetectrx_reqa                      (o_ch0_uxq_txdetectrx_reqa),                      //  output,   width = 1,         .o_ch0_uxq_txdetectrx_reqa
		.o_ch0_uxq_txdrv_levn                           (o_ch0_uxq_txdrv_levn),                           //  output,   width = 6,         .o_ch0_uxq_txdrv_levn
		.o_ch0_uxq_txdrv_levnm1                         (o_ch0_uxq_txdrv_levnm1),                         //  output,   width = 5,         .o_ch0_uxq_txdrv_levnm1
		.o_ch0_uxq_txdrv_levnm2                         (o_ch0_uxq_txdrv_levnm2),                         //  output,   width = 3,         .o_ch0_uxq_txdrv_levnm2
		.o_ch0_uxq_txdrv_levnp1                         (o_ch0_uxq_txdrv_levnp1),                         //  output,   width = 5,         .o_ch0_uxq_txdrv_levnp1
		.o_ch0_uxq_txdrv_slew                           (o_ch0_uxq_txdrv_slew),                           //  output,   width = 4,         .o_ch0_uxq_txdrv_slew
		.o_ch0_uxq_txelecidle                           (o_ch0_uxq_txelecidle),                           //  output,   width = 4,         .o_ch0_uxq_txelecidle
		.o_ch0_uxq_txpstate                             (o_ch0_uxq_txpstate),                             //  output,   width = 3,         .o_ch0_uxq_txpstate
		.o_ch0_uxq_txrate                               (o_ch0_uxq_txrate),                               //  output,   width = 4,         .o_ch0_uxq_txrate
		.o_ch0_uxq_txwidth                              (o_ch0_uxq_txwidth),                              //  output,   width = 3,         .o_ch0_uxq_txwidth
		.o_ch0_uxq_txword                               (o_ch0_uxq_txword),                               //  output,  width = 40,         .o_ch0_uxq_txword
		.i_ch1_lavmm_pcie_addr                          (i_ch1_lavmm_pcie_addr),                          //   input,  width = 17,         .i_ch1_lavmm_pcie_addr
		.i_ch1_lavmm_pcie_be                            (i_ch1_lavmm_pcie_be),                            //   input,   width = 4,         .i_ch1_lavmm_pcie_be
		.i_ch1_lavmm_pcie_clk                           (i_ch1_lavmm_pcie_clk),                           //   input,   width = 1,         .i_ch1_lavmm_pcie_clk
		.i_ch1_lavmm_pcie_read                          (i_ch1_lavmm_pcie_read),                          //   input,   width = 1,         .i_ch1_lavmm_pcie_read
		.i_ch1_lavmm_pcie_rstn                          (i_ch1_lavmm_pcie_rstn),                          //   input,   width = 1,         .i_ch1_lavmm_pcie_rstn
		.i_ch1_lavmm_pcie_wdata                         (i_ch1_lavmm_pcie_wdata),                         //   input,  width = 32,         .i_ch1_lavmm_pcie_wdata
		.i_ch1_lavmm_pcie_write                         (i_ch1_lavmm_pcie_write),                         //   input,   width = 1,         .i_ch1_lavmm_pcie_write
		.i_ch1_pcie_rxword_clk                          (i_ch1_pcie_rxword_clk),                          //   input,   width = 1,         .i_ch1_pcie_rxword_clk
		.i_ch1_pcie_txword_clk                          (i_ch1_pcie_txword_clk),                          //   input,   width = 1,         .i_ch1_pcie_txword_clk
		.i_ch1_pcs_pclk                                 (i_ch1_pcs_pclk),                                 //   input,   width = 1,         .i_ch1_pcs_pclk
		.i_ch1_pcs_pipe_rstn                            (i_ch1_pcs_pipe_rstn),                            //   input,   width = 1,         .i_ch1_pcs_pipe_rstn
		.i_ch1_txpipe_asyncpowerchangeack               (i_ch1_txpipe_asyncpowerchangeack),               //   input,   width = 1,         .i_ch1_txpipe_asyncpowerchangeack
		.i_ch1_txpipe_blockaligncontrol                 (i_ch1_txpipe_blockaligncontrol),                 //   input,   width = 1,         .i_ch1_txpipe_blockaligncontrol
		.i_ch1_txpipe_cfg_hw_auto_sp_dis                (i_ch1_txpipe_cfg_hw_auto_sp_dis),                //   input,   width = 1,         .i_ch1_txpipe_cfg_hw_auto_sp_dis
		.i_ch1_txpipe_dirchange                         (i_ch1_txpipe_dirchange),                         //   input,   width = 1,         .i_ch1_txpipe_dirchange
		.i_ch1_txpipe_ebuf_mode                         (i_ch1_txpipe_ebuf_mode),                         //   input,   width = 1,         .i_ch1_txpipe_ebuf_mode
		.i_ch1_txpipe_encodedecodebypass                (i_ch1_txpipe_encodedecodebypass),                //   input,   width = 1,         .i_ch1_txpipe_encodedecodebypass
		.i_ch1_txpipe_fs                                (i_ch1_txpipe_fs),                                //   input,   width = 6,         .i_ch1_txpipe_fs
		.i_ch1_txpipe_getlocalpresetcoefficients        (i_ch1_txpipe_getlocalpresetcoefficients),        //   input,   width = 1,         .i_ch1_txpipe_getlocalpresetcoefficients
		.i_ch1_txpipe_invalidrequest                    (i_ch1_txpipe_invalidrequest),                    //   input,   width = 1,         .i_ch1_txpipe_invalidrequest
		.i_ch1_txpipe_lf                                (i_ch1_txpipe_lf),                                //   input,   width = 6,         .i_ch1_txpipe_lf
		.i_ch1_txpipe_localpresetindex                  (i_ch1_txpipe_localpresetindex),                  //   input,   width = 5,         .i_ch1_txpipe_localpresetindex
		.i_ch1_txpipe_lowpin_nt                         (i_ch1_txpipe_lowpin_nt),                         //   input,   width = 1,         .i_ch1_txpipe_lowpin_nt
		.i_ch1_txpipe_m2p_bus                           (i_ch1_txpipe_m2p_bus),                           //   input,   width = 8,         .i_ch1_txpipe_m2p_bus
		.i_ch1_txpipe_pclk_rate                         (i_ch1_txpipe_pclk_rate),                         //   input,   width = 3,         .i_ch1_txpipe_pclk_rate
		.i_ch1_txpipe_pclkchangeack                     (i_ch1_txpipe_pclkchangeack),                     //   input,   width = 1,         .i_ch1_txpipe_pclkchangeack
		.i_ch1_txpipe_phy_mode_nt                       (i_ch1_txpipe_phy_mode_nt),                       //   input,   width = 4,         .i_ch1_txpipe_phy_mode_nt
		.i_ch1_txpipe_powerdown                         (i_ch1_txpipe_powerdown),                         //   input,   width = 4,         .i_ch1_txpipe_powerdown
		.i_ch1_txpipe_rate                              (i_ch1_txpipe_rate),                              //   input,   width = 3,         .i_ch1_txpipe_rate
		.i_ch1_txpipe_rxelecidle_disable_a              (i_ch1_txpipe_rxelecidle_disable_a),              //   input,   width = 1,         .i_ch1_txpipe_rxelecidle_disable_a
		.i_ch1_txpipe_rxeqclr                           (i_ch1_txpipe_rxeqclr),                           //   input,   width = 1,         .i_ch1_txpipe_rxeqclr
		.i_ch1_txpipe_rxeqeval                          (i_ch1_txpipe_rxeqeval),                          //   input,   width = 1,         .i_ch1_txpipe_rxeqeval
		.i_ch1_txpipe_rxeqinprogress                    (i_ch1_txpipe_rxeqinprogress),                    //   input,   width = 1,         .i_ch1_txpipe_rxeqinprogress
		.i_ch1_txpipe_rxeqtraining                      (i_ch1_txpipe_rxeqtraining),                      //   input,   width = 1,         .i_ch1_txpipe_rxeqtraining
		.i_ch1_txpipe_rxpolarity                        (i_ch1_txpipe_rxpolarity),                        //   input,   width = 1,         .i_ch1_txpipe_rxpolarity
		.i_ch1_txpipe_rxpresethint                      (i_ch1_txpipe_rxpresethint),                      //   input,   width = 3,         .i_ch1_txpipe_rxpresethint
		.i_ch1_txpipe_rxstandby                         (i_ch1_txpipe_rxstandby),                         //   input,   width = 1,         .i_ch1_txpipe_rxstandby
		.i_ch1_txpipe_rxtermination                     (i_ch1_txpipe_rxtermination),                     //   input,   width = 1,         .i_ch1_txpipe_rxtermination
		.i_ch1_txpipe_srisenable                        (i_ch1_txpipe_srisenable),                        //   input,   width = 1,         .i_ch1_txpipe_srisenable
		.i_ch1_txpipe_txcmnmode_disable_a               (i_ch1_txpipe_txcmnmode_disable_a),               //   input,   width = 1,         .i_ch1_txpipe_txcmnmode_disable_a
		.i_ch1_txpipe_txcompliance                      (i_ch1_txpipe_txcompliance),                      //   input,   width = 1,         .i_ch1_txpipe_txcompliance
		.i_ch1_txpipe_txdata                            (i_ch1_txpipe_txdata),                            //   input,  width = 40,         .i_ch1_txpipe_txdata
		.i_ch1_txpipe_txdatak                           (i_ch1_txpipe_txdatak),                           //   input,   width = 4,         .i_ch1_txpipe_txdatak
		.i_ch1_txpipe_txdatavalid                       (i_ch1_txpipe_txdatavalid),                       //   input,   width = 1,         .i_ch1_txpipe_txdatavalid
		.i_ch1_txpipe_txdeemph                          (i_ch1_txpipe_txdeemph),                          //   input,  width = 18,         .i_ch1_txpipe_txdeemph
		.i_ch1_txpipe_txdtctrx_lb                       (i_ch1_txpipe_txdtctrx_lb),                       //   input,   width = 1,         .i_ch1_txpipe_txdtctrx_lb
		.i_ch1_txpipe_txelecidle                        (i_ch1_txpipe_txelecidle),                        //   input,   width = 1,         .i_ch1_txpipe_txelecidle
		.i_ch1_txpipe_txmargin                          (i_ch1_txpipe_txmargin),                          //   input,   width = 3,         .i_ch1_txpipe_txmargin
		.i_ch1_txpipe_txoneszeros                       (i_ch1_txpipe_txoneszeros),                       //   input,   width = 1,         .i_ch1_txpipe_txoneszeros
		.i_ch1_txpipe_txstartblock                      (i_ch1_txpipe_txstartblock),                      //   input,   width = 1,         .i_ch1_txpipe_txstartblock
		.i_ch1_txpipe_txswing                           (i_ch1_txpipe_txswing),                           //   input,   width = 1,         .i_ch1_txpipe_txswing
		.i_ch1_txpipe_txsyncheader                      (i_ch1_txpipe_txsyncheader),                      //   input,   width = 4,         .i_ch1_txpipe_txsyncheader
		.i_ch1_txpipe_width                             (i_ch1_txpipe_width),                             //   input,   width = 3,         .i_ch1_txpipe_width
		.i_ch1_uxq_rxcdrlock2dataa                      (i_ch1_uxq_rxcdrlock2dataa),                      //   input,   width = 1,         .i_ch1_uxq_rxcdrlock2dataa
		.i_ch1_uxq_rxeq_best_eye_vala                   (i_ch1_uxq_rxeq_best_eye_vala),                   //   input,  width = 14,         .i_ch1_uxq_rxeq_best_eye_vala
		.i_ch1_uxq_rxeq_donea                           (i_ch1_uxq_rxeq_donea),                           //   input,   width = 1,         .i_ch1_uxq_rxeq_donea
		.i_ch1_uxq_rxmargin_nacka                       (i_ch1_uxq_rxmargin_nacka),                       //   input,   width = 1,         .i_ch1_uxq_rxmargin_nacka
		.i_ch1_uxq_rxmargin_status_gray_a               (i_ch1_uxq_rxmargin_status_gray_a),               //   input,   width = 2,         .i_ch1_uxq_rxmargin_status_gray_a
		.i_ch1_uxq_rxmargin_statusa                     (i_ch1_uxq_rxmargin_statusa),                     //   input,   width = 1,         .i_ch1_uxq_rxmargin_statusa
		.i_ch1_uxq_rxsignaldetect_lfpsa                 (i_ch1_uxq_rxsignaldetect_lfpsa),                 //   input,   width = 1,         .i_ch1_uxq_rxsignaldetect_lfpsa
		.i_ch1_uxq_rxsignaldetecta                      (i_ch1_uxq_rxsignaldetecta),                      //   input,   width = 1,         .i_ch1_uxq_rxsignaldetecta
		.i_ch1_uxq_rxstatusa                            (i_ch1_uxq_rxstatusa),                            //   input,   width = 1,         .i_ch1_uxq_rxstatusa
		.i_ch1_uxq_rxword                               (i_ch1_uxq_rxword),                               //   input,  width = 40,         .i_ch1_uxq_rxword
		.i_ch1_uxq_synthlcfast_postdiv                  (i_ch1_uxq_synthlcfast_postdiv),                  //   input,   width = 1,         .i_ch1_uxq_synthlcfast_postdiv
		.i_ch1_uxq_synthlcmed_postdiv                   (i_ch1_uxq_synthlcmed_postdiv),                   //   input,   width = 1,         .i_ch1_uxq_synthlcmed_postdiv
		.i_ch1_uxq_synthlcslow_postdiv                  (i_ch1_uxq_synthlcslow_postdiv),                  //   input,   width = 1,         .i_ch1_uxq_synthlcslow_postdiv
		.i_ch1_uxq_txdetectrx_acka                      (i_ch1_uxq_txdetectrx_acka),                      //   input,   width = 1,         .i_ch1_uxq_txdetectrx_acka
		.i_ch1_uxq_txdetectrx_statct                    (i_ch1_uxq_txdetectrx_statct),                    //   input,   width = 1,         .i_ch1_uxq_txdetectrx_statct
		.i_ch1_uxq_txstatusa                            (i_ch1_uxq_txstatusa),                            //   input,   width = 1,         .i_ch1_uxq_txstatusa
		.o_ch1_lavmm_pcie_rdata                         (o_ch1_lavmm_pcie_rdata),                         //  output,  width = 32,         .o_ch1_lavmm_pcie_rdata
		.o_ch1_lavmm_pcie_rdata_valid                   (o_ch1_lavmm_pcie_rdata_valid),                   //  output,   width = 1,         .o_ch1_lavmm_pcie_rdata_valid
		.o_ch1_lavmm_pcie_waitreq                       (o_ch1_lavmm_pcie_waitreq),                       //  output,   width = 1,         .o_ch1_lavmm_pcie_waitreq
		.o_ch1_pcs_pclk                                 (o_ch1_pcs_pclk),                                 //  output,   width = 1,         .o_ch1_pcs_pclk
		.o_ch1_pcs_pipe_rstn                            (o_ch1_pcs_pipe_rstn),                            //  output,   width = 1,         .o_ch1_pcs_pipe_rstn
		.o_ch1_rxpipe_dirfeedback                       (o_ch1_rxpipe_dirfeedback),                       //  output,   width = 6,         .o_ch1_rxpipe_dirfeedback
		.o_ch1_rxpipe_linkevaluationfeedbackfiguremerit (o_ch1_rxpipe_linkevaluationfeedbackfiguremerit), //  output,   width = 8,         .o_ch1_rxpipe_linkevaluationfeedbackfiguremerit
		.o_ch1_rxpipe_localfs                           (o_ch1_rxpipe_localfs),                           //  output,   width = 6,         .o_ch1_rxpipe_localfs
		.o_ch1_rxpipe_locallf                           (o_ch1_rxpipe_locallf),                           //  output,   width = 6,         .o_ch1_rxpipe_locallf
		.o_ch1_rxpipe_localtxcoefficientsvalid          (o_ch1_rxpipe_localtxcoefficientsvalid),          //  output,   width = 1,         .o_ch1_rxpipe_localtxcoefficientsvalid
		.o_ch1_rxpipe_localtxpresetcoefficients         (o_ch1_rxpipe_localtxpresetcoefficients),         //  output,  width = 18,         .o_ch1_rxpipe_localtxpresetcoefficients
		.o_ch1_rxpipe_p2m_bus                           (o_ch1_rxpipe_p2m_bus),                           //  output,   width = 8,         .o_ch1_rxpipe_p2m_bus
		.o_ch1_rxpipe_pclkchangeok                      (o_ch1_rxpipe_pclkchangeok),                      //  output,   width = 1,         .o_ch1_rxpipe_pclkchangeok
		.o_ch1_rxpipe_phystatus                         (o_ch1_rxpipe_phystatus),                         //  output,   width = 1,         .o_ch1_rxpipe_phystatus
		.o_ch1_rxpipe_rxdata                            (o_ch1_rxpipe_rxdata),                            //  output,  width = 40,         .o_ch1_rxpipe_rxdata
		.o_ch1_rxpipe_rxdatak                           (o_ch1_rxpipe_rxdatak),                           //  output,   width = 4,         .o_ch1_rxpipe_rxdatak
		.o_ch1_rxpipe_rxdatavalid                       (o_ch1_rxpipe_rxdatavalid),                       //  output,   width = 1,         .o_ch1_rxpipe_rxdatavalid
		.o_ch1_rxpipe_rxelecidlea                       (o_ch1_rxpipe_rxelecidlea),                       //  output,   width = 1,         .o_ch1_rxpipe_rxelecidlea
		.o_ch1_rxpipe_rxstandbystatus                   (o_ch1_rxpipe_rxstandbystatus),                   //  output,   width = 1,         .o_ch1_rxpipe_rxstandbystatus
		.o_ch1_rxpipe_rxstartblock                      (o_ch1_rxpipe_rxstartblock),                      //  output,   width = 1,         .o_ch1_rxpipe_rxstartblock
		.o_ch1_rxpipe_rxstatus                          (o_ch1_rxpipe_rxstatus),                          //  output,   width = 3,         .o_ch1_rxpipe_rxstatus
		.o_ch1_rxpipe_rxsyncheader                      (o_ch1_rxpipe_rxsyncheader),                      //  output,   width = 4,         .o_ch1_rxpipe_rxsyncheader
		.o_ch1_rxpipe_rxvalid                           (o_ch1_rxpipe_rxvalid),                           //  output,   width = 1,         .o_ch1_rxpipe_rxvalid
		.o_ch1_ux_ock_pma_clk                           (o_ch1_ux_ock_pma_clk),                           //  output,   width = 1,         .o_ch1_ux_ock_pma_clk
		.o_ch1_uxq_lfps_ennt                            (o_ch1_uxq_lfps_ennt),                            //  output,   width = 1,         .o_ch1_uxq_lfps_ennt
		.o_ch1_uxq_pcie_l1ctrla                         (o_ch1_uxq_pcie_l1ctrla),                         //  output,   width = 2,         .o_ch1_uxq_pcie_l1ctrla
		.o_ch1_uxq_pma_cmn_ctrl                         (o_ch1_uxq_pma_cmn_ctrl),                         //  output,   width = 1,         .o_ch1_uxq_pma_cmn_ctrl
		.o_ch1_uxq_pma_ctrl                             (o_ch1_uxq_pma_ctrl),                             //  output,   width = 1,         .o_ch1_uxq_pma_ctrl
		.o_ch1_uxq_rst_pcs_rx_b_a                       (o_ch1_uxq_rst_pcs_rx_b_a),                       //  output,   width = 1,         .o_ch1_uxq_rst_pcs_rx_b_a
		.o_ch1_uxq_rst_pcs_tx_b_a                       (o_ch1_uxq_rst_pcs_tx_b_a),                       //  output,   width = 1,         .o_ch1_uxq_rst_pcs_tx_b_a
		.o_ch1_uxq_rxeiosdetectstata                    (o_ch1_uxq_rxeiosdetectstata),                    //  output,   width = 1,         .o_ch1_uxq_rxeiosdetectstata
		.o_ch1_uxq_rxeq_precal_code_selnt               (o_ch1_uxq_rxeq_precal_code_selnt),               //  output,   width = 3,         .o_ch1_uxq_rxeq_precal_code_selnt
		.o_ch1_uxq_rxeq_starta                          (o_ch1_uxq_rxeq_starta),                          //  output,   width = 1,         .o_ch1_uxq_rxeq_starta
		.o_ch1_uxq_rxeq_static_ena                      (o_ch1_uxq_rxeq_static_ena),                      //  output,   width = 1,         .o_ch1_uxq_rxeq_static_ena
		.o_ch1_uxq_rxmargin_direction_nt                (o_ch1_uxq_rxmargin_direction_nt),                //  output,   width = 1,         .o_ch1_uxq_rxmargin_direction_nt
		.o_ch1_uxq_rxmargin_mode_nt                     (o_ch1_uxq_rxmargin_mode_nt),                     //  output,   width = 1,         .o_ch1_uxq_rxmargin_mode_nt
		.o_ch1_uxq_rxmargin_offset_change_a             (o_ch1_uxq_rxmargin_offset_change_a),             //  output,   width = 1,         .o_ch1_uxq_rxmargin_offset_change_a
		.o_ch1_uxq_rxmargin_offset_nt                   (o_ch1_uxq_rxmargin_offset_nt),                   //  output,   width = 7,         .o_ch1_uxq_rxmargin_offset_nt
		.o_ch1_uxq_rxmargin_start_a                     (o_ch1_uxq_rxmargin_start_a),                     //  output,   width = 1,         .o_ch1_uxq_rxmargin_start_a
		.o_ch1_uxq_rxpstate                             (o_ch1_uxq_rxpstate),                             //  output,   width = 3,         .o_ch1_uxq_rxpstate
		.o_ch1_uxq_rxrate                               (o_ch1_uxq_rxrate),                               //  output,   width = 4,         .o_ch1_uxq_rxrate
		.o_ch1_uxq_rxterm_hiz_ena                       (o_ch1_uxq_rxterm_hiz_ena),                       //  output,   width = 1,         .o_ch1_uxq_rxterm_hiz_ena
		.o_ch1_uxq_rxwidth                              (o_ch1_uxq_rxwidth),                              //  output,   width = 3,         .o_ch1_uxq_rxwidth
		.o_ch1_uxq_tstbus_lane                          (o_ch1_uxq_tstbus_lane),                          //  output,   width = 1,         .o_ch1_uxq_tstbus_lane
		.o_ch1_uxq_txbeacona                            (o_ch1_uxq_txbeacona),                            //  output,   width = 1,         .o_ch1_uxq_txbeacona
		.o_ch1_uxq_txclkdivrate                         (o_ch1_uxq_txclkdivrate),                         //  output,   width = 3,         .o_ch1_uxq_txclkdivrate
		.o_ch1_uxq_txdetectrx_reqa                      (o_ch1_uxq_txdetectrx_reqa),                      //  output,   width = 1,         .o_ch1_uxq_txdetectrx_reqa
		.o_ch1_uxq_txdrv_levn                           (o_ch1_uxq_txdrv_levn),                           //  output,   width = 6,         .o_ch1_uxq_txdrv_levn
		.o_ch1_uxq_txdrv_levnm1                         (o_ch1_uxq_txdrv_levnm1),                         //  output,   width = 5,         .o_ch1_uxq_txdrv_levnm1
		.o_ch1_uxq_txdrv_levnm2                         (o_ch1_uxq_txdrv_levnm2),                         //  output,   width = 3,         .o_ch1_uxq_txdrv_levnm2
		.o_ch1_uxq_txdrv_levnp1                         (o_ch1_uxq_txdrv_levnp1),                         //  output,   width = 5,         .o_ch1_uxq_txdrv_levnp1
		.o_ch1_uxq_txdrv_slew                           (o_ch1_uxq_txdrv_slew),                           //  output,   width = 4,         .o_ch1_uxq_txdrv_slew
		.o_ch1_uxq_txelecidle                           (o_ch1_uxq_txelecidle),                           //  output,   width = 4,         .o_ch1_uxq_txelecidle
		.o_ch1_uxq_txpstate                             (o_ch1_uxq_txpstate),                             //  output,   width = 3,         .o_ch1_uxq_txpstate
		.o_ch1_uxq_txrate                               (o_ch1_uxq_txrate),                               //  output,   width = 4,         .o_ch1_uxq_txrate
		.o_ch1_uxq_txwidth                              (o_ch1_uxq_txwidth),                              //  output,   width = 3,         .o_ch1_uxq_txwidth
		.o_ch1_uxq_txword                               (o_ch1_uxq_txword),                               //  output,  width = 40,         .o_ch1_uxq_txword
		.i_ch2_lavmm_pcie_addr                          (i_ch2_lavmm_pcie_addr),                          //   input,  width = 17,         .i_ch2_lavmm_pcie_addr
		.i_ch2_lavmm_pcie_be                            (i_ch2_lavmm_pcie_be),                            //   input,   width = 4,         .i_ch2_lavmm_pcie_be
		.i_ch2_lavmm_pcie_clk                           (i_ch2_lavmm_pcie_clk),                           //   input,   width = 1,         .i_ch2_lavmm_pcie_clk
		.i_ch2_lavmm_pcie_read                          (i_ch2_lavmm_pcie_read),                          //   input,   width = 1,         .i_ch2_lavmm_pcie_read
		.i_ch2_lavmm_pcie_rstn                          (i_ch2_lavmm_pcie_rstn),                          //   input,   width = 1,         .i_ch2_lavmm_pcie_rstn
		.i_ch2_lavmm_pcie_wdata                         (i_ch2_lavmm_pcie_wdata),                         //   input,  width = 32,         .i_ch2_lavmm_pcie_wdata
		.i_ch2_lavmm_pcie_write                         (i_ch2_lavmm_pcie_write),                         //   input,   width = 1,         .i_ch2_lavmm_pcie_write
		.i_ch2_pcie_rxword_clk                          (i_ch2_pcie_rxword_clk),                          //   input,   width = 1,         .i_ch2_pcie_rxword_clk
		.i_ch2_pcie_txword_clk                          (i_ch2_pcie_txword_clk),                          //   input,   width = 1,         .i_ch2_pcie_txword_clk
		.i_ch2_pcs_pclk                                 (i_ch2_pcs_pclk),                                 //   input,   width = 1,         .i_ch2_pcs_pclk
		.i_ch2_pcs_pipe_rstn                            (i_ch2_pcs_pipe_rstn),                            //   input,   width = 1,         .i_ch2_pcs_pipe_rstn
		.i_ch2_txpipe_asyncpowerchangeack               (i_ch2_txpipe_asyncpowerchangeack),               //   input,   width = 1,         .i_ch2_txpipe_asyncpowerchangeack
		.i_ch2_txpipe_blockaligncontrol                 (i_ch2_txpipe_blockaligncontrol),                 //   input,   width = 1,         .i_ch2_txpipe_blockaligncontrol
		.i_ch2_txpipe_cfg_hw_auto_sp_dis                (i_ch2_txpipe_cfg_hw_auto_sp_dis),                //   input,   width = 1,         .i_ch2_txpipe_cfg_hw_auto_sp_dis
		.i_ch2_txpipe_dirchange                         (i_ch2_txpipe_dirchange),                         //   input,   width = 1,         .i_ch2_txpipe_dirchange
		.i_ch2_txpipe_ebuf_mode                         (i_ch2_txpipe_ebuf_mode),                         //   input,   width = 1,         .i_ch2_txpipe_ebuf_mode
		.i_ch2_txpipe_encodedecodebypass                (i_ch2_txpipe_encodedecodebypass),                //   input,   width = 1,         .i_ch2_txpipe_encodedecodebypass
		.i_ch2_txpipe_fs                                (i_ch2_txpipe_fs),                                //   input,   width = 6,         .i_ch2_txpipe_fs
		.i_ch2_txpipe_getlocalpresetcoefficients        (i_ch2_txpipe_getlocalpresetcoefficients),        //   input,   width = 1,         .i_ch2_txpipe_getlocalpresetcoefficients
		.i_ch2_txpipe_invalidrequest                    (i_ch2_txpipe_invalidrequest),                    //   input,   width = 1,         .i_ch2_txpipe_invalidrequest
		.i_ch2_txpipe_lf                                (i_ch2_txpipe_lf),                                //   input,   width = 6,         .i_ch2_txpipe_lf
		.i_ch2_txpipe_localpresetindex                  (i_ch2_txpipe_localpresetindex),                  //   input,   width = 5,         .i_ch2_txpipe_localpresetindex
		.i_ch2_txpipe_lowpin_nt                         (i_ch2_txpipe_lowpin_nt),                         //   input,   width = 1,         .i_ch2_txpipe_lowpin_nt
		.i_ch2_txpipe_m2p_bus                           (i_ch2_txpipe_m2p_bus),                           //   input,   width = 8,         .i_ch2_txpipe_m2p_bus
		.i_ch2_txpipe_pclk_rate                         (i_ch2_txpipe_pclk_rate),                         //   input,   width = 3,         .i_ch2_txpipe_pclk_rate
		.i_ch2_txpipe_pclkchangeack                     (i_ch2_txpipe_pclkchangeack),                     //   input,   width = 1,         .i_ch2_txpipe_pclkchangeack
		.i_ch2_txpipe_phy_mode_nt                       (i_ch2_txpipe_phy_mode_nt),                       //   input,   width = 4,         .i_ch2_txpipe_phy_mode_nt
		.i_ch2_txpipe_powerdown                         (i_ch2_txpipe_powerdown),                         //   input,   width = 4,         .i_ch2_txpipe_powerdown
		.i_ch2_txpipe_rate                              (i_ch2_txpipe_rate),                              //   input,   width = 3,         .i_ch2_txpipe_rate
		.i_ch2_txpipe_rxelecidle_disable_a              (i_ch2_txpipe_rxelecidle_disable_a),              //   input,   width = 1,         .i_ch2_txpipe_rxelecidle_disable_a
		.i_ch2_txpipe_rxeqclr                           (i_ch2_txpipe_rxeqclr),                           //   input,   width = 1,         .i_ch2_txpipe_rxeqclr
		.i_ch2_txpipe_rxeqeval                          (i_ch2_txpipe_rxeqeval),                          //   input,   width = 1,         .i_ch2_txpipe_rxeqeval
		.i_ch2_txpipe_rxeqinprogress                    (i_ch2_txpipe_rxeqinprogress),                    //   input,   width = 1,         .i_ch2_txpipe_rxeqinprogress
		.i_ch2_txpipe_rxeqtraining                      (i_ch2_txpipe_rxeqtraining),                      //   input,   width = 1,         .i_ch2_txpipe_rxeqtraining
		.i_ch2_txpipe_rxpolarity                        (i_ch2_txpipe_rxpolarity),                        //   input,   width = 1,         .i_ch2_txpipe_rxpolarity
		.i_ch2_txpipe_rxpresethint                      (i_ch2_txpipe_rxpresethint),                      //   input,   width = 3,         .i_ch2_txpipe_rxpresethint
		.i_ch2_txpipe_rxstandby                         (i_ch2_txpipe_rxstandby),                         //   input,   width = 1,         .i_ch2_txpipe_rxstandby
		.i_ch2_txpipe_rxtermination                     (i_ch2_txpipe_rxtermination),                     //   input,   width = 1,         .i_ch2_txpipe_rxtermination
		.i_ch2_txpipe_srisenable                        (i_ch2_txpipe_srisenable),                        //   input,   width = 1,         .i_ch2_txpipe_srisenable
		.i_ch2_txpipe_txcmnmode_disable_a               (i_ch2_txpipe_txcmnmode_disable_a),               //   input,   width = 1,         .i_ch2_txpipe_txcmnmode_disable_a
		.i_ch2_txpipe_txcompliance                      (i_ch2_txpipe_txcompliance),                      //   input,   width = 1,         .i_ch2_txpipe_txcompliance
		.i_ch2_txpipe_txdata                            (i_ch2_txpipe_txdata),                            //   input,  width = 40,         .i_ch2_txpipe_txdata
		.i_ch2_txpipe_txdatak                           (i_ch2_txpipe_txdatak),                           //   input,   width = 4,         .i_ch2_txpipe_txdatak
		.i_ch2_txpipe_txdatavalid                       (i_ch2_txpipe_txdatavalid),                       //   input,   width = 1,         .i_ch2_txpipe_txdatavalid
		.i_ch2_txpipe_txdeemph                          (i_ch2_txpipe_txdeemph),                          //   input,  width = 18,         .i_ch2_txpipe_txdeemph
		.i_ch2_txpipe_txdtctrx_lb                       (i_ch2_txpipe_txdtctrx_lb),                       //   input,   width = 1,         .i_ch2_txpipe_txdtctrx_lb
		.i_ch2_txpipe_txelecidle                        (i_ch2_txpipe_txelecidle),                        //   input,   width = 1,         .i_ch2_txpipe_txelecidle
		.i_ch2_txpipe_txmargin                          (i_ch2_txpipe_txmargin),                          //   input,   width = 3,         .i_ch2_txpipe_txmargin
		.i_ch2_txpipe_txoneszeros                       (i_ch2_txpipe_txoneszeros),                       //   input,   width = 1,         .i_ch2_txpipe_txoneszeros
		.i_ch2_txpipe_txstartblock                      (i_ch2_txpipe_txstartblock),                      //   input,   width = 1,         .i_ch2_txpipe_txstartblock
		.i_ch2_txpipe_txswing                           (i_ch2_txpipe_txswing),                           //   input,   width = 1,         .i_ch2_txpipe_txswing
		.i_ch2_txpipe_txsyncheader                      (i_ch2_txpipe_txsyncheader),                      //   input,   width = 4,         .i_ch2_txpipe_txsyncheader
		.i_ch2_txpipe_width                             (i_ch2_txpipe_width),                             //   input,   width = 3,         .i_ch2_txpipe_width
		.i_ch2_uxq_rxcdrlock2dataa                      (i_ch2_uxq_rxcdrlock2dataa),                      //   input,   width = 1,         .i_ch2_uxq_rxcdrlock2dataa
		.i_ch2_uxq_rxeq_best_eye_vala                   (i_ch2_uxq_rxeq_best_eye_vala),                   //   input,  width = 14,         .i_ch2_uxq_rxeq_best_eye_vala
		.i_ch2_uxq_rxeq_donea                           (i_ch2_uxq_rxeq_donea),                           //   input,   width = 1,         .i_ch2_uxq_rxeq_donea
		.i_ch2_uxq_rxmargin_nacka                       (i_ch2_uxq_rxmargin_nacka),                       //   input,   width = 1,         .i_ch2_uxq_rxmargin_nacka
		.i_ch2_uxq_rxmargin_status_gray_a               (i_ch2_uxq_rxmargin_status_gray_a),               //   input,   width = 2,         .i_ch2_uxq_rxmargin_status_gray_a
		.i_ch2_uxq_rxmargin_statusa                     (i_ch2_uxq_rxmargin_statusa),                     //   input,   width = 1,         .i_ch2_uxq_rxmargin_statusa
		.i_ch2_uxq_rxsignaldetect_lfpsa                 (i_ch2_uxq_rxsignaldetect_lfpsa),                 //   input,   width = 1,         .i_ch2_uxq_rxsignaldetect_lfpsa
		.i_ch2_uxq_rxsignaldetecta                      (i_ch2_uxq_rxsignaldetecta),                      //   input,   width = 1,         .i_ch2_uxq_rxsignaldetecta
		.i_ch2_uxq_rxstatusa                            (i_ch2_uxq_rxstatusa),                            //   input,   width = 1,         .i_ch2_uxq_rxstatusa
		.i_ch2_uxq_rxword                               (i_ch2_uxq_rxword),                               //   input,  width = 40,         .i_ch2_uxq_rxword
		.i_ch2_uxq_synthlcfast_postdiv                  (i_ch2_uxq_synthlcfast_postdiv),                  //   input,   width = 1,         .i_ch2_uxq_synthlcfast_postdiv
		.i_ch2_uxq_synthlcmed_postdiv                   (i_ch2_uxq_synthlcmed_postdiv),                   //   input,   width = 1,         .i_ch2_uxq_synthlcmed_postdiv
		.i_ch2_uxq_synthlcslow_postdiv                  (i_ch2_uxq_synthlcslow_postdiv),                  //   input,   width = 1,         .i_ch2_uxq_synthlcslow_postdiv
		.i_ch2_uxq_txdetectrx_acka                      (i_ch2_uxq_txdetectrx_acka),                      //   input,   width = 1,         .i_ch2_uxq_txdetectrx_acka
		.i_ch2_uxq_txdetectrx_statct                    (i_ch2_uxq_txdetectrx_statct),                    //   input,   width = 1,         .i_ch2_uxq_txdetectrx_statct
		.i_ch2_uxq_txstatusa                            (i_ch2_uxq_txstatusa),                            //   input,   width = 1,         .i_ch2_uxq_txstatusa
		.o_ch2_lavmm_pcie_rdata                         (o_ch2_lavmm_pcie_rdata),                         //  output,  width = 32,         .o_ch2_lavmm_pcie_rdata
		.o_ch2_lavmm_pcie_rdata_valid                   (o_ch2_lavmm_pcie_rdata_valid),                   //  output,   width = 1,         .o_ch2_lavmm_pcie_rdata_valid
		.o_ch2_lavmm_pcie_waitreq                       (o_ch2_lavmm_pcie_waitreq),                       //  output,   width = 1,         .o_ch2_lavmm_pcie_waitreq
		.o_ch2_pcs_pclk                                 (o_ch2_pcs_pclk),                                 //  output,   width = 1,         .o_ch2_pcs_pclk
		.o_ch2_pcs_pipe_rstn                            (o_ch2_pcs_pipe_rstn),                            //  output,   width = 1,         .o_ch2_pcs_pipe_rstn
		.o_ch2_rxpipe_dirfeedback                       (o_ch2_rxpipe_dirfeedback),                       //  output,   width = 6,         .o_ch2_rxpipe_dirfeedback
		.o_ch2_rxpipe_linkevaluationfeedbackfiguremerit (o_ch2_rxpipe_linkevaluationfeedbackfiguremerit), //  output,   width = 8,         .o_ch2_rxpipe_linkevaluationfeedbackfiguremerit
		.o_ch2_rxpipe_localfs                           (o_ch2_rxpipe_localfs),                           //  output,   width = 6,         .o_ch2_rxpipe_localfs
		.o_ch2_rxpipe_locallf                           (o_ch2_rxpipe_locallf),                           //  output,   width = 6,         .o_ch2_rxpipe_locallf
		.o_ch2_rxpipe_localtxcoefficientsvalid          (o_ch2_rxpipe_localtxcoefficientsvalid),          //  output,   width = 1,         .o_ch2_rxpipe_localtxcoefficientsvalid
		.o_ch2_rxpipe_localtxpresetcoefficients         (o_ch2_rxpipe_localtxpresetcoefficients),         //  output,  width = 18,         .o_ch2_rxpipe_localtxpresetcoefficients
		.o_ch2_rxpipe_p2m_bus                           (o_ch2_rxpipe_p2m_bus),                           //  output,   width = 8,         .o_ch2_rxpipe_p2m_bus
		.o_ch2_rxpipe_pclkchangeok                      (o_ch2_rxpipe_pclkchangeok),                      //  output,   width = 1,         .o_ch2_rxpipe_pclkchangeok
		.o_ch2_rxpipe_phystatus                         (o_ch2_rxpipe_phystatus),                         //  output,   width = 1,         .o_ch2_rxpipe_phystatus
		.o_ch2_rxpipe_rxdata                            (o_ch2_rxpipe_rxdata),                            //  output,  width = 40,         .o_ch2_rxpipe_rxdata
		.o_ch2_rxpipe_rxdatak                           (o_ch2_rxpipe_rxdatak),                           //  output,   width = 4,         .o_ch2_rxpipe_rxdatak
		.o_ch2_rxpipe_rxdatavalid                       (o_ch2_rxpipe_rxdatavalid),                       //  output,   width = 1,         .o_ch2_rxpipe_rxdatavalid
		.o_ch2_rxpipe_rxelecidlea                       (o_ch2_rxpipe_rxelecidlea),                       //  output,   width = 1,         .o_ch2_rxpipe_rxelecidlea
		.o_ch2_rxpipe_rxstandbystatus                   (o_ch2_rxpipe_rxstandbystatus),                   //  output,   width = 1,         .o_ch2_rxpipe_rxstandbystatus
		.o_ch2_rxpipe_rxstartblock                      (o_ch2_rxpipe_rxstartblock),                      //  output,   width = 1,         .o_ch2_rxpipe_rxstartblock
		.o_ch2_rxpipe_rxstatus                          (o_ch2_rxpipe_rxstatus),                          //  output,   width = 3,         .o_ch2_rxpipe_rxstatus
		.o_ch2_rxpipe_rxsyncheader                      (o_ch2_rxpipe_rxsyncheader),                      //  output,   width = 4,         .o_ch2_rxpipe_rxsyncheader
		.o_ch2_rxpipe_rxvalid                           (o_ch2_rxpipe_rxvalid),                           //  output,   width = 1,         .o_ch2_rxpipe_rxvalid
		.o_ch2_ux_ock_pma_clk                           (o_ch2_ux_ock_pma_clk),                           //  output,   width = 1,         .o_ch2_ux_ock_pma_clk
		.o_ch2_uxq_lfps_ennt                            (o_ch2_uxq_lfps_ennt),                            //  output,   width = 1,         .o_ch2_uxq_lfps_ennt
		.o_ch2_uxq_pcie_l1ctrla                         (o_ch2_uxq_pcie_l1ctrla),                         //  output,   width = 2,         .o_ch2_uxq_pcie_l1ctrla
		.o_ch2_uxq_pma_cmn_ctrl                         (o_ch2_uxq_pma_cmn_ctrl),                         //  output,   width = 1,         .o_ch2_uxq_pma_cmn_ctrl
		.o_ch2_uxq_pma_ctrl                             (o_ch2_uxq_pma_ctrl),                             //  output,   width = 1,         .o_ch2_uxq_pma_ctrl
		.o_ch2_uxq_rst_pcs_rx_b_a                       (o_ch2_uxq_rst_pcs_rx_b_a),                       //  output,   width = 1,         .o_ch2_uxq_rst_pcs_rx_b_a
		.o_ch2_uxq_rst_pcs_tx_b_a                       (o_ch2_uxq_rst_pcs_tx_b_a),                       //  output,   width = 1,         .o_ch2_uxq_rst_pcs_tx_b_a
		.o_ch2_uxq_rxeiosdetectstata                    (o_ch2_uxq_rxeiosdetectstata),                    //  output,   width = 1,         .o_ch2_uxq_rxeiosdetectstata
		.o_ch2_uxq_rxeq_precal_code_selnt               (o_ch2_uxq_rxeq_precal_code_selnt),               //  output,   width = 3,         .o_ch2_uxq_rxeq_precal_code_selnt
		.o_ch2_uxq_rxeq_starta                          (o_ch2_uxq_rxeq_starta),                          //  output,   width = 1,         .o_ch2_uxq_rxeq_starta
		.o_ch2_uxq_rxeq_static_ena                      (o_ch2_uxq_rxeq_static_ena),                      //  output,   width = 1,         .o_ch2_uxq_rxeq_static_ena
		.o_ch2_uxq_rxmargin_direction_nt                (o_ch2_uxq_rxmargin_direction_nt),                //  output,   width = 1,         .o_ch2_uxq_rxmargin_direction_nt
		.o_ch2_uxq_rxmargin_mode_nt                     (o_ch2_uxq_rxmargin_mode_nt),                     //  output,   width = 1,         .o_ch2_uxq_rxmargin_mode_nt
		.o_ch2_uxq_rxmargin_offset_change_a             (o_ch2_uxq_rxmargin_offset_change_a),             //  output,   width = 1,         .o_ch2_uxq_rxmargin_offset_change_a
		.o_ch2_uxq_rxmargin_offset_nt                   (o_ch2_uxq_rxmargin_offset_nt),                   //  output,   width = 7,         .o_ch2_uxq_rxmargin_offset_nt
		.o_ch2_uxq_rxmargin_start_a                     (o_ch2_uxq_rxmargin_start_a),                     //  output,   width = 1,         .o_ch2_uxq_rxmargin_start_a
		.o_ch2_uxq_rxpstate                             (o_ch2_uxq_rxpstate),                             //  output,   width = 3,         .o_ch2_uxq_rxpstate
		.o_ch2_uxq_rxrate                               (o_ch2_uxq_rxrate),                               //  output,   width = 4,         .o_ch2_uxq_rxrate
		.o_ch2_uxq_rxterm_hiz_ena                       (o_ch2_uxq_rxterm_hiz_ena),                       //  output,   width = 1,         .o_ch2_uxq_rxterm_hiz_ena
		.o_ch2_uxq_rxwidth                              (o_ch2_uxq_rxwidth),                              //  output,   width = 3,         .o_ch2_uxq_rxwidth
		.o_ch2_uxq_tstbus_lane                          (o_ch2_uxq_tstbus_lane),                          //  output,   width = 1,         .o_ch2_uxq_tstbus_lane
		.o_ch2_uxq_txbeacona                            (o_ch2_uxq_txbeacona),                            //  output,   width = 1,         .o_ch2_uxq_txbeacona
		.o_ch2_uxq_txclkdivrate                         (o_ch2_uxq_txclkdivrate),                         //  output,   width = 3,         .o_ch2_uxq_txclkdivrate
		.o_ch2_uxq_txdetectrx_reqa                      (o_ch2_uxq_txdetectrx_reqa),                      //  output,   width = 1,         .o_ch2_uxq_txdetectrx_reqa
		.o_ch2_uxq_txdrv_levn                           (o_ch2_uxq_txdrv_levn),                           //  output,   width = 6,         .o_ch2_uxq_txdrv_levn
		.o_ch2_uxq_txdrv_levnm1                         (o_ch2_uxq_txdrv_levnm1),                         //  output,   width = 5,         .o_ch2_uxq_txdrv_levnm1
		.o_ch2_uxq_txdrv_levnm2                         (o_ch2_uxq_txdrv_levnm2),                         //  output,   width = 3,         .o_ch2_uxq_txdrv_levnm2
		.o_ch2_uxq_txdrv_levnp1                         (o_ch2_uxq_txdrv_levnp1),                         //  output,   width = 5,         .o_ch2_uxq_txdrv_levnp1
		.o_ch2_uxq_txdrv_slew                           (o_ch2_uxq_txdrv_slew),                           //  output,   width = 4,         .o_ch2_uxq_txdrv_slew
		.o_ch2_uxq_txelecidle                           (o_ch2_uxq_txelecidle),                           //  output,   width = 4,         .o_ch2_uxq_txelecidle
		.o_ch2_uxq_txpstate                             (o_ch2_uxq_txpstate),                             //  output,   width = 3,         .o_ch2_uxq_txpstate
		.o_ch2_uxq_txrate                               (o_ch2_uxq_txrate),                               //  output,   width = 4,         .o_ch2_uxq_txrate
		.o_ch2_uxq_txwidth                              (o_ch2_uxq_txwidth),                              //  output,   width = 3,         .o_ch2_uxq_txwidth
		.o_ch2_uxq_txword                               (o_ch2_uxq_txword),                               //  output,  width = 40,         .o_ch2_uxq_txword
		.i_ch3_lavmm_pcie_addr                          (i_ch3_lavmm_pcie_addr),                          //   input,  width = 17,         .i_ch3_lavmm_pcie_addr
		.i_ch3_lavmm_pcie_be                            (i_ch3_lavmm_pcie_be),                            //   input,   width = 4,         .i_ch3_lavmm_pcie_be
		.i_ch3_lavmm_pcie_clk                           (i_ch3_lavmm_pcie_clk),                           //   input,   width = 1,         .i_ch3_lavmm_pcie_clk
		.i_ch3_lavmm_pcie_read                          (i_ch3_lavmm_pcie_read),                          //   input,   width = 1,         .i_ch3_lavmm_pcie_read
		.i_ch3_lavmm_pcie_rstn                          (i_ch3_lavmm_pcie_rstn),                          //   input,   width = 1,         .i_ch3_lavmm_pcie_rstn
		.i_ch3_lavmm_pcie_wdata                         (i_ch3_lavmm_pcie_wdata),                         //   input,  width = 32,         .i_ch3_lavmm_pcie_wdata
		.i_ch3_lavmm_pcie_write                         (i_ch3_lavmm_pcie_write),                         //   input,   width = 1,         .i_ch3_lavmm_pcie_write
		.i_ch3_pcie_rxword_clk                          (i_ch3_pcie_rxword_clk),                          //   input,   width = 1,         .i_ch3_pcie_rxword_clk
		.i_ch3_pcie_txword_clk                          (i_ch3_pcie_txword_clk),                          //   input,   width = 1,         .i_ch3_pcie_txword_clk
		.i_ch3_pcs_pclk                                 (i_ch3_pcs_pclk),                                 //   input,   width = 1,         .i_ch3_pcs_pclk
		.i_ch3_pcs_pipe_rstn                            (i_ch3_pcs_pipe_rstn),                            //   input,   width = 1,         .i_ch3_pcs_pipe_rstn
		.i_ch3_txpipe_asyncpowerchangeack               (i_ch3_txpipe_asyncpowerchangeack),               //   input,   width = 1,         .i_ch3_txpipe_asyncpowerchangeack
		.i_ch3_txpipe_blockaligncontrol                 (i_ch3_txpipe_blockaligncontrol),                 //   input,   width = 1,         .i_ch3_txpipe_blockaligncontrol
		.i_ch3_txpipe_cfg_hw_auto_sp_dis                (i_ch3_txpipe_cfg_hw_auto_sp_dis),                //   input,   width = 1,         .i_ch3_txpipe_cfg_hw_auto_sp_dis
		.i_ch3_txpipe_dirchange                         (i_ch3_txpipe_dirchange),                         //   input,   width = 1,         .i_ch3_txpipe_dirchange
		.i_ch3_txpipe_ebuf_mode                         (i_ch3_txpipe_ebuf_mode),                         //   input,   width = 1,         .i_ch3_txpipe_ebuf_mode
		.i_ch3_txpipe_encodedecodebypass                (i_ch3_txpipe_encodedecodebypass),                //   input,   width = 1,         .i_ch3_txpipe_encodedecodebypass
		.i_ch3_txpipe_fs                                (i_ch3_txpipe_fs),                                //   input,   width = 6,         .i_ch3_txpipe_fs
		.i_ch3_txpipe_getlocalpresetcoefficients        (i_ch3_txpipe_getlocalpresetcoefficients),        //   input,   width = 1,         .i_ch3_txpipe_getlocalpresetcoefficients
		.i_ch3_txpipe_invalidrequest                    (i_ch3_txpipe_invalidrequest),                    //   input,   width = 1,         .i_ch3_txpipe_invalidrequest
		.i_ch3_txpipe_lf                                (i_ch3_txpipe_lf),                                //   input,   width = 6,         .i_ch3_txpipe_lf
		.i_ch3_txpipe_localpresetindex                  (i_ch3_txpipe_localpresetindex),                  //   input,   width = 5,         .i_ch3_txpipe_localpresetindex
		.i_ch3_txpipe_lowpin_nt                         (i_ch3_txpipe_lowpin_nt),                         //   input,   width = 1,         .i_ch3_txpipe_lowpin_nt
		.i_ch3_txpipe_m2p_bus                           (i_ch3_txpipe_m2p_bus),                           //   input,   width = 8,         .i_ch3_txpipe_m2p_bus
		.i_ch3_txpipe_pclk_rate                         (i_ch3_txpipe_pclk_rate),                         //   input,   width = 3,         .i_ch3_txpipe_pclk_rate
		.i_ch3_txpipe_pclkchangeack                     (i_ch3_txpipe_pclkchangeack),                     //   input,   width = 1,         .i_ch3_txpipe_pclkchangeack
		.i_ch3_txpipe_phy_mode_nt                       (i_ch3_txpipe_phy_mode_nt),                       //   input,   width = 4,         .i_ch3_txpipe_phy_mode_nt
		.i_ch3_txpipe_powerdown                         (i_ch3_txpipe_powerdown),                         //   input,   width = 4,         .i_ch3_txpipe_powerdown
		.i_ch3_txpipe_rate                              (i_ch3_txpipe_rate),                              //   input,   width = 3,         .i_ch3_txpipe_rate
		.i_ch3_txpipe_rxelecidle_disable_a              (i_ch3_txpipe_rxelecidle_disable_a),              //   input,   width = 1,         .i_ch3_txpipe_rxelecidle_disable_a
		.i_ch3_txpipe_rxeqclr                           (i_ch3_txpipe_rxeqclr),                           //   input,   width = 1,         .i_ch3_txpipe_rxeqclr
		.i_ch3_txpipe_rxeqeval                          (i_ch3_txpipe_rxeqeval),                          //   input,   width = 1,         .i_ch3_txpipe_rxeqeval
		.i_ch3_txpipe_rxeqinprogress                    (i_ch3_txpipe_rxeqinprogress),                    //   input,   width = 1,         .i_ch3_txpipe_rxeqinprogress
		.i_ch3_txpipe_rxeqtraining                      (i_ch3_txpipe_rxeqtraining),                      //   input,   width = 1,         .i_ch3_txpipe_rxeqtraining
		.i_ch3_txpipe_rxpolarity                        (i_ch3_txpipe_rxpolarity),                        //   input,   width = 1,         .i_ch3_txpipe_rxpolarity
		.i_ch3_txpipe_rxpresethint                      (i_ch3_txpipe_rxpresethint),                      //   input,   width = 3,         .i_ch3_txpipe_rxpresethint
		.i_ch3_txpipe_rxstandby                         (i_ch3_txpipe_rxstandby),                         //   input,   width = 1,         .i_ch3_txpipe_rxstandby
		.i_ch3_txpipe_rxtermination                     (i_ch3_txpipe_rxtermination),                     //   input,   width = 1,         .i_ch3_txpipe_rxtermination
		.i_ch3_txpipe_srisenable                        (i_ch3_txpipe_srisenable),                        //   input,   width = 1,         .i_ch3_txpipe_srisenable
		.i_ch3_txpipe_txcmnmode_disable_a               (i_ch3_txpipe_txcmnmode_disable_a),               //   input,   width = 1,         .i_ch3_txpipe_txcmnmode_disable_a
		.i_ch3_txpipe_txcompliance                      (i_ch3_txpipe_txcompliance),                      //   input,   width = 1,         .i_ch3_txpipe_txcompliance
		.i_ch3_txpipe_txdata                            (i_ch3_txpipe_txdata),                            //   input,  width = 40,         .i_ch3_txpipe_txdata
		.i_ch3_txpipe_txdatak                           (i_ch3_txpipe_txdatak),                           //   input,   width = 4,         .i_ch3_txpipe_txdatak
		.i_ch3_txpipe_txdatavalid                       (i_ch3_txpipe_txdatavalid),                       //   input,   width = 1,         .i_ch3_txpipe_txdatavalid
		.i_ch3_txpipe_txdeemph                          (i_ch3_txpipe_txdeemph),                          //   input,  width = 18,         .i_ch3_txpipe_txdeemph
		.i_ch3_txpipe_txdtctrx_lb                       (i_ch3_txpipe_txdtctrx_lb),                       //   input,   width = 1,         .i_ch3_txpipe_txdtctrx_lb
		.i_ch3_txpipe_txelecidle                        (i_ch3_txpipe_txelecidle),                        //   input,   width = 1,         .i_ch3_txpipe_txelecidle
		.i_ch3_txpipe_txmargin                          (i_ch3_txpipe_txmargin),                          //   input,   width = 3,         .i_ch3_txpipe_txmargin
		.i_ch3_txpipe_txoneszeros                       (i_ch3_txpipe_txoneszeros),                       //   input,   width = 1,         .i_ch3_txpipe_txoneszeros
		.i_ch3_txpipe_txstartblock                      (i_ch3_txpipe_txstartblock),                      //   input,   width = 1,         .i_ch3_txpipe_txstartblock
		.i_ch3_txpipe_txswing                           (i_ch3_txpipe_txswing),                           //   input,   width = 1,         .i_ch3_txpipe_txswing
		.i_ch3_txpipe_txsyncheader                      (i_ch3_txpipe_txsyncheader),                      //   input,   width = 4,         .i_ch3_txpipe_txsyncheader
		.i_ch3_txpipe_width                             (i_ch3_txpipe_width),                             //   input,   width = 3,         .i_ch3_txpipe_width
		.i_ch3_uxq_rxcdrlock2dataa                      (i_ch3_uxq_rxcdrlock2dataa),                      //   input,   width = 1,         .i_ch3_uxq_rxcdrlock2dataa
		.i_ch3_uxq_rxeq_best_eye_vala                   (i_ch3_uxq_rxeq_best_eye_vala),                   //   input,  width = 14,         .i_ch3_uxq_rxeq_best_eye_vala
		.i_ch3_uxq_rxeq_donea                           (i_ch3_uxq_rxeq_donea),                           //   input,   width = 1,         .i_ch3_uxq_rxeq_donea
		.i_ch3_uxq_rxmargin_nacka                       (i_ch3_uxq_rxmargin_nacka),                       //   input,   width = 1,         .i_ch3_uxq_rxmargin_nacka
		.i_ch3_uxq_rxmargin_status_gray_a               (i_ch3_uxq_rxmargin_status_gray_a),               //   input,   width = 2,         .i_ch3_uxq_rxmargin_status_gray_a
		.i_ch3_uxq_rxmargin_statusa                     (i_ch3_uxq_rxmargin_statusa),                     //   input,   width = 1,         .i_ch3_uxq_rxmargin_statusa
		.i_ch3_uxq_rxsignaldetect_lfpsa                 (i_ch3_uxq_rxsignaldetect_lfpsa),                 //   input,   width = 1,         .i_ch3_uxq_rxsignaldetect_lfpsa
		.i_ch3_uxq_rxsignaldetecta                      (i_ch3_uxq_rxsignaldetecta),                      //   input,   width = 1,         .i_ch3_uxq_rxsignaldetecta
		.i_ch3_uxq_rxstatusa                            (i_ch3_uxq_rxstatusa),                            //   input,   width = 1,         .i_ch3_uxq_rxstatusa
		.i_ch3_uxq_rxword                               (i_ch3_uxq_rxword),                               //   input,  width = 40,         .i_ch3_uxq_rxword
		.i_ch3_uxq_synthlcfast_postdiv                  (i_ch3_uxq_synthlcfast_postdiv),                  //   input,   width = 1,         .i_ch3_uxq_synthlcfast_postdiv
		.i_ch3_uxq_synthlcmed_postdiv                   (i_ch3_uxq_synthlcmed_postdiv),                   //   input,   width = 1,         .i_ch3_uxq_synthlcmed_postdiv
		.i_ch3_uxq_synthlcslow_postdiv                  (i_ch3_uxq_synthlcslow_postdiv),                  //   input,   width = 1,         .i_ch3_uxq_synthlcslow_postdiv
		.i_ch3_uxq_txdetectrx_acka                      (i_ch3_uxq_txdetectrx_acka),                      //   input,   width = 1,         .i_ch3_uxq_txdetectrx_acka
		.i_ch3_uxq_txdetectrx_statct                    (i_ch3_uxq_txdetectrx_statct),                    //   input,   width = 1,         .i_ch3_uxq_txdetectrx_statct
		.i_ch3_uxq_txstatusa                            (i_ch3_uxq_txstatusa),                            //   input,   width = 1,         .i_ch3_uxq_txstatusa
		.o_ch3_lavmm_pcie_rdata                         (o_ch3_lavmm_pcie_rdata),                         //  output,  width = 32,         .o_ch3_lavmm_pcie_rdata
		.o_ch3_lavmm_pcie_rdata_valid                   (o_ch3_lavmm_pcie_rdata_valid),                   //  output,   width = 1,         .o_ch3_lavmm_pcie_rdata_valid
		.o_ch3_lavmm_pcie_waitreq                       (o_ch3_lavmm_pcie_waitreq),                       //  output,   width = 1,         .o_ch3_lavmm_pcie_waitreq
		.o_ch3_pcs_pclk                                 (o_ch3_pcs_pclk),                                 //  output,   width = 1,         .o_ch3_pcs_pclk
		.o_ch3_pcs_pipe_rstn                            (o_ch3_pcs_pipe_rstn),                            //  output,   width = 1,         .o_ch3_pcs_pipe_rstn
		.o_ch3_rxpipe_dirfeedback                       (o_ch3_rxpipe_dirfeedback),                       //  output,   width = 6,         .o_ch3_rxpipe_dirfeedback
		.o_ch3_rxpipe_linkevaluationfeedbackfiguremerit (o_ch3_rxpipe_linkevaluationfeedbackfiguremerit), //  output,   width = 8,         .o_ch3_rxpipe_linkevaluationfeedbackfiguremerit
		.o_ch3_rxpipe_localfs                           (o_ch3_rxpipe_localfs),                           //  output,   width = 6,         .o_ch3_rxpipe_localfs
		.o_ch3_rxpipe_locallf                           (o_ch3_rxpipe_locallf),                           //  output,   width = 6,         .o_ch3_rxpipe_locallf
		.o_ch3_rxpipe_localtxcoefficientsvalid          (o_ch3_rxpipe_localtxcoefficientsvalid),          //  output,   width = 1,         .o_ch3_rxpipe_localtxcoefficientsvalid
		.o_ch3_rxpipe_localtxpresetcoefficients         (o_ch3_rxpipe_localtxpresetcoefficients),         //  output,  width = 18,         .o_ch3_rxpipe_localtxpresetcoefficients
		.o_ch3_rxpipe_p2m_bus                           (o_ch3_rxpipe_p2m_bus),                           //  output,   width = 8,         .o_ch3_rxpipe_p2m_bus
		.o_ch3_rxpipe_pclkchangeok                      (o_ch3_rxpipe_pclkchangeok),                      //  output,   width = 1,         .o_ch3_rxpipe_pclkchangeok
		.o_ch3_rxpipe_phystatus                         (o_ch3_rxpipe_phystatus),                         //  output,   width = 1,         .o_ch3_rxpipe_phystatus
		.o_ch3_rxpipe_rxdata                            (o_ch3_rxpipe_rxdata),                            //  output,  width = 40,         .o_ch3_rxpipe_rxdata
		.o_ch3_rxpipe_rxdatak                           (o_ch3_rxpipe_rxdatak),                           //  output,   width = 4,         .o_ch3_rxpipe_rxdatak
		.o_ch3_rxpipe_rxdatavalid                       (o_ch3_rxpipe_rxdatavalid),                       //  output,   width = 1,         .o_ch3_rxpipe_rxdatavalid
		.o_ch3_rxpipe_rxelecidlea                       (o_ch3_rxpipe_rxelecidlea),                       //  output,   width = 1,         .o_ch3_rxpipe_rxelecidlea
		.o_ch3_rxpipe_rxstandbystatus                   (o_ch3_rxpipe_rxstandbystatus),                   //  output,   width = 1,         .o_ch3_rxpipe_rxstandbystatus
		.o_ch3_rxpipe_rxstartblock                      (o_ch3_rxpipe_rxstartblock),                      //  output,   width = 1,         .o_ch3_rxpipe_rxstartblock
		.o_ch3_rxpipe_rxstatus                          (o_ch3_rxpipe_rxstatus),                          //  output,   width = 3,         .o_ch3_rxpipe_rxstatus
		.o_ch3_rxpipe_rxsyncheader                      (o_ch3_rxpipe_rxsyncheader),                      //  output,   width = 4,         .o_ch3_rxpipe_rxsyncheader
		.o_ch3_rxpipe_rxvalid                           (o_ch3_rxpipe_rxvalid),                           //  output,   width = 1,         .o_ch3_rxpipe_rxvalid
		.o_ch3_ux_ock_pma_clk                           (o_ch3_ux_ock_pma_clk),                           //  output,   width = 1,         .o_ch3_ux_ock_pma_clk
		.o_ch3_uxq_lfps_ennt                            (o_ch3_uxq_lfps_ennt),                            //  output,   width = 1,         .o_ch3_uxq_lfps_ennt
		.o_ch3_uxq_pcie_l1ctrla                         (o_ch3_uxq_pcie_l1ctrla),                         //  output,   width = 2,         .o_ch3_uxq_pcie_l1ctrla
		.o_ch3_uxq_pma_cmn_ctrl                         (o_ch3_uxq_pma_cmn_ctrl),                         //  output,   width = 1,         .o_ch3_uxq_pma_cmn_ctrl
		.o_ch3_uxq_pma_ctrl                             (o_ch3_uxq_pma_ctrl),                             //  output,   width = 1,         .o_ch3_uxq_pma_ctrl
		.o_ch3_uxq_rst_pcs_rx_b_a                       (o_ch3_uxq_rst_pcs_rx_b_a),                       //  output,   width = 1,         .o_ch3_uxq_rst_pcs_rx_b_a
		.o_ch3_uxq_rst_pcs_tx_b_a                       (o_ch3_uxq_rst_pcs_tx_b_a),                       //  output,   width = 1,         .o_ch3_uxq_rst_pcs_tx_b_a
		.o_ch3_uxq_rxeiosdetectstata                    (o_ch3_uxq_rxeiosdetectstata),                    //  output,   width = 1,         .o_ch3_uxq_rxeiosdetectstata
		.o_ch3_uxq_rxeq_precal_code_selnt               (o_ch3_uxq_rxeq_precal_code_selnt),               //  output,   width = 3,         .o_ch3_uxq_rxeq_precal_code_selnt
		.o_ch3_uxq_rxeq_starta                          (o_ch3_uxq_rxeq_starta),                          //  output,   width = 1,         .o_ch3_uxq_rxeq_starta
		.o_ch3_uxq_rxeq_static_ena                      (o_ch3_uxq_rxeq_static_ena),                      //  output,   width = 1,         .o_ch3_uxq_rxeq_static_ena
		.o_ch3_uxq_rxmargin_direction_nt                (o_ch3_uxq_rxmargin_direction_nt),                //  output,   width = 1,         .o_ch3_uxq_rxmargin_direction_nt
		.o_ch3_uxq_rxmargin_mode_nt                     (o_ch3_uxq_rxmargin_mode_nt),                     //  output,   width = 1,         .o_ch3_uxq_rxmargin_mode_nt
		.o_ch3_uxq_rxmargin_offset_change_a             (o_ch3_uxq_rxmargin_offset_change_a),             //  output,   width = 1,         .o_ch3_uxq_rxmargin_offset_change_a
		.o_ch3_uxq_rxmargin_offset_nt                   (o_ch3_uxq_rxmargin_offset_nt),                   //  output,   width = 7,         .o_ch3_uxq_rxmargin_offset_nt
		.o_ch3_uxq_rxmargin_start_a                     (o_ch3_uxq_rxmargin_start_a),                     //  output,   width = 1,         .o_ch3_uxq_rxmargin_start_a
		.o_ch3_uxq_rxpstate                             (o_ch3_uxq_rxpstate),                             //  output,   width = 3,         .o_ch3_uxq_rxpstate
		.o_ch3_uxq_rxrate                               (o_ch3_uxq_rxrate),                               //  output,   width = 4,         .o_ch3_uxq_rxrate
		.o_ch3_uxq_rxterm_hiz_ena                       (o_ch3_uxq_rxterm_hiz_ena),                       //  output,   width = 1,         .o_ch3_uxq_rxterm_hiz_ena
		.o_ch3_uxq_rxwidth                              (o_ch3_uxq_rxwidth),                              //  output,   width = 3,         .o_ch3_uxq_rxwidth
		.o_ch3_uxq_tstbus_lane                          (o_ch3_uxq_tstbus_lane),                          //  output,   width = 1,         .o_ch3_uxq_tstbus_lane
		.o_ch3_uxq_txbeacona                            (o_ch3_uxq_txbeacona),                            //  output,   width = 1,         .o_ch3_uxq_txbeacona
		.o_ch3_uxq_txclkdivrate                         (o_ch3_uxq_txclkdivrate),                         //  output,   width = 3,         .o_ch3_uxq_txclkdivrate
		.o_ch3_uxq_txdetectrx_reqa                      (o_ch3_uxq_txdetectrx_reqa),                      //  output,   width = 1,         .o_ch3_uxq_txdetectrx_reqa
		.o_ch3_uxq_txdrv_levn                           (o_ch3_uxq_txdrv_levn),                           //  output,   width = 6,         .o_ch3_uxq_txdrv_levn
		.o_ch3_uxq_txdrv_levnm1                         (o_ch3_uxq_txdrv_levnm1),                         //  output,   width = 5,         .o_ch3_uxq_txdrv_levnm1
		.o_ch3_uxq_txdrv_levnm2                         (o_ch3_uxq_txdrv_levnm2),                         //  output,   width = 3,         .o_ch3_uxq_txdrv_levnm2
		.o_ch3_uxq_txdrv_levnp1                         (o_ch3_uxq_txdrv_levnp1),                         //  output,   width = 5,         .o_ch3_uxq_txdrv_levnp1
		.o_ch3_uxq_txdrv_slew                           (o_ch3_uxq_txdrv_slew),                           //  output,   width = 4,         .o_ch3_uxq_txdrv_slew
		.o_ch3_uxq_txelecidle                           (o_ch3_uxq_txelecidle),                           //  output,   width = 4,         .o_ch3_uxq_txelecidle
		.o_ch3_uxq_txpstate                             (o_ch3_uxq_txpstate),                             //  output,   width = 3,         .o_ch3_uxq_txpstate
		.o_ch3_uxq_txrate                               (o_ch3_uxq_txrate),                               //  output,   width = 4,         .o_ch3_uxq_txrate
		.o_ch3_uxq_txwidth                              (o_ch3_uxq_txwidth),                              //  output,   width = 3,         .o_ch3_uxq_txwidth
		.o_ch3_uxq_txword                               (o_ch3_uxq_txword)                                //  output,  width = 40,         .o_ch3_uxq_txword
	);

endmodule
