// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oL5o3zdpsF8kSnwevvpcVj/H1FZmzc1oRwNmgViSjWZH8LNj7/Wzob0/XK8B
L64ugFI1s2mdbMq5wp0+k4PAC7d+FUca+MKQwDe5+YZ1dt+yYXC6rkHVCWcn
QekcmF7ylGNHDqpfgMLCi7F4xoRylc+Oel++Xf5B6b2VTBeCSjL+Ub091ck0
zAVfD5LGl8V17lpyOAEkuYPmFGtiDDmmRFhWDnHud5m9ZO7BMDb3EFAdsvF5
eESm2iReB3QFf7DXOOBua12kEY+pygUzCRbnYJxZj0VNw+3pfK8z+G0cKUgf
0HjcVpqdkBA/3Ixp8ZtCjSfk/ROyb1BySAMSbNlJYg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VJRu8zt7e0hV0rlaI9m9ly6xMfbPdO/uR9MRAvltmXOwdB5Qk6vp/58HMhKJ
YYbmpSlIsKPxDXfHyPbaku2BKdUn4TLMciNM/iujtrLCUlq9ZziKAAIrmRI5
UM2ei6ibC6XQyZhc+jpDKvxiVhoGMl6mMdBWFoUFxyG7pipVokDKtrY0PmMG
tlTkWpnt6t2AP3OUkl8du32guc66IID9G8jugt0hmmt3WyTSNimVSjgSGEmC
SwPenAiTsdeE5VmjLUcfbvLBbiuHmW5ZybhcVZ8IC3P1oVrOCdiAY2SSIlau
H6a6l6UetXERk2BpEkO5P7QYMu2S52GUN8iG1n5SJg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
En/eOUxlurWQejNIKB/YTfO6GzAHbpc1U7onv38bqDrJuBocdO7bPlE0A3Vb
IfIiwt/8NUAH98WLsDRY+Bw7heG3RkipbBfjsnm3CGB8cyafl8shDn/PcfSI
EPKlpIEHTWQEKCYA2wc4pl1NrNJnqRXDKNUum9B5v/B7xgIr7Yx5zF6Vw1sg
q805A3pT1u/Zg9tP7NNDvFoEUjNvTDgERPi8aV/YMscr7W6YVJjWW7dZetcY
nMVtyZ0mqpt/g12tj88stdpz9hIhO6LrDUEjkj8yrxkrQYzjZZwTl1volsgN
+pardji5UrE8nZuKDPsGJZx3OS13OUmFVGygQDoQeg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
V9CQVF07Jcx9vtZihY4OUKR3u7Hz1ni3GllfVlHqx25GPa2HIp4MtI1P3FGt
ZkwnUlfMf+ltIXX/r+GZe+l0pUdcgkjjz9YVzcurfQIqvqV09kGRaY4ROIrp
e1DFpX/sIn/y2/nCNy8Qownf4l9Nmwa6PIZo8RqQm/uGG9xCcJA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HqJPsDQENhG9tQT5pIddnUJPcdNZ1toLjQUUwh9ktXEf3snYlpEUHGs0Gu+A
BpkcTA08kTw1k3NlaxL5AABhFnAAfbYsTK7BJJCjWTgSs13huHq94SoLHqH+
UKLrWFjAP5ZjuNXihTdgzJHGoBwvfySszCilnAp0LQ9c5TF5Ox2GSHvmeBqQ
BQz20Z6BiIqi9TCMxsf+M1Q1otZdBUYoJJpRtdFg+cOHz5vOoBs7bq3bsty4
P1XBDqxb2xwy187WrZRN9sMSfz8E+8MoTZzF8+5ruN9GfWFCmN3X5x+qKgly
AdV9XYeviPS6ejhBR6OGGFURxTL9Hwnax0q2mIb3Nqb2lEeMM2zv9CwNu2h+
jLJiVWo6DRb5rPPcNleFChNbmfibaZgdsXye4x3w0rRGxb0WTY3PXapagP4r
opkMrRtDVYWrguc64wmpoCmnAWdruAQna6TesiK7zRUm00Hkwbu6kVcL3POI
3FoLWx1J3PfzaNfTD5c/Hye45ZXQx0v8


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YWWRjLU/13ReEB19mYOzNXJanzzPg3zb9RamBUW2EH08BKBB0zwiT4DkS8dV
kkmy12TQnmp0SCYjcXVgrtG7g16wCPTTLHoKcwvAi++8Xe2Wei9CLNXjWoLs
No4FjSAnMQ+N5rl+oej+Oz6wL750GMg7d9/92/VYf4lc843IR6Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bWMVuQERxGPJhNz9ji3uMyThxZFRg3W091QRVX+vV8xuXgZZ1zp7MAt7qmG6
ROcGr/mjrm/GAtx9LY5CMYC62izxymAeqQHpZGhTvzEKFz0AXsLcZe50wvVl
CkmZMvScEmySVvrsaFR/kmnS+bhkKcPhuhK1TAcOq8lWEURa+Vk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4512)
`pragma protect data_block
uhMKtLXnAr5/pGOqVTBShygjt1akhS42oaPxXen419X6MzS2C2Bd0Q9ZTQX1
6lzfBrap/H/oM2+GsWHIfwT856ONaNxe5MlIRCjS8MrZJOMQL6zBRkb47zk+
nk/Jn2BL6AMgLNUeZlVkh/uE4vf0WKGgTfPdlB/ObLDXLuIPOBvdtlqbBCjq
xavMXqJarwU8bf5yHY0xMRtJ94HEPAx+6Lt9OGp/RsmgcvX2zOZt1PMLZX6D
PoOlq3+37N9y5uZoB+dHceO9dM5NCbWTzh2YOWSlolc1KpCIU/XCUgoqUP6+
JTP9ehfZc7ILc5c/PT4RhPXK04QRmjheA3to5joIiaOkuSwPGPtAQdtZS0Jv
QOxtdgEmAtiVsznIzVwYg4f0tBcjcouBzA53Yg47eBvN/W3pr0Q0D6FHd/Gv
rk8cj0NSI/KqWdprErLxKPWFiLFOOwIZHWGDcocT8K/cgF5Bp3F22pZw5/iu
24nG6h18o9fN2410abOQC9XMs98I/Xi2VG+qjPobEu/0hZBMMGqIiIzyjS9P
c7Ia4L2TSpXcur/jw5j47WHthdPFeQbB5BnIY59/4xhjMMp/7CqqtB/kfz6p
zDkF9zSq++pw7lcYLEkhYiHLAqO7AJIaE1o9k/KFS0yBysUuUknXbM5HeoQE
0IbEDb4G/hRL58ZS0Bq74HGmJwoX2Cg/4trK4X1LwGEgKX5A7HMshz0UymOd
z4bSVpx4zRrORvR5t5Ydmag91Jk77vbDHAojXvl+xgMs9WSuwFtzbM8QCmrD
pLqYR6HIhn6j8VrBNrcItgIJhM5g44ImFusOq4GjJ8vM3YU0AXHbgTGDWn3X
Ys6THXpmT9/dRCGr1EDAj7z8QIvaQ0jTc+rPcWAwhqQ/si2CloCxI2l6zVj8
UlLL4A8zbQbMeTXlCz0uRvawXo8aI72LqFSfR5ctXngUMq1PwiRPl9ZJps/u
gDX2AD9rHxHpEpNUbCRTotO3oCyjQbB1FtCEbfnjRUvxIn9E4BdHO7NcebRi
TocS7gtKgEuNwdlDMDSdlil6y12csAHSM6erPMKXCWBjJcKqYVOHxVbYeB/T
50L0QZPqpmlTUsJe0hNAFk3fmRaIl2NV0O9aZ6STyfoDmc0wp7sSF2z50Un9
eBToPj9zp44oAykZKjmMXGQbP7fQxN4DFq/rW9lqGN0s3y8G5BliL7cpOJ+/
Xmmj8iDkkWY2VG3S0fFsk0fbGQ8jAkD1FuGoA/QvGYSiZArCXgKapj19iABf
xDp57rsYqp14GOfHpXERpat+Umu3hmKP+XoUiadM/39XiE/33R25+nPKqWjJ
gog6+AXpQL2iuh0xLk0kC1FsXvl09ZuIEWnSRG4wH2w2QthbvaS/tStl/42D
cM42WpIQE/uZO9oD0dtN6cmRj6c/gvvAevcPmxK0qIFYWZ5PEAs2WWQeZ7tK
/dZ0uZNMONaZOEmx3B9/CZ6arP5xlMpQssYoSJOjJNA8//A0OseVFu1mKs9M
K+oejcnee2IhFrX2wN05o9vcfWKap9iNKbJar7rrgKh9sXnROcPo3giOkVKt
pbhlCD2t565akFJphl+FD9HMqF0y9vtRFmQQRyjh0qwEcpGqQiKE1+V++OpL
Wp82CzYkus1aQ1jcI12Wkj+1eUwUUxlWXWnr7aNZgTz1HFQ0nxd+28dK0I3j
nES12aiyUHi+skIhjCvoZKVkbs7TBv/FSlJTuVd/J2ZXts1U7thsC6b9MLds
gvjShH3nRxEh8ghsnx1T6LwhayKCDeqBloNw8gQf9mJgid82mO7fxBCRtmMl
bDd8NRuoSc04pinKDbW8fH0Atcr8gHUXlLvp25QjrCqEGYj7oGG7viD7cLHO
1O+oPLcnd7ztPVH6eHDGqJ7oADdpLm+FhELtely7/AoWoZS01y0+Yl3E1GIp
ODu91VBvo3gYexqzSXlp7F5jDUbLtL7kv9JA8LQTAmJ9u9T+wwKo51aHdPay
giVrHqqyDhltssLV8pVW8URip6zzxDYq/H6+5KRRaFW5B/51re0WsLUaJmKi
B85gwBL/VV3HoYo7GZA5Bsx4qxJRNi0ijoTyX8J4iK1q0v9vvwdb/SejN1kp
yWxMXtkgmfdYALB+IsVfMazElu6frjy+MqHuaTNI4+dIxDqDVo4iPzcFfepg
MCorChlU4/KWn/WlZC/L6Fl7Fa/cKj5DeGgsafm5U7w1rO4Xw8dkkJw1pvXi
D5JjFrDbAzJ56zEAe9f5rcdsLT8NoM0Av6KNzXfJGqy44mA3nLt+A3kfK0/p
HLCuCJCep8zM97TiQpahq22bfvuxG2pe236ug0Y95q9cFlkwDh6Adjynrxx/
KtKfhGbT29ViljZHNNvLbTVwQNUW6cOtCWl3ehGelw/TO3kmTQsOp9rQn0Q7
scd8a4/Vrelq+ixb75Gkz0gTNmTAiFMtwCYWv0g5RM6Csssl5gqs/7IguBLR
PnypLyz6u+HE2upDmcy2VHcB5g5NEdrmKKwUNJDIhoCScp6Whmv8AUzfky8S
Br97gATWCEZNIaSgH3YEhWKNnarM7nL3FQed/3ZmALkzsoP6MtMfMnxG115E
rOm++Cso3RsIPH2CXEwFLw/z2AJJ7rkwLVtFewydlzGlTbK8IX9fTsNtkw0V
s0n7P3HnD4nHlW6jzr7F/INSUIavWSjmZJOOBzZW1E8zpVjYeOCQOugW7lyb
Gx2w29Pn1Q4Cw/gqzZp1kvO2Vf3rq+NUscUu9EOk0k1hiEmyl6OCPo7OW1Kl
6ChH/VGofmBuk4UoYKcQhhvphC4bnbBm6PjHzVs52blOQrBgWqysh1mKavOR
SXDsyc+WHwilgrWYRRL0Ut4td2mISjLOqcJqPPqm+ilitGiDXhi1G6ZEjhFE
fPELwqRsMkUHeBCB6DWleQHod4zk0JV4sKZEbpUyaB+cu1i6XwVALczIZ7LY
QEjhRBSR4S5XnopkcKuOpSHzcKiGgR8SawIeXob0HO/vReBUXF5qLGGJTgVl
DTEiX2LpoE4hSF1bQMdu9DF5NaQ/Ly3TelekKoBHPORuIaQRBbAs2okwupdU
EInN1MdF2kBde4fhiK+8XOX5mO7+TVFS4EbOCHiszCZNdqQQdhKREvJnAqD5
qvVuPDCYIFn/Aar/Zmdd/yA8+1Wztsr4AS5HRJuYZgbWRvDLs0ZgvruQD53i
Pj7MDOLEZp2lElLd8GI5Emv0fv/bMh/LkAJUIrLtkpyAcNFj4naWypRfCWR1
a4wQN4JB89PMN2jWlMgQSurAkb1FHUlKMtBfZzUXr6j8h1pm3Q0HS4tFGhQN
iEi85Ex4AGnS3Ij39GwVmrmvgHXc7sOIPE//xJXblmDTIhzqYtcckYb4T17L
iqRxVvH3Q8mwk0FZ7bhnjnOXNKzO0342XL2oVMArahzPZJ6YhmlFyzAqK78U
pU5+WUa3yQgCmckQpi8J+QHKGfJdiMNx7Os0ps94KbBHaZwviM9V+QaTtRAN
gTmyVX6wQsl8KLsPR2432hYi4JXKx2O6HdnnMbLaK8bc8xYmyGlzGmCC7jL0
kPQkMY3LnNme9Wk8RpyYKvW3H8o3EGlcMHWvCJIprnnt66VtC+LLpIGVPeJ7
l+SkrENFBKVUD49ax4Y9oNP1j9+NOrZ10FcYlZoNkk9xL0mRijTHpRFvtnUm
PyzSgkq4M05VxJjRX/CqXiXcUD+fZJaPN0mtI/qHMFNPGj5Ey8IrLWftB9n0
u7GO1z8phft3/Nlghx/2ybwB49lyi7gu4/oeemJi3bxSXZzz0nClv3feqspz
5GKdPC1iVVJuLNrczYDnzu74cafdC9Avi6ehGUENvNB32OTLmVmV0H6AJuIq
g0XDYDem74+9g50W+JEB74P8GAAn/8LrvMIqFtmTIfvfHJGb/A30d86vfIcD
lYx/DM2FfA1g1fG+Ya6jjGfU3wLe2JFtruV3/I0cq8BW5dSNL7R5gZNl2wRs
S5cgjI1kZ7EUakPgMHNQTfb1RSvbJUZew96Mg0Ai4vC1cYwqwZFuWWqpCDWl
OPF1JVvqdctfyeoXOq/lTk8SXVKSwPBRXJvMIRXLrYB42OiMjNT8CYeExkH3
CwuxERQ7aosAZu12kGWiU3x4RoHh89TJh8DFBCHbbuTMfJeVpRNCB5hTf1YB
6rgOmeRo7ACSy4zba6TWWAsgqmSO+dIuzhYn7k8n8rAIpMcQVufld1M2gTea
8NK84aHkfC5bHe5DN6VR7ozLtrNh3vkdxlJ8GuygiJwknfyhWueT+s1UcIUd
Sk2otkdJtsTLuM0bPZqwZQz5p98lxx9Yh0ZqaTbD7Ty4iWMouwqj51MrdUm2
MtH5u4vshw/mZngUVZQ2T1DEeAFpCdKMEPy+FoQ+QffU4M6j0OBc4QlJclU6
KGW21mdmNb1niygpHQq1CLu2FZoywF3u/iM8AI7ytjc0icu9rLNHFJVlVOgK
OGw59Y8++2CAAuaqY+0bQQXAEqzs2aT2mqE/3UCUk8CAPsgw8Gqy4DBq0mDY
FDAhTv+qQm+h+bL46GipAeA4ipt4SSnoke9JaplybfzBemWgXTscONZUE8Th
rqXD4Dm9GoGC1VucjsKTp1ItTuNyAGWYaADLjE7rkEjroQkURRi8IKaXsctO
kAwcCLagzN1m0NnSELMBebGzJjDMgdaYjb3RVq0+ACsZtX1uZ2TFBI4TSPuR
A1jKFD9+CQ3PIfiwCxXp193FOm40geki/tYxMYtZJ9GdFYwrp1plObm11SUI
NlruACrJTlcyfxWuV6ylGmoOJhejcSpJRpbk6eNdFOXlfDMittWREbrUGkC8
ZjnT6qbA0heYxAw2Knogy2uTwtKzouZlEK+AE16Mxa9rNflEz5gTqRFIV5xm
I3glAOWyfDcZTMzeM5ERbeVfcWzCLoK9PGOV8roDPzWCSk9icEAuprd6vYJZ
mn56rMZXSMuv4eQgBcKvXgUhvt5rksahlHtcv7sS47a50iqWSznwvNwH/sfT
r9qTSwjaMfeT679tnCsOqEwCdG7aEUAbLlpJWl2yqYfJ8pZXAhbM6p99pVQX
ivb6cd+xIBWAQZIt8Bq+C/BNZdZmp12qUp/Gg0NFZ4zpLyKfHFigFpquOZcl
pQIbcvplJidUN51QHZLUvWScoAsElIrlMI/CZKDdep5Y1uiqSlORkehGm2o7
7PqcatyedAgu+zjthk460fCNrORWq0BrcfOcDm4MQknZF3Sf/GUu+hiYhKVE
eMI4jPdP7qGEPyXgPrAf6Yp5gpeBYEvNN2E25Iq0kxIDUvDCZJIiakRdi4Lq
6qIUOINuGYahz3RLqAwSjwMo/8qf/2CVAK886/uNscOkLyuVeIa9A/Q6yV/d
uspJZbo0AGlkOka00/VAySSncqJoaFiP8LsoRuIrSfFFSqsgfvkfJAdD7ZEk
CyN2cl3mXSNcCbEju/FNvjasvD/+zIoKbib5sc7IJL4dDsr/WvestzxbPnP6
Mn3L1o9FUKWNpKexEh9u6Xelwex9XMfWstE8KednM4SnAdpysc3Dwu8mOwwL
RDXkdnfzSc45lKsTR4I9JRyJHz5L4+vC9HB6uzd/RdYT/W6iHHIQssEm7eOh
41rkMqSoQrH8MFXkxxu4qetNYeQuAXXqQQ8U4+Dt8Fvc4J93nn+SwC0OrEi4
s7EeK0AdP/wXEJ8UXtR+5BjCSxUdRnir5HN8mvcAf8Gi8WirBscDVteuM7Xx
gagsD0s236pVJ7xvuWoOjPT6XRO3qplXk+JY20fkaBhmkCl+eSLFemFs6KDq
tLYwO86iZCz1ziIJVqwC4AtaT/2xHwktkaVOcUfpnWFEs7ZVWtmYulxA1y6z
ezYBUVPY9mKh6C9jS2MrXHYXYo0yTnw1bclxqt2SGtVLjHqJBxwdKbvBfRPc
ftQNbYAXsRHakxkySdbzcysykaVQjcPP12uUkqhQY43bT3O1PTKO/nIrKY0x
Cn1qoX2V6RpFTUcHGrlWOjT5qRRNtux06YsSro1vEJ73B4Nw7tpzZQ37WWf0
6ZhxaJ0oqg7mhXy/

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q5MMsmE8c7uYGR752Kas88fOBzxxWA3kLtoe86Ab8LnANnMsPl1kGTYJoFODIbazNP3j87EEciLWqYBVY4A4T6jN8CkbF4I/5b9+HwxprxsxvqGivDCMPraHFhaIT8DL2IqSH/YhFOTZJzxvHyl9xbn5RJGVSmy/h+giYqNFlZS7hwshImUc4N0XvFoIYCnIJsAoc6D2LJZqluqPe7KFnWgC08AInsRmHlzxLKdlApb0MAypkDDIwxsqQeLlgvJEi11TiUliE4e/7abBApOLOwo74i3852lMvefwz6zfZX9wjAOGI6Hd9sikFZoRm+xRXhUfDFmGUDhBwdwQ+8qEpFIXDnK7WGB2oD70X5XoKIFglLhDv8qYW3qV9kCDQNqvQj/6lMhHmUt4/2H2s3d1RPjeAgUSsiGZayXEvo9MOVfxNDBsqlVZyboHJb0SCXiWGVPRBNK8WrFFAsZ+BgI5SXryBlb1HNUHXBqtKMB49LNP+gZQdnGTeWKHki3Fd2mOZqeAuX0Bbw1KfufA4+5RlPTtyMFA+HLRf1lOw2itYXP5KA4R6wyJzYK78AWrlK8lSZwUPlrPsVSuVxs7pOdYxqsmluKDSLEfG5AJpV48WNObgehrGWpb5sKIPaaxROXPqbSTn/iMmAeAm6++GSOWOc4zgVi0bUqO5WsT05zKdasJ6at7YpRmjZX/MTTu/Rsk/Eld66mzUjETPd/WmQYXQ0W/6SMlp8ytyG4EY43uwHtCyiD9CkUlzGzg7JwO7bvog1R0DlNW2dyWhF56x67YZVu"
`endif