//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WTEBmYMN8Oc35Qi/4s04fQRvAqYDvhlX7+A4bxY05GkxyHF3WeDIvKDvePXc
8w7Ky8/Umbp/jSc+B0WszQvyV0FQ/XwYo4DSqtkgRiwturu6PKIbw0ADecn7
mxWZgiCgRMdRl9yuM792dSMuhQ4hgaElpqgMrO8eiN2nrgJ7Jfl7UzYEiOVT
NEdHza8xijWdA+nK8tZipGI93k7M0/QdSMNGeHiLU6JnmQZm4fAZPsODJcSL
8ov2dQUHgeq3c5pyMap7n5iQCdJG4Hn4VuhbGtsTf2OMxZdlwb3p1slM9ju9
eq8j7tdBoAk6+Qj1xJOoCrBuwcsRzgmeSBk0d4SoNw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OYIuyDsmsPMVHGQWMK5dVExNo0rnap90TK+u68P+eiOgqUOt+v4PPWT/tGte
aWActWjzM4/1LFluDxUY+YWRDBGPqRSNmCJWFJeWon9hdJYiWTJ6Hroz0D97
IYIBy9FinTeMzRwFoTiHvvafhY1dsFJa0Mz5iPQ6nu9+hvfLD8OfvY6C5L8s
lzcsZ0HrtN5DTs2+mb8JaIkwgjVIiIUBy9x+rno1Y6hlwSDV3XfqDGMb47/G
llaq+ch80BowZJCvCcOak3Di4MNuKOCsaSBrWQCMmSuNkA4sOCsbwvRLPsCr
swB0xCfTHFb+D0AN0e+z46VIpiboki3GJcBcvbKndg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HRTKYKuBTcCTNaJ2vmlC8/BsiIXJjl/9AoRIwPAyfRzke/7a/XfnpwxfT1r1
/O1p5ASILZqlaKd8xcBxZec+hvok3jXdkoIkHZTK/OFLky4x7h4xSBtCeF+5
UYWb8s7pysCTvyzHfwBHSl7BsxIleiHt6iXP8dpFVWOFAnIeLt+77S14fyQk
6Z0hAX/FDb/8R7cd2QCKa5TcjDOBWPdbCPeeOydu6i2625WQAiijGv5h0d60
anfSDHJG/stGG2lV/rOjaveLQNv7ySkvNbIbV8sqbT2VRylX2IQqb5SmI0Nt
dY4V8fSJ3+CXk3KXcN5RD3t9DkdeQ405QThm13cn1Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
sVWezz85FACFwG0faKuM/ViHcKsC0500tI27jlbqg5SeIpCQBm99Sw9a2wcb
kwOVU6nv0I8n27zXAmU2CVL5vp5V8Syhk9fMsjzObaKQSynVc9R19ncVxK/Y
jTNwJtHMqyk9i00UhRct42+G8LLbSHK2fhtUug0rNQpE/9e4gFM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mmCvvaJr8HwWegPC2JEDIyRihMsgvuGYaKIjGxstip3GI1CDJeYOPSdBz/Wk
D+VI0Kls/if9aLpnVPgZbdoNb40FmAnEQo8FTQBMJzdQ3bDHSbf/fsktRIEO
w0UvouOSQH0jdHFN6tKgSOq5UDCt4rNKRynA0gleceNkw4UygtZsuqzvsgmC
WEIcDDg21K+WVJ4T9zPfKFRJshHu/XnOfCyEEr5ifbLGEXOA+mg0JOSwRhoz
haxy7WuHa/TfnHhEvYk93MvsNJwIF5y7xwLaP1Efuv++f6iCe526jHekRHzK
iPeXtkVKX19VaT6XiCOU8oENGPF7FiFY4KJsRufvGe6GDnfeHDy4e7dRaXTh
zldlaclTjLgVjq1PwmnGRFIR54fTLTl+TZiRfsN+lMNLEQyv/7hrF1HyU46t
snwb/TpifuJPMEO6LxkCwX1r61rIETpZl3EWQKWEN86mJMU/7RRjDYn8JX2j
mf1sLelFlUheaR4aPZatPpf0jw7NYgpv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ko/95L+pjaKLUX2hy7QUfgBzzsG7vmTj4aSXAKjASREw4aQ7JXDNrzhWIFjm
YNEEfiskUYLJXsSL9ZWqFdkRCjR4dieuwOE7PL5dec4NzfyExwjyed4D1wAa
Vn2qs5NGpKvfTE3SP7O6EV2Qw1fqnK/2xBSIClzcJ7ecP7pAhsI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KkHEPl3kC/wUEF18eHJS0WcXyVX+fCnZTPA473teDZfq+DYfKOxPxdqJNf0o
dx11tlw2JASCfUojwxpB8PSv1EONP0j4qyUt6V4j1mXLE2v31LxM9USTXrXo
ZZBF57e5S0oErM23mqahl6tZ/UtX6JNmJ/yCavFtX3QxaiC85DM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46864)
`pragma protect data_block
cBTQeEtLhyM6cy6nlNcw61B5gj+xfwtRtJ1LDWpXzBYgZutYtdKBnScMpajT
hHa/tSUnWrTEDMQFiskQRZ+630XX6KfTZ+9yUleNswfXDoyb11wBvx6DHioW
i9HqK0R/5Cw8WVUL26Mv1AQd/07xeC0ZSAujZwY00nSdj/OcJhWBij0/IziD
qyW7znyPqpay2e0UhYNoyx8sIL2KukJVLMMOSqo5ZgEeW9+Zz1+r54yVV0kd
EX7pyqqjqGzx7zmqvjgdDuKz989JpR1ZEnKUr6e8wW40FtzodOYkvKedKOOU
EWjhkQL5d9CT/58sjYZEwCvgKfDq/I4NeCLkareDU6MwAzl2jCkLj5eA0FUj
LT76S/PH9EeRZhY3r7XrqucYugv0hfFhn5ziK5CeL76omEJU+8q3Z4bCPp2a
oOio4BcfdyksMUnUDEYpnBkpL8rZXpd45smP/DeGv/7u7QjrRP/OZJrDkPvW
Op7e49iwWc8JDRnpuA06Q/jm8WEtspG/5IACtjyoZlIkRJ3Ly1bSO5lFXC0v
vIkp0FePO0G+wHgxy3IJW47QNvAZOlp9o+H4z/kzcrVKGKpnXnNgaS3KwUQB
Bceowa/Qp7tPMVBDR0OAM56P8uRNrmZLbpGFGLEoabTcLFXTFNVfkKRUKlNR
UaG0ivdcyWqAW7C8Mf6TEnrQQc/NK5zIiALrHh9MG9571vY2XyCFiC4BRcZa
nP/WTHztzfuvDb8n14ZHP2+CFKxkTqajxgw+GkFZOc5yia4l136t+Iv/qIHS
oeBkG1Ik3+6NR8zuK1sHWDyv5roP80/g5cLagg0/mZYo/PtjVYt1Boh2D8uk
waHToly7/HsSvpLmJea1RPjM1Rrq1ScAJcajSWGjTWgpkBV3qCJ45JCvcIWh
8OpnUTEV8ebCA+HYF2i6s9tb++1BehyuIVa+yEDdSlBYyUqitTuXJ8evQHnF
VRN2BBwIGPBL7QtCHgfTvLNc2YXjNRugZJ/VvcVRrCzJXrN9cV2tgZQMLF3G
u3XFcepPeJDr3RRGXAGz6UQUQZTNvB4ca56sLe9hyNuWYvoBKghkqG25IaIO
60AiNcgGLGdUXnhZ6yCCdwaT6aVBTMmo/3aeJSZZvUpCcH7Q2z6cffRlB2rS
GreC3V9BUUxME/Ao+ncdN6gMKvr9+Swr9qKuQGiFCsyoVLpcNprsnIrxIXSd
izMLzc8gE1mYk/VkBRtfKjxZ/l45T047QgP2UhIelIrrhn/m0Ux/3FiGG4an
KmxkT7jgRT3oXiMcMwnbSozZgzpxdiJXQ5MOcDI8ZQN2VEl2BpllSH9nTglT
xuC89/FI3tl+K5gx+LCzfcWtcqAEGXW13+tAHGFiPzbeKfQLIr8C6LmI/J0H
nilDEsEx2UkSDhOup9QTd1EKZ14jdkyCwzEDwH0W1W8VQLZQtSt760Apj7H4
bNC2dxkr+dGjDYgB4ooqX6J2SvBz9BedzTV6w9YzQun4WYqVDYog6ELEE1Zu
dwH3HqHTWWssM6aiOgkkAQiA5RzWVxgHvidqYc5ZpRM46pYy2rLFPr9IkJu+
dvQjx75VHzeklCMGQkp8bjDui4JMxz6zaKvNKvRKuS/dWCdaR5k4dZXxCj1U
z9PBr5rTeWVO/EE6E50pDA7ftgeGECzSjyVnKo/cTvGabf9SW/+cwpB18tnf
DhKkGjjStHBuf9UUdSU2aQgCEpAnQeEP7YuWqw2JiKliWvOe/4Z7P1ZyaghV
TsxF+dpoAI5dkrUcN3jd3w/gaF7I91QC6zhV+bJNe8toDXIw9xwRUnxAbgzz
ZhKsxHx6kgRbCjHmWYjDQrEtXLqEclwTtPkFkPiglcXY/k8C6X5gHuPcojIP
B4uLuveZATAJe6YiE1JAk1WlK4XyB6rlCpmQQHoIpbIQAWZFc/wrvt5tlWGN
3YeTZQINZfnOGSOdWuGq/H7VVOVRKKYt3oHcps3ieXfCgmnyuOzkhXwb01cn
xc71wtyGNoMcA00ATrZOzcRa7vq7RyiSsSopeyAjmDU0Ezwn7gFkCKyAlzd4
kfqEuH92JPLjkQZFT7sE8QaCPlzmLikmiAo0gdzdsrMtB7QS/Seu+4YdqYs3
wEPmEFAFC2SrC9I1zP8IRxsz1R7Qw5nPCvirBjqQwCdnI2zd7S5azWhbdAjA
DMuMkv5RnPwoGfQrFYG5Jc2ZyZ6ru/EmiPsWbUExACxglXQWqD/CEhkgBrxw
R6bGUcZwnIxae66bosCpA9G34sqvu++naoBWPlMSz8+HZUpZbDYZVPjZY+QZ
Yp1dObpXBzeFd5QsaTIuwMDBD7LLt4pSe4BNEaCoX9MApoyY6qQ1DHq/ept+
rQcg4o5YK8H/R1jEd0tF/GacZb1BU+dQAu8e5K3yqUUzVEWWBwxY2vO40xWD
Q567WYWFn7wjvI4XPTMrGQ1CkA643evB0bXuFePZKMcka+ExJv2gH50x3/2i
o9wZIXO09lVnV+VOhkWIeZMjrD/+tdz/AicThIqNCcyI3hfFby4L6Y2rt+BW
2CHj6rz856LrS1OMJp+1oj2C/9WvkShUIQIEeqFwCGKQDFM1LiS7iDFhfeM/
+U27syQaTuVtAw2D4sgDinWAMU/4C4CVZpQ9uiAKhImNoCB0UNVRtwciCMUx
3UInik6mNdejT3dOwcU3k7oBAo2c9pWV1Q4ibE7iWnF96aixLTo8o0cnlCVm
G0BXCcMZtWlwNjyVovk5RRG9tBAMnb8AGeCJ6I4+3jHI5VoEVSh1IrB2hdkE
BkNoW1b/Ghk6sBKcXkIZ/8xku6JnLnaRFJSqMsrpryGGRrF2msI8WDuqtYBR
8U9o8VvscWvDx8g8XNIjkAiFbVmYqo3Svv8KPqPUBZqUItirI5goOnTinLJl
tDAngJJkposJBneaQUWDbMa+WFqUrFGYvYZVxGoHusIbXvibA0N7M9jbCaXY
YXueXcAiFnEMw27WtLo1g2qB8RGBog9Dr2IMvlgAU9ThCLNOuMn+8IBgLZA9
9wo3IEiPY+a/4EU+g2LYW/Le8XS1B13sap0A5n+Hfc15YaAaZjkolqggSmb0
nnNPMew+ZShrLU5zd0irVSsqynbLTyQjWcmlGnE7IOyAUoe751Vfa40xm4+h
uf5FIBKCUGdjfC+I06PY05Emtnju0wtfVYP9FFnma7XX5M3DbL37YMDw9oN5
ZqXuUi7QvX/CjiDIqPbIglz1USaDO0I9QrqRNn8mg6UwRmJhP26BSJ/Xgr6W
muw73ViMKC+iy1Wg4d0tMsWFvnHzQ5++NvJb0iZMiJ8H3KD7aH/rEcC6ixWt
vY+aa5mLHU0iJbq7LoguwByXXZOMtuDHjpC3C0uZex/qitiPOld+zfAvOo8R
bgLXVJivrnvoAJpZd6m3Yyig7wpV1uwdphFAKZzL228nMHlUJ9XgPRWqfvh8
B5I8EAYUma7LuHQKEEY0bDXpgYOpSICs/NUyydlDsFpuyokaG1hCl1leX1pk
+bcgMIVHKx2FlRCyMXVZeWSPtUHOQbxPk1vjv8Lo47hcMg70YgVkfoE5Ccq7
8PFmh0mJZ+eCAbZ2yQS+/p52ARil+aDpJcX8vGtXuGOxXO/HcQZ5HjBwtd2F
Mdk8YBii/ZnQwqhYjLOv8ye6WUk+gSWH4OCx/HzYg/GkitE53Hi39rqYvKAC
galcqmfIEMqDPtypJy4lyfcW0VM+3jIr0rdtn3MPIK7t7hiifLKV5MzkgRke
cclk0zaYEU1MEA4xpvbuGh/UTmddasvpn/DBMf4jPhMkKkh44Fed9ciLoAvX
iGaOBHOLnR57e6/HumDreB6LBPhRfu/gZ7S3aOxE9HVlhwRrCu86jX2UFaYy
T9bmeQfDH7O9JTwp5LBJnlplg/49BBChfa+/fG3EnVvdyrWcQYbBuTMTEsJU
JXe728LFnJxkou0MVOvOBTiKSm6qSYBwKtjKavJzo1vSwn6bWqu4F60yFkmT
iwf9fRbOXRORX4cpB5P3s4E/NHNSDTkd5AnCk8kY76HQr6DguSjvNY5oy5Cl
o0YK3Rvu79OD8KwSIvLVTQi91RBrDyezNyXkyGg+a6CF1IvBqDbcwbqEFUpK
yDUuKlxIdlgWQ+y6sJ8r8SVgP05DNBIVEb/2vBXzgN5qgbo7uTKTxHA93KoA
iTmh0k0VFXEZHfiA5AhX10Ejat5DE/55cDhap8lY2jv9q4F3PROtdn121R0u
MjvCN/cF7vDRE5ncub7tInUzEZR+BSXUgcIjtb4L2WNQQtXXWQ6V4eKFAl4B
Ddw09toYIUFBn4OGs6aOB5dQn/pZ1GEdxFl1mkhhWXGU8Mi+jjqCinv3t9Nf
4jxctMEi7nPxRkv7418KoXZXIG6ONy0POfj+wPo8/uGdLNTUwQxyW2QxcPPq
2wsZS5FTx6Z7pPqYYR0CNEidxM1udoXPLg3yOuo5HQPZkYE4FOKhI2Fg8ZcZ
0poTDg+MkeJP+vsyyz2zCSR6Dh9CyTbf3D+pK1FEvfn4ZRARjDNn1jxLtMKv
x4Z3XAYgunIrElZEzJyva4Bbu0W/QATSzn4bQyt6KsB/2ih/m8+JKmc9Ov4b
S7BUdPeX3HQjAQJRM2Sq+AB3yXiXD1CVVUTrz/zrmdY1HywkIQMRr1QDN1ub
h9cBMAEBdbOAiBDUmmt7SDA11JX4zduTT2Gy3/pnLnFnTIcO1OulPXoPT1G5
ksTSjPHnkn7nrgEtCpRELnw+2oxel2J2eMNAsWT9JR0m+vQqj6ftmKBpdziT
Imbv8ibv7BzoBdAEos4qJTLe5eK2hxEFNYhPhP+D4DLp8nP+Y5ESizHiovv5
t8NiPoFwCehZeewfPidJWdPJJW6CETg+zS57b3DzSFaX19JbqBOy3SsTC2Av
bARo0OnKjYDvK7X2FJxaT9/HpqW2bDBSJp//FRYJTADg7dycIHC9un776lGY
uJgr9hb4hrIp6g2qxVJU5fJ/17b6xe6tjc0Aoi/lxhpXN8wNBDNR5pztSaGu
2obmQVxzNNgV/aV9U7u+lCKEs0mC95JLwv8WYDNo80ky4nCh2nWOHKxPTBr1
9jsmOEfWsvIqL9pug93P8nOmsiQ1zhOQPdjeTAuRd0aV7uztQnMI70EsmhHJ
9EMoIftvblixUWx1JwHD9nvT5lphxD1R2087B5zwp/HKZUJnamrHBYDHfRVI
+cOv2nfR7NGxoKTqf3zwsf1KFSFIGOdkGkRoaVsJEbJoCn3RyqMJUUIejTS5
72zQ4GatZ3v1+5MkTW+Lh05usPrmoTn84l0rle13+7DlX2wUkGNBkHyQIYn1
QSlZCa8+j4BXZjFDUpsRrLwlVDcatW8j1WbBc8pq04HNrUG5dPk0IxYVTzQS
Pzstm21f7h1xqQe/wE6oqYKJOuWGecd3Jx3AqdQT6h6JKn6OHqNSUMa610Ca
1oAsYo57D566c8DrFf1eHtcA+9qcVgW2rQqwnQG8YeKhOYJ+nknhKgh0dwqE
KygUv6KqDkNmnW8s0pNaAUlJZjbQZau1ZmikhYHi3b1RTqpW4oDy4YDn4VWf
QNqimH51SpqqHTGUnJH5zvF/SZrZdkqKF90jS6kOl3hIlOaTlLTHh381qL8L
tbMN62NS3da4/tZTRzsXEcGijJADM/5OaZ/FkS85Faz+jc4/zjvA93tJiqaZ
gVwglfr+QUVAVO6cN0Vmr9xBVjt6bpN2Ciuc5Yfi55yXoHaANB0EsxJClNV7
1GK112GrD+s6/7CClcMF0K8W2ftKe06YUuN8bVds9aadNCsu2mVrWVTtgcuU
aagUQv6s3BoZGwh1U4XJBW2VcMvxZZe1BSb5Hak7TbZVJ2VYl0p3HG27M3iv
G0C3TnNiypJTMGX9Agmfn7F9k217FARe1kixPelo6+Xn0SzyHqnsogBykymW
6yPB1rjrmLx3Sek5fK21rSiJa2hdCLsDzbitqVOigpA/1iS25bszXoqhzX4m
1hV1fML07fTS+oiuTybHWuFrJdgJo2t1UbFhajbhCZhzid8TblLvGdUKBOcZ
XAr/zEPbimPeNy8ce2qhaCwYHPmUbx3azTS45WIn1+eHyaKPWwWWbM57nAho
Fiyjfi+Zm/AITXlHLPubqnISzIh+4LIZM5LLjnwTnYAdNcKrIcAQv2jDMEcT
/+zOD5xw9FGtBCJOjx65cwtGa9K0HSxSY3xKN7QELQigiNj/LpqAY1sCF9nL
t7XViAI2K9palElzj1t/BL0E9eP9P7kdQ/akIGTrUrSqMBspZFQq3KcYu7TW
GR5fjejQionkcJPGV3HmSd6sb9GNFye0zz3cdswJ7Ij25hduDFucjmzXR7nD
xSbWZhsMMBL51BvyGFWv0SA7Sp+ybe4TeA69U2Gk4WV851LKORjYcbhP3jbl
4CHGmWf+7J6Fb0WkmMYmQuixYvlr5K664qE8kpq6VtvCD55NZrB9DLvvEoq1
L90Ij1/FI57DAsDJOlVKHiXA1T6hksQHXAWHL8PnC+gKfBKT1Np8z7yw5lgh
RDZQFbQRcKoPsiV7mzE9FDVViqQGpxTFJ+tyFR10VMnuHbkSUmFaymeoHrKN
at9fv0RuK/64fy5jiGxwjsKNahfgQmUawlPHmYUk0OFehbzlGJDHwBJQ9bLm
PDSrqLLi0XbRyY2yTnqitVHI6d4YqU/EjP5Msh/w2xxPX+W1PX9kCa4GuYyr
eF58/pz9oItir6/8y9qhDhr5IyZt/+ojxkmdiQF9J4CnM2oe372uAu/31M+o
dV2mTIG9LsvSBr3IeWVWBD7ih3vAuU2aXoE75s0GimSueAAze0Djac6lgO9H
TK3q80s9oERVCXyYnaj4PY+7go129vU1LpmqSQiKob3ZRgbz7szkOvKbeaPc
axZYKayKfnhOGcQ21LCEwWH1hSEjtNSmHCX+8IJODDRuntD5Pkw2FfSQAa+6
TAbVjvABg+MQxpASTWqIrPcfveyZYGeFEyCLQBucyC0X9fAIBw4y+XYGoQIR
U9oCDlv6pPejAxsqZ5FDTwegnU2kUpEqQ5cMkUWWKQprWIGv2sR6Prb1HS46
BN0eu3KN5ODquMLGfZ9nXAXXVosBNLxm8ynBrqXaoYdGWcRiwtV2sf6CTZSc
gK+rVIM/dboeNzhC2R5Hrp1iXRg9pFu8FVZlj9DoDY7UgWRX05c2pc6YTVAl
FIdjKStsZExTDt/ykWqNlx8YF0jqRZDr4GGuyrV4tVeSja8ZZjIY18MHK+Dg
p1Fn1NxnBOyeoaB3cVo2yYvESwrmUALtD5UlLVof9+xpr/SC2eQZQIeo0DUD
jXbap0ySP0GxbkELWSCb+GqzCfYoEdz19nuYlWqfS6PfcknEsY044IhlpnAM
h8siETxvYne/XeJ14nCvlW5XCTd7dmJwEwpvgdVUvoH4XmaPz7MtiMmYOzCY
jvpZOxtUz1x0qMFDqd9zM6Xmo/4DGht4pS09PoBIrvy/zIUprWAbgg1U3hME
qinDfW6kiDDVRxmjXBJNrNKZXsTgkmcdhNWZF4TLe6IdyTNDG86cEZactk2v
vvP4EE7vUmyFLnAcPRUlBb9aqEDJmSq1iVDfaXyzaRXIcWrNVhRq7KwcylCc
SC49N6DqgULglMsiobovJKxSUEhirx1xVEUhbxsVUJzWnMIAVavu61YSJmLv
DLpWOV9mj/W7e5hUit6u+7ND7tTH75EKMznCJQmQcHcsLRCh72YjFKhKO2qc
gtmd7oZAcDfThq9xjYJlBmcLVPH2pBQxJ5FErDiY/+Xi3x6kwV1LgnYpTVxW
NWmBsEs26gXTuP8x08vvZLRvpL+n6tq9wd5G0/h3lTT7VMoV9RMz7cb02MCg
GssW4+SmiqT3i0FNrImwszeSU3R+ortcZy2BHmwiM6LV0Kwe24lHvHoZUR/o
w3w/U3wLSyFC+YuyVxlXmacbsKLf0grSRA+CV2XyXiFe/ZddN8ASTVNN+Yvm
cjPWZX3656pEPq77DqtjOR3103TVSNI6qVpdK1dfKE1B5vQB4Bpmsa15iIyY
UEpILF5mGjB2bC5KiKP5JktUiFNWqKnnlEItKVKJl7lYyZeYUb4W4yjBsQKD
wwbFRXmNRrFqSGuaoceI+NI6PNTPqRasVHelMhul64yzb75i7DgUoMn6qlpc
eWIrGJEYwjBYdh00wxPfhbUL/AjeqK552FTgGVWrKDqfZ9FeGHrE16G8gUSJ
hhFIoO+CT3SpVdt6001d7s0urK+wFkmKqeYroFrdLyf6EBfd1oEpPQZ9SZjZ
/nhDEBCF2G16hG43W1G3oYp6h59vTdn6Xa/JdlZFA6TqOZFze+1VS5+I5cYV
LbBmPmM6XbtPrDB9zuMbKCvn/iqb4i54V/zFAI+8pLUNwBJ8TRzPJ5Znh1at
aQsDPN6FUPbFJL/NTnDsnsy0Jqz1tPx1um+r4Kurt5w2FBi0TdIOAi8t6lzB
gfUcZ7vqKB3ktGxyt4ZKbwRSxSCUzSSf7v+2tRoPX2+MEsXS8iKnEY7Rol7T
HBsyxDCN8Vyv0OODeuLTuX8QYytviQQQB6c/M1Kegc7ZEmiKoXiCMWe3YsP+
suQOI3BxqWE4LkqOBDVjirZIHf/J8WihfqcJdFigCPQHObro8tV4j/vm1OQI
lBLyYs+OzOu40FHivROF2QlfixBoqKh2L6xRNMQahnZdDj2gKd3g+nmDDJnm
U3dZgS/KNgvMAZSR5yiq9A3ocvKAqhz7+UJxjCqQzX4nEgsSX67zrBqwFuS/
Q6VftTYDDBfByGAMacUET9R5itCaVkfPaRLLPSnxDYdyvNs8X8s39op3S0C6
zUpGCuLA3ZoTIil3UuPpsAw5d8qmdfWTjg44Mep/qvDsz+Cw0ILS+3Va5bj4
EzMUPOPZuXExtGdD1srbcFwMY09wc2lK/FWVSmFapuwqJnzKRJdejvSFV3Yn
5Ta3qToCBf+jWXRPpOn5+s7XkZTpcQmEeczcWbiMnn0q6+3h28gtC6sK4aB5
sSfAtPO12j9rz/5isaZs58DIU7Evz15amd/xEg5BvrBMISL5GM2kE/Po5qM+
iwJcbeavQ45426P3azCJxKfF/e9rMHBr2voHCl3X7pvk8I8e3mknISpfNj6X
k8eIhCjAZfdWpsMCaf0vNgLnNqCrCDtnJvpYlnH27ZaLZDO2zjtntTaBfBh2
FAsSthRSzQUf4+Hr2QKnfZZI5wm9im3x/1Ia+cp5aOhDUyVEuSabJa+eYnqg
ge9HukvZVsA3uhynL+GMu/W1qMHuIyWLI06+AiY3iYdmy/xpR6L9FhJ45X+7
p4bklaZnwVXR7ogxarocDWl4CuM7HLpJMBr3Ga3NMgcpetJPWz5sNEfo2BzB
6KBbBC33pZ6sJjW/Qhf5Hqm9RQ7Ll6DGuAkIexfPObYOBlhJl64Waf+zvKu3
cD5vnCKoR9GibZhm0qHCDLaiKyNaWRws3Xn+F7SIXOS3caadUP8ithdkGAdU
5UFvvaSMOTTe/VzUbSfFgdzPGWJ7qq0GjHkbwDO8M5r8X1AP4/GpnDDe99zH
kZfH4pxT0DE2fGgrwczBv7BbEzWQn0VBOazHdDWs0Kc+0E6RULbHuHl6IM5W
88LiAWwZx1h/yvoYzupeuRZBZktCLX/tj8fgwpNQeMk0QN4zTb7XJ4QLj5bi
r24KLm+HH4XKZ6ZaHDd4EXIF4D50FR0r8zDoDFAnxKzWqkZijNzLPzcIfVoZ
1xsorW9aZMnoWOlFNRkO27wh9tp3l+rNUVOtsveaceXtnX5UxsrapLmFuXbu
WmdR5aYYOaL0M8elRr8EumBeiVSR0dGZzeZikRX08bilMK2D7MmWOeA4Hicw
/qlMM5rjTehzQ+Cf7KEyT+l1t7sjggaJjHLKk0GdbKucKSSFpwC+COyLPfzu
wPVKpnMGfwOMpqd607lP2nyf2y8Tr9rH/Le7ZAxD7bNac/b2jbjrwGE+e8t4
SEVMTCxjffAd3R0L3OZEHWzKTLRwJxI1GKXC3/UOwv48pcX5LdpW84vICq90
hzyY2EWZrQoQDlC1SKVyk6kX7gwRv/GJZof6dZMpintjqHSqMXAIkPBzRNvr
5MeU5foy57CEIQtYsUI0bNHjBO1dYi4Aea6otn/IYltHlIBCGM0BUEaq3FKx
Vvzf3Q5yW3h+rTi9ValWPM4FYCdRVKtt9lJ4LLbvCMzpfgY2HSUNhNkluMQj
eYgEQwbcxxpmmmGwE+3xgvyGqCK+1subxK5/mWcaP+fkt+3L4dkgUBIFAicw
8rlufxhjiBQ4E0Ri41fX5paPU8Hl2CxhSicFAzPfOtUUIM/SYQ0PTgHmSpJM
gF6qIboyWxBLH+eBKrCAMFupJLZj3yZTIR5V7BEv/1lQyKx7Y747Zb5krK/e
PI9RPh/mzq/doTAkGgej/0CdFFmOvEsB5VtPU9Ud0d4Ok8utpbNQH+js6VEn
jWi6ESG38qMDSOlTdS8T3vkwn6qrDYh3Rg7vWra+qIySC1dyxtd/mVXIuUaJ
BsjO7ioyDN09TD/CYmKQlXTwBzx2AqmPul4x6HuSqYZm3Hp5NFePhO52DoIh
OGqkl0A/k73Wk+29kqNzfTtTcCbn5ltrWQX09rPXuq1K41jRBllz88wjSLLh
V/gcpgLkx0UkTA1leruP3ByACjF92YVtZAz5dqvGVpxmpXSCLH3QOBYf5Tl8
gUyuUu6VjkdqyvYcYlST2cC2Qke+opwssBrI0X+R6rTOCAKaTmMV8mhqlIho
EEk478QAScpYP/N9JBvt9tOhe3n4l3eMRMH7ayfdt9paRz00qIG/wy/+s2kU
8rfIBfm+uaDxUNlKAgatab5vFvFoOOB2CcfNPaofUsOmIq+3Jyb9MOitA45E
gTSaWfHUiNno6ED+gGYJRscQY1lqx7W4O4SckysgH8Bdw+9VwzBvtzcOk5gx
kb2Mf9adLvkWCRhFDBbXHe1O36WJef07A1yaGw1f8zmIgbW4/D6RSyTYSIcL
g5mg+o9G9MKu29Zxeojpv1LMWm+RBDU109RZOm9fE0mCi/sF/fC+3mJ/ekcs
X1ezhSowjVTpIHI4LkAPvmRpvmsCS686kh++NLgY7MhYd8Wp/vtVrLHZ1sYF
W8i5pC+qAWkWWFApaqOSRPQFpOKoCAKDm1g73cEyeI9UeGJMysp2kuqgYJIA
DHzmcRPT0VwVBVIYi4ExcWq0ajDItiWxaJZdHkU4UHFHh3Lca2CN1Uq6p4oZ
vBdPv289Ifi1+ClMiDSYF2BdMBQ4fh32zCP0NOpPXsPYry9ymvi8xlXSNkKe
Cnl7wnV8MduFqAjLkvi4R3OowZ/A8XhGroAeNOjwTH6P+o02mwkQRFORGJ6/
pDchPYZtJm7q1OljC1eRRzHzOxAtfd4/VAXk/JZG40SAEuOKyuM+FpL6Gx/O
tRVc2xkDXWQOnIyT5lZQX/fZWXALFf+YU5gHuSWLfxgjPSJBvaooyo6D1J4d
6xtjEEhXwexA9ks58BJrbkg5aCPXFh2OjGHBtVREhMU/enQrNQJ+eNM0UW4L
eXYiXx8TbeOu1xhJE1bBdqDovH1tYItbYBwlZBSkyLm8EeOSuQRbCn6RumvA
B3/66qGRP5fdN/juPiHEdK3b3oDewvcMgqDfPFE8fVncz+X7SQ4mUAnFlHz1
1QiM0IvsTrXiN9od0BvOsGadWj5WGoaQKVqYESt1c+7Sgb/eyUHq8gnYoBV0
hIJT7gUT5iL38V+YcNr4X5r1NpgkhtIPoPvQvmvjrR3dsPxOeGususqM/FPr
tCS8KDaeHigDjwzf3wt3850Gh+LJvFAFNgyGCki7BigATgg18gJDymHNzenA
09YGx3/zVKtjU/T4nF+dNDwigqeNrw0n9MwvIWH3rSKFy3FAx+iSm5JYBANY
4kYDJAoy2C9S41amNTICvhaPJiF7A3uUO9+A17kxuC1bZ33jjGXb19HcZu/h
D7IzApEfQsYG6ESWg+8fArUIdThWkiNQRU4laXK1ZsP0atvp0jgBdfy980Cq
AODy5M9jI/i5oUQmJoXiXFto8/OMbsFBJ/lxkeCKANCghxMo0oEa8Q90eLUq
F0S2mVxFelGbZehaSTqz3OO2KL64r8e44igZlAFNPM7ANqw7fHB/hlmcWtXB
zD9hRj+fCT35qWeTV/Tx2vELg+rOIkREyj9F5G1BFbsF9oMd31qkSmdghsOO
LI/O7u95uEv3RssDsrtMiJTvD40nYl8RWGKSw++O3y+O9DWLRhcH9PsrgtxF
fpas+c1CkWnIEJ7rrapBEJbAQdkXsles7xb/eK1bnbhj5BzRqj064FFaCKbo
K00PgLYc7bXdTRQ6lQC3Z69QfykUZXiH68GKkj4DRljWEjF2rZgrPps4pp2t
4ZHgyeWJ0An2grinAUFqjSfRGPXVrb3/o8jrrkOBHY2I11W47rUnRHjuB2ho
s2qwKtBx+AP4TTa+w7RNEoctSZo7oZQEAN0v5NVzcnuOPgghXmPZ7vTpTMSH
CgkjNnU6KvU0G9WXm2wwD0cCaJbLxhC1GFZ168JLlIVGIJbXnAm7ihYc+cdZ
fauuC9z/5igBGSFSxds2jznos2sXgJYoQYmMoeZkkpyL7e0Sm3g8Wy0vzNez
v6Rcj1mjRTGWI6lhap+opO/nORAeGF/ZEvm47agZOTaBsAuYFmXi5W5vSvJI
t1bHwm/UWFSjquwDKGmVfITV2XzvUusUD2wMpcYlzKSS177+9A2sWleCmKbp
uQduxwlx1Wo8OEaf/oJJp7qdEMCGa1t0HY/69Fr9iFhFF9zoPZKn3fm9wfW5
dJ9lHZDJeCSIuRsXrRXuGAbrQPoyYSMhBXD5TcoJbcFpvXbSgRLZHIykNYNe
zOlFu8DEaWFs0T4ub0W2w2Ild+PBElGaMIbQwh5pFydnyQxywjoouULH5KN/
XjFBooBNkeseGf82Oikj/XfUo85AoKQhyRbg2IfVVX4iWGyef2FKZ8ZQhWBX
xksjTaKOl51jZvUSkygrf2xCDNmvSBBXOR0EssX5K4NHDT/X5WOyX5SXEXRs
3ByN5HtK8KP7BciIIIDBGG93jHEmrZ5yw5HyrGQJow+D97AL2aFHKpkMP4SH
yfsCxqiWkzsW3DZGQNPF6+Vfl9Z9FdFLFh3J+2G4VrkBg43N0e+Q89dZcroM
ONNHGIug8tGoPVIj0mM9UMV4cbKHAcNrmrZy6Vosyq7OcNFjpgNnOlFG/DMB
NSfa1OTIK22PeRZt/+lkg0n+Y9kZBdgTsciHpBllVyKkNfl3AiXfXtsGEyI3
vcpfmGlJEmzErscnHzXMZlig3oTr/arvA/3OlmefHJ8pSS01h/MITDa6oVes
eSij2fE2lDOtCycLci7lPH8/DpiQrZt5KApzW+5Bvj8SBMe55UhOk/sCKdoL
cjwpblDgNopwVELmyzEpIye9MhdDFSrElnRLm3SGc0/tSz7YawokAXszABUq
8Ou8ABLRUkLoo4VgyReC9BgIpz6a5OO0Rzuf7kM815yiYR/VTNfkzWVAkDzs
MIADrql/PEW+FCZEV82kycYFb7PSR2U3gVzmAxt/HYjfMyiqsbNmCGcHpQWU
yAgtBmSc8+6XXus4T69KVeOtGFrEHFSbMGv0E7TI3+mghwoQj6N020aPrrxU
Ct0r+We+HEQOmlR5hjL++11/rjF96NDi2C0jF5GzEn6aUEdQwohirNOVbGlX
00xBfQeem8eOqKiKfYQE2+9NVdx4AU5lOc1P8jpPuJ4XQLSyuLxDcU99jMDf
g24I6fnuNiQGSjfZiogvJRoDL3WuUiYQ5Po1WSfFfM1lV6UXmSD4g6h8t5h5
iJYB8lMHSwIB7Wl7Du2KPxuh8UMyPZlQZyefy8p5NbcPHHVyMj8WrObi5EfB
XHXIesdRvh74eFYRtxfPSZhzks0iTmqAAyL3Y/0F931UALgB+DgwgP4gyfNj
MGH1TJMr2I40w72aCUVJ/NCdEZ+J+f3ypSvbH8Jf8qXY1A+0bQweGhVah7qM
G57l19afJ8AaCIRwSsgjWPEq9nLtV6aLDeuJMbcpWzsKboiwFr3DuQ99SrxS
xu2TJctIyr/Ep81R9efCLzKPE4VnR3aDtqiiaFqYKB70oG7KlF2zzC4C//0v
NDL9WboW61M3aDklgdyVxa7pJsmLNN+Phcot2AeEDSKZP0Okmc7hdEWbAq6f
zHTyft/BQKwhaNFaErPfrYjXLWFkTakj2logurgI8g2ixRdaA/mfkolslRcr
NHTjKJLh47wA5mj+NZGSczGNLH05KpRwqJfHL1P5D9/A2hKchTeS4T8F6Ujb
TsBZrlnL/vYE9Q/uu/SIsjUikMuDe+Z0lOakuPmNmYDsOc+jAvPc8ldIRT3h
66kgUOTIYgwIYr+ogXxFo06JG+qiWpb5I/P7Jdx5LAtPmCoWiVaTeM10ojq0
YKS9eOV5AufO1e6TIvz+gkMZO4OxWV/GtVhfBeYgbfmj8Pm6zXOQe96r8WbJ
7JtkXbIrlZvarCJHkQkun70f4mxw50kxP9UK0F9DvLvukOCxLMSzJllRcYNA
1UgT+UwElXJvi8Ku2HgAcg2HcycLpa/BWFwVyBnyT2Fvuj0aLqp8RSNt4Pfj
1fTrAKmyd3LgBc9KNiQE9GQowp1DO9aSX4bfgsb/ej34PDePN1aj8PG+Xb+M
V/eoe00Twet9X+Upr9dhD5wuJsCiJQpkicTyDNMYtUIa2brT9hcJhzB3ek62
h2zkUsCJCmSLxFr7AbI/p2amzO4527pfdipyNn2hUM/VzvQAcMA3qs/wNNPE
pHP3U0jNxyv4qHIoRl+0ZwErrEt4B663yWaI9MjD8M9HyOK3J5k09WDQ2HCq
riWNdnMEQ6HP/Us2wi3/kMA+s6FMZxeqPxe4sb/FDNJ6QR9luZXf43cq3sR3
swKZUwFHLrbONulMRh8/5r6XlBusCHJBSPvnkJbWNbxt2XT9+YKODMbaN56D
ow3NPK181fyA+5IHemYJ2fdaB96VG3xj/CDAIO6DNdnfrdLvFL8hDBSN/z7P
fmAH5Rw3vO21FNwHz2NO2n4GOuKbMdksYZ9y/SAffRIXdWx/tEctz+Th7NaX
6tAv1lAmrk+Fbjoe1KLmyly3ryoRBJi9nn6yAD+ddHdr1T/w7G//DHZg2IEd
zC+O6Ox7tUKHD2jAV7hHgrGPTwfZvkeufDFcvvaHMvr55VajMFLnzll8dFfp
r2wPmc8YayCUIzhNybfn6Y9Mer6BBzqU7cubDCsCpH9V9vWQcvFNhtB+c6a2
AVwaIJNXNNpCOyWu/4ZpStM7TsUqe0TSGRKVm3gnmFkx/e2FBWK6AwfhFG42
ib0dSILsxKvW31l38J5LlSgos8T4rEPxF0ornCFQBiDMt8606E5esMlNBv10
nO3iEXl/qY71oLSM6kIWjwBSGA74jMJx1LlzR/HqbGAlLz0Zi2AP765C4b6o
DhfuzE9/pDV2PJsnKpUVpwpXFpC/boI80XgySeglA82em/OUURne02sXmgpU
GZPFweuUrSeTVrUNcQKSvSdSYVVozGVC/vWPSZpo85In4d7S6gXL7nlEsMDR
MAvuBvNmu/s9+FYKTGs9R5JFHCiUwFvHK0w5wu964N2ZbqquEqL0yHthS+tq
mgXERSQ/vw1NJktHqGVB/UGfHAJ898Z91zXQFPdApY8jGnJ/bTmF7rZaSlq8
NBgi2myBaor+2GD2qxVS+6T+/lF23HDs1tNXM1ZzXQhODrnVbNPFOjrm+VtK
EyiRhSZyiiHn3kNDV3oDqr0wCaILHVDmKraf6trgisp2OWevIL1Se5/ZHONk
raHeKqSVCnGeTz/OUIYEQlpQSrp9Xah/nV+NAhttZd2kd+bNV6fZd4wp7CIs
clH53Hn0plTQ0CQj5KKy3XX0WozLmiVfFvOrcjESkk4+nQQLomD78bRG3JOY
pG2nOeKc9Lq8gigftdk2P7x8F33hRttQmtVbgZwd1LZK6YHiySF6V066jpah
76jU7y+vu3CfA2HHPyhpbSbS7Va5Nc/WX0xBLAIhOHjz+HnxsRTMgenK0YzD
Bd20Kyz0mlhQgdYk28G6a9vaTNdaYlnWg3E9Wl2e/cDuzkIdWu/hy9RBVLzn
aFPAeMZPkxfr7SKzRGCmDCanhyVVRr0M9XNzC3NQm/AtPA7igCnTNjzbrwNU
ZzGoqRnyaYmEpnQ/uneSpsMpyHRoxkQX3kzIBe16gPOFVxqroSEadFxfXyXD
tT82Iydj4uMU7xvA4NFmq7wytYDaqHhANfkvfsiUVG3+eS/a7+3AQrlZ9Pmm
g7janL7P/6zxT/2v8d/P9o6ThoQ6X2h0pCxfDtxuQJVLhJaD+y3yNeMXMNo+
DmgTql2qRTtNuClFd04gmn0dDpndGls/55BqzGWWFel9mRRSGmbQgeLAQ6J4
qQMuFWs5Dq02v9n7u6K/DPqvO2C/DOVWhQYEQ1xmnDSm1XmGfg3Auo2EHt2p
JpFzhnBLchYTxRtPx99qs2nj9sRsKCPlMbEskXeHyY8/hzjosq8knxUvBYsA
jDVFt040RmN//DGnUI6FU96BzLuyaVe0QIbuPygALP/KP6XK7kyN2f63CUGR
Kn+P9YHGlux8J1nijUE5CVTedA5BjrGE+LytjnKZm1Up0cObvw51qIlocrmt
ore6use/8z1TXydQpbBk9fGEttDpK7jxU6lBEF5fp5RUVKxNdNEiAchq2sxo
Ro1blPdvNY+E3rsVaoF28oThLosvzTUUZiqVHMjUSqGRNP1H3bTzUpbmUJod
JOegz4P6uiH/lW44+Nq98n9aIDDQdwC4coAiNbCq+AuLoR0ZJlUgxjLnPCkJ
iTuHpR1Qo3Oe3cdYEYxb1aKls10KZrYn9tWysrznxFy5VnARpOrR00MNKedd
bWj/9PYcozha1aYT49InsBeXJfMQFaDZS8vsY6A+Flx/Rc6ZsfmiRjzwfGNk
o1mwNiPr3JCoFaqkUEjlyMIvCYSxOqcyMBQ7CkCzRrF10Ytme573NVVWybQw
C7HsXEVLbBnJIHzpwJFkrU2MB27SnGEO/9+AdVVmzdXEnvcaekTGsLlh5q/g
VZMTg50p/Zlual+aMSemrd9kBxzrNym9bzqX1yORDnkYsDRcbI5P62L0Xevz
ttoEzwODyFqJgNv3kq7ok0CfKeQo4dCbvzs4YkEEqDscQaUWfq4DqqL+UcxA
WG3dwvJGtkdQvP3CBbj1ITEuXMnNIVV389pw3BCr+8s3tGZpz0x5CympscvI
vSMwLZVTIuPWlnF7xT/D0xfoG+k/JbUH7SwCuCaRNOShK/WbYUAYmuvMRNPC
qKjYPDwUR77e6cMqbdb4lCo8INKc/uIw85c6HGZuYKsy0PBGfbCOt3Hgg6Rz
e0lroP9eRbqoPpCLDAsHBa7NFeNXaVH1HWSRLSahuF35Q2b3kFCLIc4EToPr
3/PkgWD6Apng9EguPIq7IRDF8jiXo8qeQuwxnl1itb3uclz/KVNnCoCY8wLB
iKAoRl3Is8pVvU5wc436VUqOMGLgwdLItF5A/y7olcubQD7w+aEhhJYdyUrw
mDEHRkcu/m5DyGSvjH1+haczWk3wsQQbPCUbs3kMoyPqxbDLOfT++14TbjgW
+wOxO3KIbjQ9J8Xl1zHqrVpwocNwBv++h2bMcF2MNBonm+lvfQ4AzSNVWhBi
zRltWIGredVvJ8dPTcfrBTI6hCJs/0s9vtM7b3y5ovvqHf80Bn9vUbXF16ct
qaIWUZNwxlIiO4oTZFu3JZ0Qo4Z4uum3rrTZrw5W1aKvtS49Ikpvhlvr7A6u
8P50puFtFH+fWIYQmZMOkxij1IlZXF6VeJb9BfFXsdgQxpVUM/xZn5dL2mV0
6BX1C7AHdDccxfx8FNGpcZkT7np9sPSYy7spDMPmhaXZ3j9YzwhT3xHJ7t4C
os3Ipmj4a34wZpeQ9LH1BGe0eoDrEgc7F2LQShRPe42jevhOfoyi7Ceylq/O
wizhDLnFACPLWM2ylQW+u4oSKay0CCKjh71qYqqSIHSfUZ3UxXJsgCdh7JlC
WxKTZdET3nGEtWZVTAiKS7gHc9628ic3HzW74Nb54lzksbZZmE9iA5ITh5vF
vg3WN/D3+a/MH0g5g/giX05IDYDSz0J7ecyp5AiKURkEZAccZdMBkP0T19JN
RXtrlcPWsmiwhEFFCU8zdW8eZAyMaZDFttL1UyGKUFFyfB7F4nVu5/KyDtx9
PG9dMluVN1n5QiIvgmAWgSuRPa6uZ7UtTl0s6YbYJgaAerRONlGkrFHJLhcg
oNCs5RU1GlsXCzcHTn3sMi+NjMR+XrlkbhExI4OM8noU+BSThgqENLcBuLqb
FAbPQYmctESWiN/QE5KUx4ajoSX/gqkiXxvIiBZBlG32869QpGiLs/oirz3C
s0zkC2+Nc3dgqvAXfHPATXtwJGnVda+VLgELAi5v/UzoO/ljCjLX3mL+fSIR
u3ReVi+6QjcS78dUWHDLSWG7Q9gJ9+Bk3GtZHvAJlFa95zMFPEP/9VM05lv5
nR+KbuvBfNq4xQPJNMCkH4ZaOFqs9/Rwd7e2jf1EMntxywrN52ixDo1jalK/
1nW1qWuFHk3ZD9x3Jqq5KxeB4AhW63476yE08OFiB5UBtBzg/7mSH+0Uj6v+
iydX5C6fFllprHKwI3YpS9vCqeTf0KSh8mTSZdLUIQne++Gvq+2iC/K55ePf
G7jxlIO4I000SXhhseAhC+9aq3eVShz+esUKVNkB18zhkTcxAgj0OJSbzpp0
95OAabWrPvg6lHOJSMHvYXxPYCOfdr0qj04iPIzamRoNN6RHLn85qUyIfXPe
vRJnevZggUUsYzTBw7Qi8Jy69ryaYPpwQyE+bmVhpl3awAmBWqjVu7k9CDq+
FH9acL7TKZsm8OxwbXxOFy3ML/hGAaWGCs+gzFPB+PZR3Z/Mo9UeAnS6GBty
UdcLWG6+7hEqGFFl0VuIYstBGE4Z24uIiB6E8tSbNX+nZw0+M3sqHK6WjzLU
xUOJU2z+anv1YWETI+lL5C2xvX2lsWC2+Jy3laS5fIr6DW9/SgiqbvxUhEWc
i+tMiIV/+7zSPi1dR3Rr5VyNuhoN1TZr0pqEkpnMNe9ZTHnLAH53Vbo+m2pP
Z63aFzgaf04S7oFVmwoauSAWyIRva+cd8oqUvJqNMi+kpeRETwADPe95VaIT
71rSh3xerpdYg136ziyJp57ttNt2dZSl5okumAkprMWqsjNxLPhkk616Pqjm
KIMPtDuehIrbX+eUiGryhyS48zrCXSJV6c8/qi0Rpf6VJNYZlywHw+CGepgl
08d7313W3zZemvDjHvt0obpIzrUMEfFmVZzL0sM/lt1GtJhPQctqucfo3Vz2
hdiPIbJpyAnu4MBjn3vmfsmpJcYNHU2csV0HXGt24pqe0lGqLKV7Xb9Iaip+
ArhTrvV7CfWWCHeFtc+1XLs1hu5NERH5BpnVuZmzYDcZr6+og81DTyhOVapK
dLEktnnl0mbkizg6U7PqtkzdR2e3Ix5ElDpkEyesZwCpHBIBDjpIxAyeTtn9
4xpERmcJgXn/+E4IYwm7k1SCLp3sbCVwD+vJx+xhnDEo6Rzfe1bu43UU7DTK
rNLPv1MQLMGuIVDNaTjJtItaVBmGw31jocq5yD2+fIBF/SnHkGmnfZ1vcVB0
SJ4ga9RTZvFcqREW3MjZ/XmxF1ycdLNOPWRTK1bkZ/zWL20FFL9cpSO+qIw+
9Ytd2fireQjHYbplJJcg/IEf29i+18zvFaAsMYRjxq4p/PMJD60Mq91WItZG
NNjuc2hUfmOG8XE6jhsS/3jV+OhsA7QoUlUULAwAX4wGgT+YsMxiIK8HlGWG
hy3rDClSRlG7vtD/KIh2M2sxkqb7Hk2ed1u76yY/bJRtpxUp02V/U2dI80gp
2+rpjJ+iS9/ZHJ6vVskZ1AzVOsJSbw0vvwWmnCTpdIV1mJPKqHnvG8WoTuSi
GUFmSg7dm4kdXluYtOy2M6XW3kJUv1IuG9HQX7sjByzK2TRJIdjtMDltYx4b
wJxmj/vSuXKLXGsYW8oq5i08hQYEtqslFTyUH6+KDtPUuI8MqMdNEfNUOo9f
USjewaXy0G9ghmy7+AzIzHduHIQ2zIXKv2jeBePsUe9/RC8XwD5WrZl5PTEv
ioG+oZfufLgKzaCN3NdHo8EJ39DxdM25HdTfaA/VNE8rbxV4yTbFAR11bmHx
HYkL/+wylFoaHQ0DIEk1wGgQqpYUUEq+6tA7WkizZiV+ZgASGbZbh8bKb+Zn
GDbLFuLSrSWYy/MwhFXSHOv+SIIaAEd7tr8gfJE5PQgusVuzfNdxxsLKNDX2
4yMnrDZUttbSYT92E/+QNufBkFn6vRDPfkhsxI2TFfxFwqBclcmj5QGtwAG5
dJ0kxE/8ywQyhqw5byLU0GQZ95C3NSHeJYiRhYH5V7PYXvBwJKiNkcl2M2cr
LPA9jSwyOUlS0fRSbmYg+uCHXGzEzwVIOF1M58745Q3f29/N8zrGz+V7JFhq
H3j2UGXfFtoSoeixWFTBQUd46XC9BJcBrHOLVXkiyfrbyLWt5l8CiB0xy8iJ
ML7Eoyh9MbVXG/yEV/Ck4xvTf3DT3qWtrCf2Tl4OJv/9o2739iWXk/SFKzI5
XtTHxuagy83aZBMQBZeQIo8MLxVL8QdxDhWoMjcc17HHNpJ3YMUe52zhNT8l
vhiNRckguyAFCa0Wcot/gAPmnCyY8MZwns0K5VlUuMHREbl9+DNR7QEqwFvm
8gML6JwnQPDIwLNa3qRKSr2lAL3XkD3P1ubGx23ubYzv3YNR3Xyd6oWxndrh
Xzb7K8i/AWObk0BOK/3ovAZkrZsBJ+26LOtM0pkEccp1Ff0YPS44iwbwV0B2
gYHNSYq8JJe8gKNB2uyHbNj8inia+mV5r7McShBQobbIcRfrImHQTv9bimwN
RKNhO2BNlSUgroKGcFdjO4SN3M19cn9ckwKLZiAKpJpBICoNJj/9v1nMigSu
L/6uZfdo3qLCMzvDdWRT2J+qAxvRLU8BWSuUNaTLeGzgQVWh6mC77RcQ/n5O
A918VatmU3QJRKbHEyoz9Uqa3lDNCntbUEb3NiFcRqQhFCo+ESWe+DS+8Cwy
+F2HfzJGn1w2qVQgP4QjaAjrNfDndhR3gpMva+lmn+6Ip5DdIc6PPSALTJib
9hORDVFAzUFTY21r/Ovv7UhJo7KsZIrHeF3L1uGlcIyAnMCBSGCm9FlgfSDt
Uha3VPIQfzlVh8TDjhhGJC8uNk52hh/kCbkGkm5jXKmS6+MWDvPkSoHMPVk7
QeaVEFpngeErhYOnrPxhuVwRyfEL8cfX8VDAwdCeFhoiDc0Gowgn8X6l0iIu
eUVlCaG0YOESKnTUzB5iA9HmRh0Yk7S4sGAixRuI6kzNLpNtbZz55UDB6k5z
t3uWtx4YFFyh8/QTdRJ0CBSmuF2pxOJUDKibbBnTziqnAeD2A2utiJzDaYMH
xbhnIyYg/HiwY5m/qcHcqZkMz90xqKbHcE7zi+SX1fwVZJc4dx4d8br/CY4f
3H3Xn+QRYxSXO3HtfcktwTA/t29S7Hbc9QOTPx5wbOpyip6+wYz0XN8ZoQMi
DkMZWQu239JZUIPgt6XphzhoeHbCY4BNOxRJA8aBrQOgxZxeYTb32uofjkt8
YoM7+KvS9qL5Ee7ABDtRl+6TwUTnVQYIFtnmA6/V2ZzoSPebnSR9AYlWUHJB
GT8wtXl6sD+ibB+C+qRIo0e2PZiaQsvFqtMlgiT1GW/tcaGRfTZkWxCNxXPL
fpcpJWssDZduXoBpQWjNmXKP0JwnJ8sEiHSDzAEZpViBdo3B5p/cdpdGC3mg
lwXLDggx36vB2WXiufBhyx7dhV5fdiE+V9FkoZNjUKTKZDsRda9Cr3izpDAX
vzQecHwDBC/bM34n/MMZRF+a8lXmULdrep2Uvj69Yv5Bf1rkqAx3UNIlX3qX
BYYzU2HzkuCeohlAz4OPVXTK0CF7Wky54CXuh35lrP9bRclfLqZD/ygsNJCr
QNWBWh99vEz7sWdpbyMqMIIrf6hADP94gFoWv4YHr9TtEBeragCq4pYUC2rN
CIMNd+sS+0reRepLJ0sV2ZahNN2wIsvLqhFgQ66NMrLDpizX4ePYUgQ43AL4
kcvx/VNgyzhvBXpMHAvdE27tupJmfZtUxR2qN6PB8pAV74NzEDfzPJqid3ph
zTGh7HuKHk7QM5WKSD6vRQd7BTgxnfoFdzU9ON/iMfn7r7cJe9umQuCSh8UU
2xKfzz3VsH17/cLuBIHTtZT6Cy+O5/e8m0jd3bTi+GXqQQDlkkh5uSQxpo05
hbxq/grjtyTvank1dTot60M+DQntdd2fBSaSp7wgbrj5xWvvGDKotvWkLr4j
nDsuiqTYKdZ5i+lugO1ObUQQiH75fvlrPJRA6he9f9Yn4Hp5k0DBqSfiVunQ
qxROEHAhJaQmtDfI5gVyUO6pL/FwyHfVgDt/fTw4d0ffRMuQd79sh+x8y1s7
bP7ptGh6EXZ/vXCftXqkCPAsuX9XaFQ7diulK8+QRH29ih5ENjW1xMOmVXVF
1zHqsSPofkrqSYCUTdLGvo4yJQiG5WsCLJ4UIDz0BGkoT8COZVEcz3irQVfF
26XsOqswY26NUJ5JQmdJZ3OBYBEZl4cOOi/UrJ5sdGvKmRidTJ7qeYiWGTy8
7QPWI0sxx6IqR+RXswySf2pV75kDWEUAsukbYM/x+ZoVX0dhUwlrvXKUIUL+
LiWOa8ItLMsxotsYcxPxE5JTp4RyXBq69nNUBvfmC6FLdIi0I3QBsbBGh7qu
4c1xuiEn7LgCIBXIgdw3Z68C9zJVYTHnJuj97pPnlEexOXdbY28TT+Jt214I
cw4KJNe0jvx3y91OcxTqijO/RmJA++k4WLyCJb0m9ITW6q9rnb7ACUilHgYo
gi3MgQ6Trn4WavL1SRty5U2WjCruuGP11GSJ/Aedcng7KjGdrPIYwGKmt7GA
eEX6SkgA0832+p3/7bOrz+KXPOoaQJ6/GIj1xcix7RRYH8ZXOtb4Qlh0vHXr
qSRr59B6zYKttwq5AnUcMsrrjTnjmd6HpqSj2JHXWDhrkA6A0QwKkmtEbSO6
e16ZvPDmqnQehu8l1Da7LlNdIaC0+yCoDtfrNsh+3NaVxMHJAUgIiV7sp47n
/RKt7ZcRJitj1PpN+nTU93wBC5DHfIxbr0AOT4R2hM2MU8cTt1sgWXorBoGf
rdNyGcnbQ1OHNf8G68ThbrHJIhP7EG7fvxJUs3OeUUTGHHYrB15dYbZ9lUDq
8tDhgDgrUeCz6nmtr8UMwcdfLtGhhElavEjcC8VfE5cCVIeqOJXB3rfns/8D
ZGZFW7mSPgHm80FDQroYvXSlF8XE36IhCT6IWq7lfpJ089+Slv+BOU4ZLWLS
Ng1YewALK0wHgKGvfNeW2tFFz73y7mHx3m4XrmMICkaQeLP9d6KwpAZ0xN3Q
lMbn6kgTfSoHsQX1SAiEXXUkaoXvxRgRV18qiiANcAr8ziCzcnF/kbdho10i
eGRjxBz/F2oD4JMPKUaURqX2BKICl9MEkyliDLnuAhcrWXZBIWgSAhq1oPot
YXX0qCx3U8OUY9GvVh0xjW3OXiHIrJ0KWq/IaNkk8u74c/aZPdl38souFRum
O7qd9svH5jy9SMyc4SNlup/62Jg2W70k8xG1GI4iWSDAWVWvckQiWBxG7nS/
Ofwxnj6taIxtKZOX0kHVRkxdSkRrB4ftpQHC43kai1FBCISzrzOdEbc+EodJ
iC1SPwT5/0T2H+xV0Z+FQR5K0eUZ5VK4M7i8q6ITJwOtqHLiB4azoNOe2KeB
4FvOtl7rZAS2+xwxtaAtjQKXtRDgHeF8eKA86yGNAiUA1saJ5mA7mfRjTiG1
3m1wmX/SvBz6qg1XjMoBG7a2hmdqgEE/wdn+Q2gP7mLEXo9H6kco/+3amrgn
qlzJ7c9ByNaRdJQ99iYoZSq845W13hFqbxDNByRG2GOBoqOr1MLZfcwkUeu9
LMwbWa2kzh6+oSVmjpFc69By0dv4bO29nrQu+OxOSA4e1Bq7lfi7Zn8jkoRU
jRNMmzRD6UEa1iOqqxf2edHBRj8JFA5ovFNM4HwCedsykDesoFupt1je19Ys
AAfp9+r2BOMpIkw2dBHJAHvCHU+fJXeqLA27Er/1k7QoImmdZf0GdoTsgq3A
WrhC7VQHbO34Ze9NBwvuQgr0v1wY8ihG7DaZjmQVXnX83344fCVp1NOWyF+E
LJEyCUgTT16TBhp29/pb5p8UdG+JUmyjsTcFNTmo6fEA9S//A4Ch5H3YzJO7
XLF5r9v8GwKiNwHb+VHPDcJ7PtBj2OWcOE+y/XttE9uFjKaWDXf6L0vb/IBH
EJla/yOyYMTdgVn3ps73eAUxgPZNR42DXia8ELqZd/CVcqhp5KyIKcuwhsbn
Iy0sr4i3DMoi8ATQM4DJwNDtbj2F89iQOA1MHALGSdkCkEGmoDTNe0Pg2ve+
E4rgSJZKXPm6MCk1sltxYUy9Af9hB7fN3SYFuLXEIcPQ1p84T4tzjFsoyhdm
OksJ2Em61aXV/SU5sTPZ8Rh8AbGjPONRhjLAGl41ppBoKp5ru8obfRy/X4oH
TcayewbRC9tDKYyyiCNjGLuahkt8nPJwp1j0whTA3mzy94X+Cg13xMpcBSVM
ta4AvhG4Zc6CGQQ+iSAp/kQGF4OiHXHsoJfVQXb/ui9972m1stsBIdDaYiXn
rvUowwIMhM0FyJc4tJohfjX1mqoXCr4FSzsg0qF4OqrnWQbxcfFQwpumICEE
4T5TQ82SoK5x0pTWoh3hD5zHSlclU5n+1l+iuPQ9HbAgeQh1q5gOD+SYnXET
3evT6SzgzLKcSMKGrOSToMysswIgCoY8p/hvNxz814wtSWICDqA/VYUvnmOJ
po6etYHvRxZkOa59UCZY66Fr0mdf2A1NGqwqoKO6A4Nuwpena0XzgWyC1sSW
dV6cpLm7eIAa7uuBGlXAoq1Gbaomivbk4coyZAWAeqNKRMuxFi1DxvN1eEs8
x6eQ+ayueLhq7lI1tG69VvMSPFy+HmqXX/r1hKsxCCxELuNAmq9k4XqGprht
R0bzJGKXggUtBzaP3cez6J7NrfuX0c7Py/wzBxrQEMvnMJ9/ReUHQgZNZ4yo
5QLnnOs6qG8KRrtVl4pw7jkBhFsSIk2lQfZspN37yzhtXFy9uVDnSn7cTfil
NHiV5HOMZQ4+tVgOLLqDSv7cD+4+Il7XGdCR7wp2FQyI/q/HUi6KRVhw6RuW
snWmoV8VtWzFxt6Z3VkyqfT4L0k62QQvlcpAM4pj4w2kqbEZelV02sw+wPnB
OKBXjhoRUHxkbU8Po6CCF7bhbkUJi4iRsNfgqYK68XaWEdiYcLRR7BxDgWJ4
/yyLXDJ0pMPD8jXy4swZeniCDuwWMERciDGtG+PtJJzLNSfyW85xs444Nd2D
cydHKyHOeKTbwiMZczTIqC78rTexLVPc37N5wnyVftMqZh2XGEXjZmk1LnQf
75TdNZ2Noeq465Me2pp6v4yZFwyGePcf1afm0WQ2BpKQUSYp4KjQ8nzesBvq
wDJVGdUng9bXp0X3luzW8Xo4wgkorIXpXHsCxzyuUEB5tPWVXPmxcy66BePq
F5rLlwS05jZ7l1/pn9A0dOV6P/miZ8blIiKUzdjl1B6qqzs6qUWirsvIkmzK
nPdxnVLypXFUoNylkA3SkBvoN31zeGvUwlXnS1Yqrp/8Mh7A1MPIoEKzwvXi
COYYnjQ9HQSa2+GxZsx3vdpS2erRPrxgywQHGOzcd7eT0dlcP5KWHSa34y5K
SM0o2Mm5X3GQneDAlCtvYFa8y+cidC3OmVD3L4Ms4a2xlSxDq66HRBGtqWeN
8jJaAW9xgcLCI5QeDM8ScQD+YRyp/uEOXyYJrQaPjM4c5OFfeE7YWSiQi+43
OEjqQ8NztTjfQYpq6vZ+Y1zN1ehFZtZgt5AxjOweRVz2fKveP82Lz0oJznMM
/G1g0QD37OY+/AW4XIjbKm9wIxXRvD6qIrKdJC+t9nU76TV7rExx1KyUB4s+
IDezxmsBmN5jdioVl8toNkQG9LdS5WqxdpORaUcgc/u1XFx1vpn3RAgXYZgS
2/8RvxUkEekOLfkdya1Lf9DJ2vQ7sWCYlJgqZ4qImVe01G2LXQza49XsBaFN
oNtxVi4PncdS0U+mUmy2Z4TV/RYe0S+NWBUlLQNvxs/aEuPAC74C98brKjy3
Bc3DTThAhpSywi/WD1gI2WAjhn+qfAdb6zRBcYIs8gesfgldbe4JHZzD/5yy
pNCnetxEN9AF/u9+z0h52aCP+3tJxv0Usw7AFgfBuxX1Kcr/yy2qKbqxzA44
Ebp4yoDxuNkUelFnhc1et6fAEO7O8/XtkEzNNMxTwXa6zOKo1E8BAijXNRi9
jVHduEIW+FRJDr1u9hIiG6k7ksCvD+GakxgBZ03zljs3bCjVyyJRUG+RnH/H
/oYiVtF4Fc/G9dePn8PzJ1QKRFHgYzz4WKK76NU2MNRtuTTK99F1f71EDJvQ
0HeLotcHW3ZfPjjf2dWVUgaNl573k7XrwwuA+ApfDK8ZwAVF+fwPGxcSl/oc
5FopbWcM9OCBIs4KVS6J69Judqv3cDxsKHrm3uqHEEydWJ2y6s1pepKLzob4
qrgjx91nxuPbjLOI62DkP1lorgYA0gigtWJCjdhu7MRn7MIL1or3BeQnNxzX
wrwIfm6rD4n4rd/npC3qCGgvpU6yaZYj8J1NWzmUF+P+28lnO269XXh18TuY
yOCuKwDBVVwTKhpu+DFJeSGN3smDiyF7bgYktWNpRDIZrm4r0bweScxpj4YB
iDctdugYlP6fTZE29nfdYK3gPtm30NXtPMiS4786itPJjvTAQCQruDfHxvDr
WRUQ1Ob7QZqIa2zvdH2oav4227MKZ7aeIo2ct4EjpRBWptQ2rcUeHSusVRKD
9QS2Wz56WbB4DcznURjAjWnTSWDgKsy03v4nZK1EHkEQjFxJ2KwtFeuBWJLf
4valf4oZKt1mWhJdSLThaMSOgs5ylng86eTR2xR13MUi4xr97klEdg/AdXIs
XZFKr76Mmwr86dkKu5zZDzCyYSf94VgAfx5lpISeEpdmlq2jayrbwnXdUVAr
2UlrTo+TJwMTrHWs4NHbU5tvHiHgKZOU/+S9vBDoHQ3AVxCi0RHhOealDyIR
x2yxajD7TJiAePk3u7T2TLs6sxo3HJaTI2V5f33uX8sKH8+ljvQWx/voERdk
0O7qg3BKlj7m2zb+qnxXiwI4DrtcfDbN5WaSxAtZLd3Yj8Wc7xrZeCGg+Tqe
OFGQIuBWxg5BWO3+94JNiTyDMnIQVXD81TthoiRh7bFzBtfsbRyQEOElrHiQ
Mf1PEhJ3SZuJ1jLKk14gOJsatWfW5uGXoeRfVmjpyteEu2Hu29l93SQwQHp7
READbC3pbbQgy4lL9e7XH588pzo2yFTBLTZ/6O7/227pzl1aQD/28IIOhPfR
5f0Qvw1cbz89T+aIGDhkESIUU4kK8v9/IyvxnUyNbGT0zmcxrv8yucAu+OjT
tbMF9ihypUjnQRhD5Nb9M1+30WGqdY07/dP9oPtVUgzr4OpCHRLyg0HXsDL1
Jtxwvb6J3yvQDiAJgtUcjiqhHEsvdLWXZmQRlo0tcCHGvQHyObSwEZRLhwt4
3AjYezJcjGMXnx/k4fMQE1UeZXvWciV+X5lhXhegf9Ni1Zrbep6IWgi/lW9y
nHuyhBeDUK92lNjwjHWiuWKS4rhPBWq5X5YtYlaA/aeqB4X1Tvya2r71dU7a
sGGjMXkLzrXKHDmOO4wCMZrasbeFZfNqSj0WLAuJomQz8HJKho4ojoPD0043
KTrwg2SkDv5reKyp5NpNMTqI8ubp56sQVcbiqNVPrH8D4UPFlX9fPZ6k2kg/
rbdIDTftdcGjzpJky6LJ3Yxp9djgssd0Hci+x+2Bco5ks3n2Ad4S9NzH7EUV
0CtDbWv+SdELISuswgXbWBe3WCjJP0oZ0O6AmndCpzwAmBUfgeGC1kccOTiV
EWMvx+imv6TqRJSQNDbuj/EX7ciNC/qf4J5gHj/gMeUIWNM7vIRdBb1PyNFc
fPPKiCphBMF8XAxS0qB9JIl9PWU8bc6UVotR9k/mkEuOJJfJZTgFs8qZDA0P
AZwMHKsfYPBOabcmJFKIkEO+fdEqO1js9NuN30aOBkHGkQWOyoZD4EQ/u4Gu
DA1x+KqkmkmboJnnzkFSsELfBoyotwn2NUpx7WJWPvqCW1GzsEgvXUQphygG
9Sff1LSOarqk2SoxVMk2uGkFSb15lZ0J0JEIWyDGO3WKuEKPdkcDhpWYpf7W
/MzAdiDAnQx6yzNbQo80ejiztDwXSvk+9MSKb7Qa1b0m/3DlyRYNN9faA5ix
JZOz6VQ17aaxvyR4Q4CWw0ZyO3LtY30no5zXLN2cfNmvdeYTws7P4UPFcaux
Dz6jppBW+nBlne01hhamzyZ7g8lJ6GNE1E9DXVCYx6qj2RAF5/qUo04wzdW/
Z4Eyogc6D53t+Pv0HUViO9EWPlaY+wLH6WIrHM/+LL0Ip/7/sb2BBL4Z3WLY
UvnUgZFMMkW8tkPKRCl28JZxHLyvPb8rZs3AgU0Sqs1S1iy0jJ7FMrb3GXmH
IfJNa6HHLxJtI3F4ZMrGgT7Gix/rVP7+hx8sonx/Qy1LgSTSyr99hIvczzXd
DFGJKRQn3+K/GiV354EURw4bFNluTNzQ12xXmmZJRCE1NLevOMVVoX0Nm0VG
uwa0Z+aUs6u/IURaAgPBvRgfCVZx7uGqhRxuoSaz7KbVzrhY7HXBrfV9zwAX
78Z7tCEH8IC6NY5xs1dWI9aUL93YtErc7bdXCjdozg75NyCjfFE9sGteZImW
sOdS0ih5BDCSDfOe9NO8DDMJ2SauSLnKdGQwjSdmqSXH3dVlWH2DClkOF2ep
Oq9CZ5hPGZjM+54RWPgaKSyCS5/6MgU4rk2gy6ybks+fdzNLuenayPgNx8cU
IaWWofWJUyxi1CLVuq8O6ZmKuoJt02hzz3Rbx/PqkjFOgfAvl76iKpIqUMDT
4fhL9B2sh4lXavVXlR9ZdTwz5ZkGzZiDLWrg/+TQq9uHZk7rzewJNMhJu9qf
I60bk81et1KAIjiEokJWMSH9oG1Onih2pUQ9tNpmO9I/RceaUUunLqSZwsff
cY7gYGj4NOTfpirO7xmWJPU+1kSQvk7ALJrrINYueHSXGXVk+MdlHZjodxZj
sLavDyD14efqD4E4/4/lBq8EFzw8VjAVhJQfRCC73k39MhV6JcdVjh9SpZBA
1dxLxHWX372AChxbY61xONZ/nLo1lEa24QxKTFP8/L0p3droIAR2MzDNK++y
nj9viSHavGPaD7G2xgZlS1VTdfbVIRv9QuVld40PyGz6iHzSxtul0YjkBYjI
FQWEVIQ7hlTQaT1G2Dh4JPSue/+LWA8kP7NZLv+HFJGHqB1tIQb77094jLkw
BEBfM3egd4HjLeE+2j39JxMSxGxxgB5l22S45gRB9vGnAM9+rgL+xur3R6Ll
aTLwcCBJjG5Ws2yhpY8a5uxjQqVMZ/85jMmAjeu7YUp9pL8Q3PUNfAHiQ3HT
ddZemO+aQhz1c5fEC28ET4IteHevd6nalu9ivKBnppsmEyq0BK18msxf7C5W
yD2yU19oMY843vnrPuyCmRNQe6g7l46CdhPDl/EM4oO15Ql+Q2WnNqKprU81
uTnUH/PWCvuuOEFCUDyzzJx29yh/v2C5pDNu5/O8LLTzcCcwWpPozk1s22kQ
RcHwMtpNFvg8xXvJJDvvI6vdIdjd6EjVGPHeme0HqvTHpOFH791FhmlO8tpf
nLSqIbNIoRLc58DESRZNy73JwvPDlXQavbVc2V9hXCNu2yn2sTpTsTPBBgxy
UgYnsI9+C88G7C/pbxGwz5R7CD07RfTXl6kFs0sBYIYQE5soUXp0v5lttDG+
jAXY/3oNUugKvTxiVBx4/OzWFkNAPEYH2ByA6bvXhmitTNpOyqFZWSeX2Nys
ayxjKWhW2gtRAit9Jw6Rv6AECQYgOiaSYxX6hwQAkA+jzJYuWNDyu5nAOxmb
ufrq7pIdI58z1+bfyZkmASot5n9bIrHd4/Heo6Vs5RtgaLwcF2dwjytDFJ+P
ng4W6CcB9v8ZmsCpzznTDT074cPhc6NOrDwCT0RRV+qOUrEjzNXluQZIgcew
99Br0KJqkM/sZ0iHj5PGrQ6JBCqRG1WB0qL5hdDPtKXKxQXJvSFQ/JyURNPO
b6WxsF9fOqSuSXb+VDxc3SHcmqnQH0HQlvd4FfzNKK5XlEQJUpYS9DbT7VVy
4IZATyzposB+4Bxd9iT8T8zYNdkGC+/kX1+Bnxe6Q02uyQ1ek7jsfyAC8L6i
l9+US/L2sBPXfW9sPeYK36XuY5oqi92IhLu6H3DcspnXjM+Db3qIleMx0/6z
Ho1tyrm29Yon3q7NTpcOLCJQ6NDHj0HypTMcXPGFIIphAFIBM6As7Bg+G1dI
oxuXi+zHmg7YeHglyBpoGPKtTeSiLTvoAY5vAQbba/dpG4+jDJABbN0DYg3C
w4Q4WJg4HxCryuhPSiXRrgUzk1VIm4wygtwnlBRO6kodG2dduZ9DmD5ZrAPb
7BZG+T7Dczgr2RlYYZxnTpM8uu3PxdbNQkNKMRN7wPKcYN6/ixiiDMHgEKJc
H355RT9yQ7+C9lH0hzSmSx9Lo/hd7Mh3vUTMmwmocGG0U0pkmgB8vXbA3YRP
jWo/jarN9QsNoayeXnGZh8twTI6rJuCnNiLXxU0X4XgZmcWNHHiTbHaJDdd4
u3oV0zGqDncu0a0nZ/C8c+lIzhi4hua6kDDeFK/c/LV1myXHQaLqh7/+dqBJ
Eo9BDe0WyPFzBE2lRYHHlYEMeY4MPlrJ0nuHhFFpxN4X162W1Wvm8i4iY1I1
RpQ4QJFRh6ZX9vZYyIULjt8zAs18prDS9uweNxLxCRj3mxehc2aESpRwq4tA
6JofIRTrWXf3XLXvE0e19tZ8K+bwJOzuhwngqmfZry/JQJB14Og2AHNabFty
87qt3QAmSPngOfc11l96XkqUrxKqvNRtsmUNw+2yHNrsSwds3gCSUK/CZzQO
fs0+ZTvHypELRCjvjjN3eOd1q3JI802iz0JhP7WbayCwTv/VA7b4VP6xeZXn
v3TGXQJUS/4Qs7v9Lk2tfPsWvLtF7jb+S1lemtCtMpATqQ30n3AL3TXexm7h
Grm6MP2JzVZ3ZainO0kIGOZxpMxioEvu7SucZBcN4JqIEM4vsc7CyYaTE8At
GWyEZo1/3bF6orcN1IOMceXzX+OZiTjfUN5eeEf7qeYMwq3HtP4M5E8CfUkj
bjfY6tMCIgMj2C3Swi7KnbOcL1agNh0biWztS+7llNDGyU0g5Rsf//jIsdtG
2l+WjLUBSSIu8n3bZbErPHwYJaQmOHl+hgjWpuzLRQUhqxUxnPnjP4d1Y1YR
BiiHR71Z0fL9BnZZ/XWBS/vaHvK7L2NOuEekzlUL3PZNPDlRp6q7tzIuM62P
iBB7EOeK3I+WqCF0X+uNRpTu9QM8Z35FmbXshDjQS+1HZ1hI8S51PqnpNa9i
Mn6bzdwLWm0omxd5/dJfzYz4XniYsCUuKm7D7mgyliuQmqNsf7O56lLa5Jmz
HqPoBa665jffcULQprAggtXPzbyTrrGPLQmkx1gilLSkh/jkjEUK8jKIt3s6
1/ek8fvXQangX23ttkPTpui2CB28q4j1sW1Ti04AJpu35RouSpfpP40DsnKR
94KgjusejFH6Q9IQsnfEc+kvUMc7BFe5NVZcjwYFlWzwStWkwMjej5ns8Qi+
u2f47XNcDk2Gzr+8THmCiaUAFgq6BsBjyoP9Ue0m+E8JSDgO61QSlbW/Dc0r
f1g4jQtVAoXdvA8m2IXtjC4FtYLVZDDDeTEheQqsdGiHYIDgjiAIof/Z9KuH
GUoc/I7OroN4k/anJwozvNvGDdT0fhNlHeaHCVRvgLwRUwCE2WIdoE8w0qEF
+Q/HQmVGeMx5d65wikZLWaGUzY7+xiyltIc1XG5MO+dbB2qn0UbmkmV19KJu
HrrEwr/tfZaXyURSANqfREJ75E3avnD6D0WJgZeE0le0sY5LhUrzPASiosSM
psY1okdJUDDGoTpwo5q5xWfuftTCeaDyURsaP6/uNHjtAH/MdxFadBm/Qx56
EeEPvLXwCdm5PVMTz1irUN0KslIue9XZ2k6jV2M0nC479Fokxa8R8iirFgMH
Po1foGzXur979S4ght38+m/lAO1crxGUy5WQ5/f+XK4zlpplCKWkZwAOSxwi
vdGPbBYUMUAqc/sQ6cx2607bqzZEbpH12v3RPYP1MLrg8Lg8uBCoB/U/Pvqu
rBUpcrSiL2OwpVj5Bgc6UjAVVIz9xJBh7zmRSsna44ONZEt8+TdHbOo0lOGh
/6tFVNAqcIYn11/OHlBCAoezQMRXnx7WKDsye1hN+Ogz4i7LZIDYha1wWt0I
GskEC9vC97NhnLAt74wgL7iP2s41MgZtbM5tNv1if5XHE3qeWLhbDFdGJ6ZM
IZanozlWo7P26hvQkYD+ZS9s0SdIYjlew0wOpv1s5Nr1bguBm+QYpRtcI7/W
fx0U6aUm2jfm1J8gfAK39ePHtcTv+RWEtyshsoDI6Ce+B90p5kkj4kMRPqdA
kfa18QjPU5oc4TTJrlrjzdsEQSupEBBrJPZmAxQgeU927NInNLP4j5+54bVy
Gi+NpbOtB3tQsS98JQGKN4J/7bDc8parRyws18GnwVhXa1ZfjxN0y4I6VdEE
D5In/0YwWlS2hg/IQ4cZSdLmmvqVw8p/h9ZePh1TcfIGGg+ppAe3O6QV8Oqj
yW5x6zDdTtmCw26KySrp8lD+uZyzOa/jEGWJeGb5dQhcAvLI3A9DiQQ181w9
ER1LzXQX66cAsU2iZcHowFq7VwDWUrLoVz4dxEJIjHGn9VJDvkGzG40a2leX
s/qMghS4ig/FmcVKrH81r6B0hXmE+/LgH2U41+1D1DCmxMcWyuBkebUgn6Qg
j7/SwoJyzWAtSBSFwGtZAs6QW2b/C4JLN4z+a2BMTp8MNbNxhVCz1OLTz5pG
tcXSomnnkm16P3+0nWdX3biCQx9IwNuJ24iq5Z91UQx40KXYOvEdNmdRw85R
fqkrVwPByCzqMwvWsUZY6IyGzW6gdm5kiA6gzBOPy/sIiXmHrqeTFM89JPBY
UMWzceUR75UMimjb63xLNNGCnDW2zgD3zqMJN2K+LUbAkPtaqKA5FIQu0khP
Ij0vlmy9fVia4tMxGzS0jdRnC2RSz73UFMSpNqv6L5CDTKqR0T7+euSnrSSA
59K58c6AmSN28ONXBTGbxU3ULVrDb6hE6cIChwnFl6MAXqu8ue+kv+pUHt91
sbq8EYLmxVxSuAPYKTf3zeQQU6315K5rXwjivc3unTp+BXofH74Atjh9LW5a
j1ex7HhJdsPZe9AGF18M92cQ05Q8fdV6mp72FRFf7+G8OWF3szNil1x4GvQd
Yv6/ZCjP0jW3vUjm6ZY3PQJ3PLM5ZhymsE7BebZ/qGtCWXQ+VxOdBL0NOe53
Emzc0wcX9M+1Ct5vVf85r5yEdB+Q5eLfTpG2CkkNqq9mA1qe1MBT8NXkOiX1
Bu3zPHcfDxgQlbNN+DKlxm+kvsdDmxkpelwZZk7sDKcaNyExyuUTtayKHjlY
PRYzi0xF63zkfUcMME3C/c3JDa99o6dAGJQLTznm2N4WZdqtMPs8PbDa1mGL
CJbmbpjKw7oUxkydoigzqv5QGvr6ijzFPbLBOiJFojFpqXVpi2ocTLGfdadg
vPHuSOdedfROtYjKpKIXA62SgA064KcPJkRwnB6kcVVDJs9v/JlL4qAD8Ru3
Emiu44XvZbiOlCr/g2FRKpi5d4PDO9Rb68KkqroBwxG3gsok2ttAXTdrNqcO
3CNUCJC1gbSOgdZICIm3NGLoqzIvPGdgYqCm+43seIpVE1MD4OgpkZVcMBP6
XSgENT12m53OsD9LDa85/zBnoXlW802TH5Ef2d2YIZ9R1qktU7tI11G+ujmS
pxOO+cZiTB1OkeqU5tDKb/TpqoBldVAj4gOg2Sz1HnLbDjYVBU+UohVBO0/d
OEytWXM8ah7fWEbxeklJT/X4kYy9owNjOh7YVrlwKJ+DKBg2pievyGFWM3YE
LcrL+OsFlU5hVUiMOLk4prlmKvMEstsder/eMWXzdVyHnZZfwtVrWR4tGc3M
cINpKu38oCIglAsV+bszCPMSjbKZU/dP43jP5VT39+sYPJaaql2DXOGjEWMV
Zb9NBGLHta0GogUajDa3f5TW/X7eLdkFzoM6lad8DP53GxYeUFDc3cwJYcX3
gSu2dNRPlDv270RkIIFqFxjJkolkz327tgLHi8bV1OjsoJ26XGvaYcObxFtB
BV/uHFO2FG1O4DvCZNhnd9NTfbFU6L3XjxyUNjSH4qUbybeEmHpFGbPNwjPL
KHzVr1TbtmDnCbkjHn9Um3C734GJlSYrVU92ATkwCdLRa44CVJBXXNrGZ8mv
O+/7U2ULD7r3gTaVs+zxcmSxbGQZ9MkMpJvNrKN8HydSgtjWbjCcHSLHsBrg
WnvMeNoxhoh8KMDkQiIy2qXK7lGeY8eCzTY0BILuQc0DizZa1Fonz8gFzLK0
zBPsN2CGgXLC6I842OCCd/khODXLBraSAhaVhhbDhcDfWJ2KiW+2+RuY9sNa
gdA9ouTfL56rNE1z+iQq5ZT6H9Trj5lqWCmKV05rWcwXr3xvJ5Di4losFOkg
Ixo0CrJnaKniqTGpt7Z8Nhzi2snOK5vRxup9ft3lhOdF4orVbE95JozworkL
5DLTc0zvzIxYbg4FjQ5OzPYL1b2Syc9thCa+C1jNzit+umnUnYFw3mpTST6f
HTm325BnpRB/zHVYQfoRskEt9rZ5muzxTj6VfyFjOE6XIT+50dDES3zucM+s
p+PQFjOl8jK/qUHKTt96CsQNYcDzvopufd8iGyzDKwQHNeaLn4TZrj+Y3eMr
eEB7fe1O08nQnqq8h6JsBh4vE6E0JbXLNleKxCBEeHto1VLTgEj0nZknwkWd
JoX/wycRD7sYzfLG1AwCyvtjqWCtuK2B6do5aPzPdIH5t/s9WZcEc6d1RSjC
R04CVapCN3wlgyo5R9EYvKt9lWo52KJnAIOznwaCy9zW6EkYI2Jl9UDYmUgY
vXMaX21gODsV9rtObSHCn8P5NyLCMR8+UB8avWOGeDgXC3xp4RA7XRMO/xQW
cfTSm+yHMy1OncylyM/Vh73VfAfqQNfifzW8FAyB5ppWODVT+1dEvC2OzidI
zlbz6VfgGumFogy8Fbh2gpV1qbLzEgtoXwxblqdMO2dJ08DE8I/eSkpWcGNE
XE1eN8lxZTfKAKG80muJO5y4BtqPFCroIMIKcg3IQryYqCC8bPXh+3aP/05M
WW2ViGb+rvI2A4ydWoQYh976V9VNsLACBVEYxZObV5o/A+U/0gaNFOIOSisX
iW5YJN/vNqQLro2NEai2h3UzrAkvDQflQRSPdQKhCG89umeCSU4Eg3X3q7Th
G5gxLfNg4Jdkb+13p/+9LEgUEeg/kPYNHtdnHOjvoB7QTH/oB8QKqldaCXBm
m48Er1KOfd6VAWqh9C9qoliu4PKDHpXQy8ju3xjrS6uXVvhe12gl0ZWMYq4x
+U11qUn/xyscTKYmUg5ffP+ozOsvZuW28j7UoNsB1HjB/7z+skXDtcrDRinS
CWjIhcv+Ny0V+4iG4mmF0ILMXSr4K42/LJkRFNwdZdHpeIldcBMqrdwp4gXM
kiJ7gaEOobh19A5ysLHUcnyPEupQr227hNaIPJDwtgySu+s7UwyhwSNg+jAH
jRpiG8F8I48/v5ynmqclwf8jr+TcEMGuod1ZwtVU95hfLdgWBf0vAXhTKtbc
6wbmHdJd2iG25CdrKnZ7DxkcMIsxhOx7/AjWSbVCrmJRHvTtp5xKaB9cneNQ
dANsbkECVIZhQmoroE91DO170EwZDdl9hov6UD8zVEwWZXBBl43V65fgdyox
NhBGv16/uYGoKi9p+GfcNc+ZdG3GKSmX/Z3Mg7rzXMUTx2xUkI0gyHiWEBKy
KZU4gL6BKF9+UB+2AvVef8Brz0+LRLQ5gBwfxsWpUdVgHfduTiZ2kJsgvXAz
+MaQXRYoPP3V3C7yStBfuXf8HMNDKJqmR7c/UuKvjd/5rpbkADCBL7N8o9wA
36sC2wPMo8IX7Dky3mB4rMeSZPhTeAGA3V/0S1ejafV1F3II7H/9ywkuN3vo
jyKPE49wEfqRaT/LYI1aQDLZWCDiLTvLQUAbPlrDWSv4Cew5pGnzoCv7heVu
F8gm9HFwvS8WlNb8wTHSQPIkuSq6u0+gw58KA5cRok7nOLvO4iP2nYKmpuql
BWzUO6p/VO63wWJZwP3+iF+6DjIQVKx8pEKT/yhcaOL7MLFCwaMO9uhPEzXH
jlIaE+61MPMJzNyq55xV/JF2o2zPlAAQ7jOalrjRSspxRDIQ7ZymX4rquF2A
KtEezkaoSswUyaC9KMxIc4UgQdn4QayFVL5IG0wp9+MN6jTxQCSne8/J9JGI
eUQJbqerN04cvS0AgUp7TihVJO9pVC4jbVf3lyAX4b8iZFzDyTFNJFiyj/uf
qxJDIbZD0jX2X8I2YUagXiL7takokC6HV+Nb0nO9w2DbAafidvsEz/XKfU8t
g1OD3pBHs4stZapDukaiT/S4XYChH25y/6cUg6sK7sUo8EAvDUGzyA6IjKSU
FcfUaOyAwiuzLOUMKHQh0IWqnqFhWFtCqg/b6lKw3GOhKJOr1KQicDkZf63T
XzZI+4teqRlPz8AburzaEBgg0PE0/OnDvcsnPNt2tSeWWq+nWf4dbK6fqtoj
rNckuEJAYsA3scXdlVjKfod1JXyJnNqmPyJ9cgbXwFi3D1ln2M74DJI/CPKK
RXyGZnHoapgKXUipw224NJ33fO5d9TwK7MA2V3fdf2euUzOES5Mh/RIK5Dkb
XlHJxgy0FlnCM0ROrb+VIb8oZh0XClqiAOqS9SZaC+O3PgqmKtlLxOf77SHS
avLyAyjaDTSdSXyVW/JckdOcMDVicaObRwzityK/feFLFW3USeSDT+uIGLyn
verJx4BX1HLLihopk+y4UheDkxCHZBuUjfnyhdWiGpMrB34GX3/OOd2vIpSB
TgS2GIBZXyzkUdZqUB6CBzU+hd7N8wOpO4fG/FGOCB7AMWzYlC5zuURHhX6t
gNxL4vi1+xJQPbuwlXCwC1WX5CGW3GMkTGSwCU9PFhSAVyY6Ju6xmM2t7n6I
Ok6OqlAj79yNEEUjEpEDfxWBJmqBMhmMjzTxz/XcUCQqMy+r9ZSwyzM9u89O
OJXXu18N8u5dBM8Fkniq7HiylvmHxQCPLEZ8rqIXlJtV3fkNRRQkvaXH90QT
DCK1fFwU5aQuJRIvp32kaLrVx86gZVThjrZW8W9Q2vB1629+U1xuGw0f/QfS
0Hx3EaD24nANbbN4ffXWbnS6KiZcx8V0s6h1khAK79IZbk8CRXIeI3S2UA1b
jzjPOnXrbGFOkPEgXDbBoZKNiDwNZ5RIgAyRfrYNsgrEpkfR0DRmRtt6Hbgh
S6jubqHee1+hW4Dpa8eQnRNZPKzggW5fPcqKXhQgCAXf5JkO6QI1Xp/NBndn
7AqC96IoYAnHTR3M7Lm91WpEUj8aeCEuzKcO5zW/ozjgxnSWG3sbQFihKW8J
yhvTOCnmr8+GmPG2aB++1sU4aSPowtJu+6vKhCw/He3F9/+vKAGH1FbmDha4
9DbnZJ0fzEOTaGIubUSgxNy+Pl5WeWbZlpBMpphHwv82J7YCXzTk2dtNN/PR
33yJI0p93fofrjTluauQ1nIHUWpKpwV2KZ2Q+/Xzd3e4AtBnrdTDNws9iLL7
h20ssJYT6j2leSbxBPQF4yfhA1MY4fDyYo1z7OetCdMBIteO28dblL8lPNOL
zL+oV9/sWxUT/rs99T6WfRm6ev9aKaAefXQyUJvY8RD3oZ7/rA1YiwrAajYA
RdOoNyMvpInW3WUvuzAhLRq79KhMSSHng/nFyLcWHsaGkHNPXjie0pUCff/5
CnUjpP8jSukffG2KZftBE2tgG8IPXbxXwdw57kwU1DM0CrEeBQ5TUnJici84
UEH6/KC2CixKAMeIaoQluq2VCE4krbpy3gYTVFBDDOw+fwCf+HpDVXouaWG5
l/HlLact2w4MpRdhOx0BIz0wu8J5FpAi95sl3X/t9XIO80RR+i+bx7V7lNVv
T+HJz7KmRl1hrsDavThys+gmmu55VQA+rDLHLUmAAmgrvZaFm6eFQ56COOPo
CReZJ+IEa0JldCFFi4nR09UqiRJLFujEqGrg+cG8kVrxNaF3pfXALhByugmY
oibGkVZ/+MfRdLimDk6ufVO7evHAEbntGP8Qldmyd+Kyerd7VOlgT2jMf50J
/MAx1Xr7PsJqrUTJP8f0H/xE9jaoMqxg7vLJ3fxbKv4x+3IYVEkb7WW2Kv9P
ROrbMzFQ0FMz1tXbqF5sCkLugNmN+BehaAQb/a3H9m2bQhAHmCPF8Sm4oU3w
U5sRBeYHUAQGrI8S7eegggIanlzNrmTxJXKP4NWJ0pi8F0KmHk+05VBckblk
8rF35Au7Jm8J+aTeGKWrNtVfFHAfF2fmtiuhC0VIii5/M1ScgyOUVcWVwzhZ
3rmFJ3y/jg6qj5n46xZNJG6wWUV9psps4MMC0xGh9lI0fAFjIsDB3XsWaHJ3
IuJ4Z1cIdf9AoZgf/yxvUqS8TBFQfSjDWanreUEgP+l+FjnIqCOPJmVppr/L
GfRVK0l1AUPvyXwOfcB0QsAJ/5CSYnhz1Hk8yRaps7QOps7Im2Zw3al3uZf6
56L2P+eTz024atj2wrmZhAG+C4PT2ul4qV2YNRDOMXyt2drMTETJVAl7bGqQ
3WSMnaMwdVWOlik6UElDhY5LToJkpBy6iPRWchSnZzmh+TnfOX2zjAtpvf1r
Wv5pv80k03ml0lH03XkDdiCoyFkT6pHIQA2yIClwGUbH7xb4+V9myTWa0wHa
I3hydZx17kiCYDl6p9nfdAGvmspDeG6t1E4l8dsWBjWhDOopb7DZ6mHpHUSu
sFXNjhTP2ratSOlAONQIUWvTBYy2nkjVQ2jJjCYqZ/6Ruyj9zz2kgCDdUXsQ
wGQ3nZe41zwkvkHsy/39ZzJo6dhWUdCRLiswmp0A0O058W0SPQAaTr5EA7n7
5M1iLGCYKoCuXzeYxJeGjZmnGeLQwSxf6XeK3u8qwInLjwtOMs86NnuqXs5j
8veeDjKrRPxlmwdXM8rK9KvJOJ6HkiSp9aKrADV591u6sJ9D5UXHtc5zSnkr
qEZ0nmnK0wtLRziJ1G550ueQEFYPnJMsPT/r08HhQ2vNC2Cu+O1clKF51Ccp
kDdKH6x1srLpP5HxnWDfIVNffkAzkRhbRhEkMPlQ1tL1hcD1hlFBtC+Ox4h7
cprISvu9ek8X4cRoiSuNAMMoCeJCe3/EhMuMcAZ/jy60quqMmL6cty27I81X
SwW5htZjXB4wqTKOs2iBF3SVQ3RMj9gc5wmCXJxdr/vQpWygMklE0mqnclUo
6UtKXOF3sEA4nNRcR7WY4aPsvb/SDHlRFBnJH6mvqylXMiEj2xhwEw0H+hac
ml/yaNr+52D8M8Pp6sROScjy0q56JcuWE4L/njRfKg4Y8cWt6Ejl6/8YBjvj
YH+2xdk+NRMbk+YFbZRkZ4L/x0X8W2GdLmRf6+4LwW7ULXGVtQTpK9PTQ13M
+6CJjg0FQO2UISyBxn40imLra8pcSwSSzPPVqilCK8G30SnX3KOPksH/F4TY
C+P/7X17eIx3gwqzVBqNOB39yAljVUJIKUUb/91U/4F4hJvLYuLVdLTIVg92
ZKpOvFZB6rn9CnqHbtFQd9ubE54p6++QJmnHMarznbhZL6E5X0veWfmtMJ8+
b1kjkrPkK9PK17nsyCmEcCoIQ84nvd2/pXqIf0J/X+C79KXNEtcwhMndvaDL
om0gSPJpLUDKY5dt5HVXu6oK010nwj9Qkvce13bkDw8H0OTq4hXla7E4eQ0a
uf6tF5vRYNhDDrUMqZ03IK3bA02egp0iLbqFVxDTAbObgMJY7hC+DISmQUM4
3T3nAG3BH9WyezbQ7E8vPElFmNusWtPghYEee9d1600Nkj1LoI1vXGA11qcN
W/c+EmH2ixNG/CYK9oKe+1amRKBY/lewgelr8ffgN5BlawfX2lo/PfBj2lPE
eHP7EuIIJWAe4ejG/Nt0WYgSvYWJlTu9UWPSuZSXeuUC5s1gPBKEk9RhpVbf
qHivdyxjva+c30HCoZwFP4yPAJ6St9FPheOa3G89gRnYc/FX64vwyTbcydvr
OEJL5/7KUAH0avKpBb34GCLy+GVPg/27BCM5oaq0+UFn87h/doKMt7BGIG5b
nLA5CWvZlImlf6oSUGOZXOwW06fhC/xDOCsebUvW1v7eS1ZaVSca9SocTa5W
s4e/2p74NoKs/uloqmf38VRzWNXlzsze5IUrFDugQ6JksZMCqzZwjnHOh53N
z3rh/wEoInl1/cxhP52fkU3oHXHs7KzOpp0WST6bCxy6lSWD0wG7tM1qfu5M
zX3It0alqKb/mOc/oaX7FRgjgxcT2vdnL8kbNLaOi+QpHs/LyyJuS0yMuDfh
Dpmhn33hwExtduMiZIAHb7gJ1xn4oE+z7mv/SIHMqGYF4rl7UGUrwOlhYmZt
jQmvGt7FiJfz7daehXPT/3aobMLqdmuPYAN1Rei4LGLeXaMWsrkAGuRkPHJA
ZygJ1D38oqzNP77mm87Ri96HG2T9jv7Bq5lxX4EKhdO2eaYAB4H8WPZcwAn0
1mnShA2GfV54mQ2FnRsP7V0zggqyIsNz45HSdFGfW1lmrX94uufkBU47qAP5
JAWiI3zQuCJHVtQ0gy79zBwFqViGPk0GaPO1g7eALhUTlaRDs252XNFAXu0R
fN5MTp6I2Gb708fPfIlKnZnLJlGHYV/l/mpvQfMi70g4WEMUT/nGfq68mqww
f5qq0jrwKTGyNuOF0huK1eqkBBWIDync+GXdjDdu+Wmfgw86XvTyuGdtSTBD
1QQBxK/5288q+Bw9wlLgyuB1CJmlNQ44B8pt9M0O/F4YFcQ3bB/gnRq6SK9M
oOmfjrdM6IdkwlF9OedCS+MgDB37gs3murpfmxVELzgUeAyy1fL0SJjLAklq
ndl3hDLZVw0cCooJvanr68RgtiS8tTZCjSvc7fd02849r39WhkqlypB6lUGf
QiI6NRlUgDC0hQkn2YIjoT9rRDMeaqhv+VdhaP6o6+W2WXLtwx7diMADwd/H
BbXvzC8JRgNvcxvyD1HNBHba0XCrFzA0/DBsg/wfsld1p0IY5XIF3w6l7DFI
Us1tyg5u2ac+RbZ2cWtW+PEbDUzLbONk7DnyzIxjzYM/9rEhKV8US6yvVIIQ
9653IJ9S/5OUS1yGHgnoc1Lz8iJ0SJTqHiZ9KAxzCebLkNJybPomyKq7lfED
yL7xIru+HvEpyt9LxFPjAqxIluO3KFm8685CguWXsBe4wAXxAOhZmpw6ZYO1
QE78vrslrPVg3T1dVNVJveigs58l02H3dOQjpn3nZccsZYF6fU+Rbw+RTKpW
+brUxxKknj4LarXiCDPPRH49KoRhOFDCWiQsOBTGzymsXbrR1jSxgkCW6Eko
x7ls3ox2lMQ1z4n8joN6XuDsY+3wvMMmtsp6IVAvwRy7WQ3qOEETdeGXVw2k
VLUxd6tYXxGgEOBepQe3tEBXTwf9QvV6Izfm5yesMwh2JZlvlvuykq8FMq72
j2jXfZIAmCIrLnC8IJL5MwYFoieTNqNJwp7OCeaEZscmhIxxivUug6oqd9UE
TqaFttXCYOj1uRvKNZBl9GrO0ZGTl32UCGTLHdFZtKh4c1yXCdRVNsjTYguV
jg67FQt2sJ/LPIb2sL6pR8nIxjYXsYw/YFjZH1G+3/rROdT1adk+xDtRgWhj
/wrVGTry/A2O2j9867+i1YYCUXJ19IBdZg8yZJaH5L0R8R52fAjrOYdJ/ipa
dc/Pl9KDFkkqClU5z+6QXgbFIuqKeOB3a/s5HbSDQOrenUsN1IZg9hE0Z2Cv
G+WHztU+GgbxcTBA0I+kA6gYzUJ9EtgOypKs+gCLKDm4rUd2YRGyworOT8DI
sGz5TghmFPovH7v2xzFpeeO0J3/Uu1Gvft7ZdH91OUt9DeU4BN25bI0xRJDv
zXRg6EIolJVyV9Z9H69wG6ilx4y+oO0Uwtq1W9D71ketBGNJhuzFPqRSdIos
rhB0mRAe0xwuEFam3sgKFw7jh+rJxgisyKScADuzpwsuwyTtFUZ/iHzmvzfz
aCoN3Mp40VBOuv0S8nO2RvzuglIl3RgpJhM/CF9DSEELNgJJGu13euza54oz
JL0SSd5g1ivnHNnAlaik76af2RxpZeCx+u7PpaLwNn0QirP6Q4NQQUrHyw+j
LQxgejIJ3vXWNtbE2/OZd84WKTgR71kDua7rDb7ZTeO9gkvHexJ9GeyB1xPn
OCu8Ytr5cAw2V7zoJfNwN6ke7H4kkjcfio9SSNDxQN1IsfuQPFDWOJMIfHQw
OfRz083EU8BGVnqydqAeKJD5WpvTqyrnSDijVKAPIzgG9VachItuApfMXIzc
B4AxcoZRAWHw7qS9BhsiNCN5GwyvcK4hedmxftoH/1+KtfH1+hJ+gDMLKxzk
8ZxweZ8a3fwR5cYV6p2DFNxti0Jnuq4SrkEOpcIfqjU9jEIlC6/J0CMm1/h3
6O5WM/0vEFuRvjzvfiBTL5k523ouYp5eutQP4h7lw8wBmUGeA4Xi5OFh7cQi
pJkHDUWsn7QhE9ygWzIq6xh2JFJ3gstLdOSdmwYFOPdaKb7E7g4Giy6qhlhN
SKiF3GI5W2Je6EcHbIWgEjIXMqOPocbcmS2CGAyF7k6Bbue8/c3JqOKNFRU7
Hab222RhQ7VyAW8RTqybsKdw7r7DYuLnrQwMiDdwWX8dAK0Z9f4bFk17F6dV
dtGnw2uGQyUO6TmXc2D0vs8uA3cFUb0MGAO+k9sEGzlvNCjkpRXFOdZ1MTai
rnkk6uWeuMgiqd6z96H181nJ9mHu+UyaYpYHWKOno+6DBo6rICMrcyjs8enB
ZuTJ/A3PJfv5i4j3ExvUeLa1rDO6WqBzwD5aTwBVabB9eKmw0OkWcyT+XyTJ
9CRshalOoBi5zz6gJXeq/7TrlvQVRee5H//WcqynBtoC5ji44Gf8TaMm8F40
HVJ0uzxutr9DyIHNDPyq3apb2ML1tpsLJjfMS4fwpGrkYLlnD4H/kmE1PHla
ZV6zjrAegOk09fVpz2ZlI6ab4y6BEtbqB9NBf0O+qLVcBIErQcIuSVjtmDyn
dvlVBt1hVVQMPDy82JlmWQdG3QCMtoec+Bwsb8c1rjoXGrjWcZQcbVFemGV+
6yYnlJUkq9CURg64wPSg9mJ6CpkLBAABAGv9Jk6yPLjTkkjAV9mJyNkEIBAr
UTMIbFLfoPrSb+u0Hd46DJmzJ5C9gJqHfmJcTV620hHWfIFC/KiLBq+Kt7hY
4+lV4CLxPmBklRwxTHcMhYJV/aBPHN4BrYrQat/rDyP0fQG6myLfJrY6Zw2F
tB2MB/83AIKwfEs+fzY+dYYHo5bPkHLH5WOTjogzFm2woFNAvfEQV963sIVh
H9gAvsvu8eAQ1mdrx7tvrpSo7sl3lNcHRtdEnXG7xxUYQnZn/XfmovfCgwy8
mCNcFuiN/GdkbnxU/OV+32xm+PhpHADgG36oj5XH0qyxrjAAHc4ZseRMKDm8
IV99KAgUen59WMRnemjkvnguDh+bQCakw5o9tcnzZtYc/Y6gGofHdflbFr7m
ztX7nhR3qhkU4vTmnj6PpyjSUqQw1LLp+lM9pHoKJ2KPInSIjR5OadRagy9H
ZYX/yq1cP/c+SWmVAjLAou1tWY8CL9jl5/uZ7oS20ylZDEzV1EDkWRmHg8TV
xrh1vpNUpJW1nEjjwrYTJCX7XRxcqOMKq1HYHN/gxbnjhLIQf/8e6esidmX3
qT8Wbo0vCQndX9ymmgu+XSIGfwodfneUOs38Y9u3Ff9mZV3jQarlAtZb3kvh
oJYlXOtGktcA6+y0f/N8tbe5dFAfUAD9ClMGVaNqJG9Ekx8C7d/ycnJVVEia
p7Xpx8dciSKh7iUcyPOmVNmBA0efTq3sr3ZdXjSYGBiTFQ27T4/e3XLX2BVW
RzzBMhjc/FvrgbOQyzVwpVcyw16Nd6dEqpRw7RQR6s5f+rGiutjsciWSMeUL
+3bMpCmo1/15eFresdayGQMraVAO+qeX9MXj7YrPtSZ1Xn+AUa/DXcfwv86v
xZKrFkM5CMGVqOBAZkOVTFBV6V2n8xKzZGD9vCen0RP6UugPfdg2H50x3T3d
teKW4NFs+7YYAigwyiFX7TU0p5NXrKsIbvDgPkMnsWmBQZF8E+EgZFQm/n+V
oTRl60mf7/MoAicXMBYbhPnFi7o3DS44oQ7aiClKRuQgWeVbUrTvgWw5h8NY
7qXedimHE6n1znN2vJX5KXcXFoj1KwKNGQ9jFqml00HG9pEmGooOa15HQ85w
MBOav7/umoPqnmrn4LT8dM5OCfUe8bztaHJp06t7QEJDtTq+i8S9A01sxujc
d7cek9Mu8J+N1R4PhCUhiVQDsNC+fHAAaObbO+gJPUq769SOWbVhm8p0xcjH
N/L5yQOcvkCIi7O4bXBoS/W3zcGEzdF3VfpKEJJ8UXORZFD1iG1FTHVvy6TU
npBViO+ptGrXkgp/VfCbxb9m7lnzpsj+YCt4xQgiLqI2sCKO3jxC8VaZQiif
nRwhMsbOei6kX49RJ89ET+vyb1ql1Rb+SQFxELUMR5JqV02E3Dr6sx/v+mhU
ptNziiEPhFYstoTQBy5Vs7ygfDBUk+VEMlNPmPnSe/BatDBAkvsI+DLf9MSH
6ZK+kLvrKoU3uNnRBvpPZEsCbCdkQIg3ww+/1NhRPlu80wpi4W6DE6ubBOHn
04OsI8BPXmGIMyTq+PXkZN2Hki5PuV7/kMnOFYQoiFCHvUM1kPRpUyblGMta
VtPN2GXMYe9AM+i1F8XDg/Qyf+uLaENyHZCE1JTDp/APTe8z2+Xyx6xUXuvb
ARXPW7qHpI8estw93c3kMcUg3wEveNcYJYrLoBDkW1PNubpIZB7IHu0AoBz0
OLFt8FkZ2P2FNlL4wxxTo8L88X0OhUcDJ7fzI2+l4DCebaePIIT74DRauC8r
VTonaMJd2AqH6w9nMZke1EUUtBE0z1YIM6lOQq0ABPa789smNwxcINXkedH0
+HynOY1Lvq/xeqZ0kk/m1wuxgr/DH42OSaS8Jhs7SmKgFMkayRbMQUjsfsKW
XgK85TZNoDdvn6s6RISysmD80Xax/g4dsx1+4AINNACHvOEpfZHWix92zs8x
LUgNZYHL0eWuuLdSvz0Z7DkMLX6/BCR31KbZCEx8FbLFB10hDFr3i8v2OooJ
KvLbCNVxqVGXZN54ubr+hsAut2rlPGIjU910LQoM6DxaVxTuG263q9R4IZuc
v/Htvw+9zIYjzhOLG+gkGf/hdQKy38CGmYBmbuu8WMjjcqC1/eEKdFXvJ7I1
UMYXnvuIJzEmUjW2pNR0Zx5I7lVwT45XHz0YEwCTIFRjM90gUf8wcVeDpXY6
9ywx6EM/CGo21kVJOW7aw1XAPcwGAvmk6sTpxmp0rUg7JqrdYtFO/u82tvc1
DPlt5/GgQyyoFTMsHDVKKUEUoayZVVZmC5isb3EO1fN7jJk+/bY3oAUwzq/D
b9+I3tQ8pez5hA5oln7pRxw/U3uNwclAfkWgHTdoUtGYTtpKqudASTkeYkPA
P8W57OuQg1vSDzBIq3ZXgssme3E/PPcUc8oii5z9H2ydVFK1P/jlYOO077xV
N+VFASxDi5LJohxL299mFNMlWJJE5zjXZ/T9NuRPeNAjJ3x+b2BvF3XbQHop
mdn186EWgOcx7Py0lkbPKz8LhfgoIjDvBplioRKO+vO2tSAqn6bzvo73ftuS
5T4Y3NiMUT4b7xTk5olULquFp2bVW14E5UDBvfvD7srShMhHl+eBLd8shaBr
6BN93GxWjYui1a7RVJAzq6xQSDn2FyrBiLPHfJsa1gWlbzH/xFDEuxtpKS8g
5XOwH6CdIxfY520NWbgivpmXolluduBmNHiyVDAUCl6+YHg40Czihhwosg90
D7VeqMvKQcQILBNlpnMJo0owh60O1pjvRzAJk3011g0HYimpiI+arGHahARF
whvU2AklUQIV0bZ01oq5/5aArdQtZ6XHe5GkQ035WQTai1JLRz9V331CPcY4
5jaRnnfkrCUbQIIHmPUP4Ne5igfRgL3f55MPt/yCrCTO49U3K9IWAD3bS6St
4PbVvw6J6/d48WvS0SycfoPXvK+ba7sD0H+H7OkZnW+PjbRgztlgQRynUtJq
b59jFhnRreStg2nBVFadNgaURigkZ++NfC3paicjUAnRxkjOYxn/LsmhhuB8
asFXWx+IUVdrg/jQDeNWTFFJ9Z94DCavZMXuaXR/Fvx6OhxdElIrP/NLxWx6
TdQzjiZTf5dpdYpoZziMJJknejg4N6+awfIq99Vu8jpiIzxqe6SPThlVOK/l
aHr4KGT3JGT/R17bZF0meYIUBc989DPkwcQvnnhUiFlxYamYaN4xnbR+NEa6
N72juXsiONOJR56ZS5P2w11Y6y6UqF8LXMgJWK2XuQNLUgthk+HBscYlYXbv
aEDs4ZYF0VL3enpfm6LJ1xesrHlqpKT0/uHHHreBrgQwRoKYvdc31DZaA1YS
rA26y9r0i+U8XVbnIjMocQldF2QMsqqUak2aReUSxMiAnel+rXrILF2fUIcp
PsnRQOxA/UdNthnp65HVtHWDn6ir/WsndCSP02PgwXk206Ev78tETua+3itp
5rpwsPecxTTQJV7bET86vKU70zZOX8WI/skvkIiP5XVc5Qh9sA6HoMZS9HPA
0jcrfwEPqeZUb9IvcbSLpocGKAOd3R5tamJL0MbaBX6d5lAzTRSKdXtmWpCM
rs6nu3j3koRKIar3WdgTwMzqtXjl2UMsR8g6TtERwOfTdWXcJnaztnMTpiLh
+vXmTk5i4fbphSPWYHEO6rUJX30aBjhIxBa3/dLv6Smr4bNjZ2CEs0QBsoDu
utCZRgKhcQoJFh2OWIcHwb49Ra8dnpXb9gOEZ2aXS8QEsVQZ1sKWqCk/hjin
xlGan9Bm8rHEW4hambCFqykxpxysCOWCD1FM1xMGkOtpHQjddk8M+iJ/BFgv
uDC5ByuFeIS/rGeEglYHhjFsrmMitnhuSBUkVV2sQ8Sj8Gy5WUWMn7yfEEbh
8GGFnCcrf0ueOq7S7wSfCVFBHy1vE2Y8VelFid46gBGYub2QrKXUbmvJrRfi
Ft5JDBXbeBG+i6m9ehHfZbUweLw+UcuM9HHUsPTHPxSJCG5GaM3eM5nE2cub
pFkwGDwBGav3x1Fj2f9t8M7d0sqAr5LWUTk/DQWxqAtTCkeoElfijVH/r2jM
Qhdj/NXRmO/Kbvpo+/5SytAhc//GPiwYgQfX6QVhhYWEGjpOy0ofsw2F1Z5a
dPPg7w0kPW6KiHAXuEf1bctMshWlqtQQCTxKLz3sMOtZJ+c3Kai5mmZLSnBM
OChK7ykZ2wdyqXsQEExbXSJr3hzSC3xkR0DOhwuUpJd/EP7E2WSWLz7upgw/
dbnv8w2OkALyWI46CCkBYH/Or49KAIPEE2sEcVD2ZFe/7+jiDe5ivhrj3zLl
6TE2gohuvgxQTs5cjx0fGV65OB0o7ZzUBof41sZOMjiM0FEUyK6PD2VBCMUP
MGY7mRRzqP4/id3Gt8JRZaGewMmMD8aVKaTSaAA9Y+LwCJH3rUHCyImbynTN
2DlbBqBBIkz0ekBuLMrDzzrfKu61tYPCl57ghig7ZXQotAJJZ+quGs1EUOlq
LCrYeZ1a7RtsrqtNqlkJZnbn5HxhUxyiGwfGKrubsrLF81wWJlb6p7ov4QO2
53CBKw8d9YVacluLyUZHYDSj7HN1oZI3E8HCiBGmNTfMN9p8YMS2cg/2esPp
qjOuWu4Fnqg5r6YYMfSvuUJd8shOm0J2VHJJwVSNZSZ1V+UX/hlFc/x+sr9y
y3BfJOCrNpb+BV5Pr3yWWVUYdu2XlIhQzzQvM3OcSxtsm2UEX3oHXj0M5pfR
EOTitrFFG7vg50CzTaCvH0xKfx2A6pDyaW9bvyRgRtkukfQhLPe/VGcWux5X
O9ZhIhFj8iBkO1sL69oiMt9XrQZxxpRyR2Nks/pffXIi/bfK7gyfXwcyZXT3
LfZB9OkKJCNFE1wL7DL/geq/lPCmBBD5ZuD5w1/1qVXAfrdLMnSTGzR++1IW
oeaytVUG8ik9QORHEAsCYBhoC9UN4FIfffgY5hkIf0JviSif0pxmbUxLOZP8
LcwdUZ5fm2bnlO3dHeERYdBDyzdIWtDxDp1iYJYfoHxqKOxPdZGBhUQDQktN
tMjecDnpRT9YWI+5kB29bcZnHVjhDIqHvkZpYEsD7A03mU5SUG4qdB1+FOF3
i+tUlFwoEbrh1QE+Iwh/DXcl1N73KjWZdBxG2AFfUBzef71JC3DwzCrakpL3
B+AljgsnOlzltz/iJRCy1dzcsc2R4QKsU/8oe1EAKUWpRxDYN6lZ69tRPQHG
53ZMVVZ1EVv4jKvgp0kP6NcD2lPgvwPoZZBIgA0Bz3r++POwlKatcZyrKCPZ
plLI8HDpykSlFoTMb/4vZUp3MxDLrUzfK4vHyAEARQrBWzv8Njyza9M3kjA9
vKsyM2iI3vU8BNy0Qn8bWJrUiPjQRSd+i7KBlsl84nl27rOaAXwXzWLqp0kA
4Vev44FqAwC3+Kj5Nup4PaGAsZpDELKxhH42iDpIx3nWbM3xmok+ET69k30R
A07NV3f7F5kBWfkfN7Ty0t+zE1L+ckg8jb+ngrQElJA3gbuF1Al4CXPxE/kN
ZNSSb8wCKMypqo9O2FXHuQpUUn0Wzb8cI3l11TPwP4aSigE2sfPAMU3Na+uX
7h3OnS3YYHiyWaxrp5ld9ZZWQUsOeRnjEJu0ycsPQ46VW1DPT8R28grNA+1e
yHChuJh3BHabl0vbQCDtCHlb+e1L05PA6BB83sUAQuMJ53tIGeJegaIpzGo9
gcu1Th9hid++n7hcjVixu2jeMvIuU7ba9kZBhnewDaO16/mESZWoJ62avjvU
I1jggFzNkDQmrN02nnKDf+1yKI1sphokKe+orCsGhFQDP2Zs9Nji4srjktbm
X6gcl74AwPRxDTvAZfsUA6KarIVXnIR0pAFLR0DlGQwj35jtPMH2mZEKqitd
+FBKaqmAe5oUbxgW0f3K6WAcRqZ/K3QFar/tptxH/AlM87G3CaczzwFHebgr
cdF7BHCzIlPMllKp5prsIhrPzGUGXlVM2axXMOvvNbQKwfP6Ld3QC1hpwVS4
sfrm7lyZqXchxgHugzJZzQrarxyZgX5L/Xj3Bz8oIR2Ahz30rg0b8LsJMflD
xoDOXzNwH5SC91mS/47gLedGa31Y2cQgP9fD132KwTnF8Ip0E1mLMfuFnRYn
stmuDXdLGkdUBMyudBomRstafls8WajZ1gUCrjgwynV7KJHBcuahWPD78E66
RPZ0LGB7uNEdWWQCoxU/RyhTOjI6BJJJyYXpZiNikXLzLbckstR6ckPiH/lz
fVVmHdPLPtGC4jqQISemR2ZU/uHkVOyR1O1zeKSXO7M2flxfnxveopoFRCiQ
nTTqyHYPKp1EPNsz3tuMrB1eXb9N5w1du7ylE0sy4RhSHy/XjQZ7Rhul0OHg
/HI0L7383hLXev9p7KQzMA3eI0ykLdmAhgRa0HgUh/8O6HdUIn8FlO/slahZ
2pV4JFzv5XPR9IPK6bZvL09BbfXdLBPbQGwbe66mnpun3ADmeNUuAdW29Rqk
b/sGLfprl31wGV8u9GhzSs2oOjvrs8LnCJ2ooeAHoH/xWhRcJf65GmssjhJo
mq6zv+8Ctt6NSItGeZabfiKWQDnR4F69mNEYcj2gibcvBCF6E+PUNpRQ6SXF
mJ2hsDONiP9dBBMWcLspAvjapFfwcX3T1gg7s34qGEM2dga3QvEGMMtAw0zq
DzKzjN+Iifmp97Y65WgTaMixFdOzuC760ulq6W4YwdY+kdebi8s3vDycannH
y164hQtL849w1EK8uIQVBIaXaY/8wpd3/awzcT+/ntlsxEwWshF9I3YVsbMR
g6meiDohh0gh4HFyS4mjzmP0Fr8bsz+3kKuMsJ0NrrDNqPrKVBbKmp4SBS73
lqnyUeapOBRJE5AIi0V49197ln+N9Kd5tzIrdDTJ+2rfNM8tdqaHbp0MiOMN
ytoafLtPCwZ6g0LO6ojXgV3e22X5jk02VWJqVFNir0pMJh8sXtb4OjpM5SWA
p7K/InaAXoQv+RmkUPkFm9Mvrl52MsLuKF8QnlSl3L2aWRBEdEetzR+zqWQ+
LX+ZeZbMUADd/HP8PgpTf+7e8Riserj2NHFJC7o5gqLQdhZgx7pJgqh+ySFK
0WfvBvvmKE2vxA12sjQobLSLhLxywiF21M/YO4MSZTrllapp83Iyf72gYmXN
BfZFSiPKWEQRlcTNwnM3o3h97Jksa+BRkqpuJ97GsqpLrHS4yLopw+xuDqyK
FhBY+roT1u69XoTu00ER1Tmrd986CY0qnYXu9NBBHqhlUF36JVpaxymo1Pmv
3fVnKYdNQ+rYJ8fWtFBaaJR3MHbVMAV3CmiqbKGyqwpaZHzif+Zc2EXHKxbw
n5bYc257Cz9uRjR+0d4HeKRIjFYxorvkvXWrm2CZlXvOBcc46h5h0fNNWK9W
KBAysaO/Wf90n/8HMppj86i7edZxtoZdDZ//VXKe7I7EHTR7eSMbuwmYRM90
cqplo0YNVywDghQx1H6380AQV03ztfAA5PTP81ViT3/7dkQsOZXUZlnznGkn
PXcxwq+KxcpimdwhjSCflChyUfashXJGfgs2P9hct6UQe215qg9WwFEZN/qv
anRQRGDb6qzbrUTrbqTmuBaXuY8FKu10Qb0/QnoBQ583J9axOcASXumLryff
EPfNkC4ir04zViElU1qnTGSTnMxbxuzI4yQ522q8ZeBfulUs/sWy/n86Cxtm
8DpnecFFaaGClV5+qub6KjZdNBYUEExipQyQUiRLiFZ/QDu6B3YUMOfvOEYp
Y5z+xbO6hadxnEEfxr3OiNy6hkHANmtkncxhcFw78PHK7hS9LhPQe5ezoSHz
1Ij8j8gf952zG2Ob/X9UQMPb5/MOl7TfaQwdRNKtDStbYJwjijtKwPbsoS9l
2l8bNyE8YDC97w5qS2BBHeJmCpHTfr54Ri78Jmjh3VuYKmduZPTFSE+to+U3
TGDAaPR9fQxyUrBuQPN/kVrLtqHMYDkMli2DeuQlqaYFfYJh2YOAvTcYxgz2
aYH2nwO+UgW6RfdjFAHZBz4Qixq/vqYKohPylUcWKTow+flB5UHkOjexy3Fq
P9VI84/0PFh20GQKFydlPq2d5kYs9t4KHft2vjErAFxmezQxg/A3QancslAI
Q25aUhwPNUxbVpTjIGMI//9s5kRowxOEK7YaqWIYpEyIGPL9qJOClHkYek7P
c1PRmvj0WpbppAGHA3KFzatjAetidnetjuyMA9X5Hshfm0Vk7kLch5xtKK7w
gSyZY1PSpTggdEkxAv1S97fXuQN+3tfGqo8LstuXBkdizb+w+zfNozyKISwD
/6m3rH4/o+THkMrZXiTPTf877Ung6Qf24tunkFBe/q8NY2peFs3mzt6tRt80
T/7xdgYTQNB/h/ouCuJIN3DUyc1Xqr/Nmq3qYwzzvncoveGMUi3hIhPS9fs5
HHifl/incM4o5zF3nbVWRfEMygaJE8APtcGIyCh2sW6JKdL2cQz/j6Dkzthp
Cia+MAOvfQSeKLWQXMrpPxgKMzd/00LnanO48WN36v8aBd5KEwDJyJ3I+8Cj
R7OWCG7Nq7+dr1EcidsyHpAkaPFIp9zlhVWwJp5hfC2ml7eORw2xueiCqjMq
d4uF4bMo+m2aYd/voaa1d2Q9lS8PP7JjjCiyjRz2zNd7qkS15TuhS2OZiSy6
kDtnJfUNWiRfxTiNPr2cPbbuyqURu5KpEiIKvr7VDaSI82GfmDhU+AAOfV7u
MDCG1nmzpBkd0KfRpAcY5pf63czJlYe2ZQvCvGv8D45rhlflCXCclMop6Kx9
yQK55YJ/iHPXJi5SUfvHx6Q/chJFIl1Z1nwBloz+ByGOCeTZlQ0TvhCTDVdZ
0nPdGnRhQaLT6PH6CFxH3zpyXkrYDTP0dRGnnAaN2FvAT2CIVpMDi76LF9Yp
csO3nmMshYYw1KLFHVfF3G90P9yqpXd8XaA9TDyVd8F2QrQhHmu8L3dIKYYY
HeLrq27vDjW0elXehwXkLepEmUB+BIzc6/VcgPdypg7MnNfWsKAjnH4/BzPl
MukORaRgHOcM5Vvz2jR/tdfYo2bkrlkXrf526/8Y4WWVGZ15v1M44NqV5GrV
b8GLKGdly+xjDFdnIy2kFkNtXmOFzDx2BTDbuBt2NQukyOm2/0q2CHemsLu4
TBoBLuz6iZ93n+q5yMky4i6CJS9WPbwPlGDuRECACgRT3vdBGspoMTxEbF9v
ZwkHMa+THoktw3LQQ35jGEDYsBqclP/IRCGa8p7v7JRtYTGkk2vBOxyyXOPW
96hq0IVpNGeu0bORHwl3/DPI/q/btgRyyUGrTlBb16ETAqSeO3emyGvGBrDK
I1gz1WfiIgN+n0cx9yB79XP2sem+GjXXOXlzOhkSWLc9Lo/3P0YKEyj4casR
oCXimI9Vbn4qw2XTpcXSJocq/4zO8WHhRhuE1sjT8J8bsA7wkJv3VlVcc+Wy
3QreOhm6heTAiOSkPRJltggpttBRkVKnzUI0ZQRIV/t2RFoN9c+JOyrxuyLq
1H3Q6aysTDT4SlYLtFpF1+9Zt56oTWRis5XWrCdIo6lhe+CfA57/bHY8gyky
jfaFTjLYKg/YX5c8BYbK6UALxQXzKpMjbF5vJsVaO8mh8CVsndCWFFoN7Nwl
eZ0VvnDWqyRdM+ByodNggiLK2e+7Az6jdHX4D/z8AWd8/c4EfoGzd8/oTPiE
i04H/qgx823Gr2JLZfcZOXeIO46qXILffg0aM1EPnHz5b29wFNvBgrN6C/V8
Zy87WxJxLqXnnXyyAbZpc3vIfFMZdE71yejXlYsyK1cuJ9RzdXsZn2uo+U0P
7eKXHFF5vejF38Dv1FBOJXxHJgjXvxVdeI/UR6XBdCf44hznOHkfIX6Za8UV
H9rrY7lKc+87EYB/qTF7TNEesbU9wcqBAZu/ENOVJlzfhpBcFEXjHPYdmUfB
s18MMT1jfCO5zkRWOMN1TMINguzhyzmaHxwbbMU5fEVxAP2Ujeg6wBSJMyFm
DToENMDRe/c8XI+KcDvpH8KdzGZ0VVvkdLr2ltisBGT3IGNgPTHPHyLFo8Fo
CEcCot7HtiyMlIulbvLnu/Zs/uVaBLk3nG3IuLGZtjQKVErycgjWG5iyrTqu
5zKXEvYvPRtJqRrxXCD1KHbhi8vImsLUBnlcOgtb3uvkUv+44o4FT8sRZmi7
x5w9vpEfZ7RqDRphrQRvPB0dn/Muy2Pn0KPx1Gu13Q0x5KVGlYYJhBUmqnXH
sN+ymY3IsOobj1cFzAfjNcHMDnZM8a7asWlJsL009zW8epVJwNWNvsEqLqqQ
mOu40gtgGvkXejGXdhkZCLPixrpZMyFQJiGfu7dpGhe3iOgJJWluLAZqQPk0
WIgWW2WrkMMysRmPJXujM87dKn8p1bL6XXqWdryO6SyEsbypdfztkKRkmIkV
3mHsPhWujzENDUJxA2FnwdI++kQvoRAJRaedEIKDHoo1eQoTSol2Niuq2Twf
Nv651NWmExQ1NfE2tJvsoeC023M+a2gksb6Se6NI6uxfcIt4A+cnjgFXOuYo
T0ETZwXQVflEVCPbtXzMhXZCT33uwBQknGK6VcUjVZrBKoYleSQ7rXTxEzf+
x2FMCiTkID3AaYYVZsUMlRJpo3udX5AvPLLIYUy/5DkNNF5xs9wScKE1Tu59
HSSn7JO+styzho4KUyNlm8N2MitOKbpwTQ3PVJRnbN/zlYM0RGlzxr2g08+u
XExkPLoGppW1PKYuydKReP5kp86BORVyyGjof9DslcY7WjSlDQ6JWPwE9oXX
bYCpFNeybA7ynd/cQpsujG54j3NNYAwDR1YoxnNTXL+oNBOpEdkPrBxfs3qJ
E+JwQ8KAyJOlxfsO9t8A7AQPtf1aBMOCYc9mr0xoUPeqZLZ8iv7D9NrdkHwc
5PlJuXvCUB7MP4MVdDYL4Ji6Vu0IGytSTeVBHh56kEhp2nX+KmTtAGdfcfpi
hFJ8LiCP6GyvNoNJXXWfUIKn46DpKBGuxKXmRNM5k+kquadKtLzaqiT4Wg9n
xPhDOa6y1Meu6AsmVKW/y+plz5++YDDvVRZNr9ah/X00AwamwxZ9goB1Oz5Q
UYUymZJZfAGlbYHRAOTWXtV6bIRkNyKva1D7YgSUtmHKKqCdBjnWH06zEXL2
+o4ven7R9cWeZJ5gF2YanOV2ivjnV/S8MS+l39vl5QsiLSqVKQlZaBpfnq3A
XHAtQNXuCpeMHEGk9Wg557xR0VOXhm4a9qDRVrL77x3uOlWIuXPIwfL02scU
TeSKGU2lQw1C4VAunqdmMLqhFwHa7mTcV4k8LGSlk+nghDmvqCbt99ri4TZD
62a1mvoTAHNHLkbdJXnCVYtH+Ji5BxRqbxickIbEQ7F4zYh8xc0HdtVldxxh
Nl+A2YRlpY4jTM2WYuzkEC+r5VrIt9lIOY6uP5mOxlud+EKaB5B8KSRjUIcJ
p5OiZvRPGbw+jr6OLJHCzRERVDC+VAOgY3Tq8vEobfGMr+Uj6OQmrBIShs89
dojA74KgywZteAIerIHYpIZYQYdubm38Qq6qEniU8gBj50RoxeNjx2RndmU+
/VWXaINCuWzqUWY7Fbmwr8nUrPj2weXJLREcK3Oq5m6ucqaMHZ9j9VhjY9E1
oZtGWwA2ghMtpnrAO4C4rJg8U/PIrNbgY2Ypv5su0m4eadNPhmYgKs7p14vh
HqLxV2Y/Z6tIGnF3dL1Fenf7M9eELKlilXyZqT8D4xQQ0VbbXgCk5RBIwBXR
3dmxFWBFlO8Tolz19uHBA+rikAjAnvfAuJFnMXZJN+hppF84UHCA6vF0pSMH
SAnHhG2Z1yMJi0/DIhOm6P9vB7Ydu4w8f/etPy8VpW+/x3Czt+OKGCXfkVKZ
Ys/9oG4l9+UIr/ZmZ2jtSGt84yhYE3zsTFwwyDmt2CAxqNRQQbXYcCVGydk9
Q5jbBSf1OqUmgQszMpHZZ0v8dnrqz+wN2sBHOR7pgLsrFXsJreU8oUUEmz8i
P8oFJ1porZarwqoP3kwGAOvAiDCIIPcjtVjUpxpBr0wRmpgJH2xhuJy73mZO
Tqf5rCJQpx174s8P1BuEHYdGgeW1tVDWneKBsrHUUiUrnYCFPjjmXM7L9WPB
+GNFWxCsmN/1ZAGEu8qlFStqktMqucftvvOZELdq1geZPHpnDSazuKLH5HoZ
JTDyrRLS0OoXaWk4fKHuSn749wpwkgwIIctnYc/lbSmtjRxG90INCfBxP5NI
Qu/Gj+DvUrDGFlOI8nsAlgBT2ZGmvdqn/Muz4BwirqkEbQqqayYgdNcrQZAk
+XCdjvWzWVQwHtAvbcqKm1lPblA33zRTjiuXQ1EtDGIi56dQPVJs7us+EHNj
A1qCj2edhO2y802pMW2VZbZgI9ugGCJoC3VZb2nO/1f0R177vZ9PsZC+JV5v
cqtEk9b2vZrNMvJF/ZIZQkhuhwiQ9V7DqFL5YCPykfZBDiFYJxshIdMv6Q7E
Q0/L7I0DPo4CVFpY6+0xBbYgQ614oMZMJUTfBky3UZIn7Qr79YAbtF0jki0p
fbAMQnnye0fF7wg7gZltPFP+EOaIALGRPTvBbgS1B+R1v7NrPwtIFHBdgg/G
uh9XY3bd9zVmZVfMBiD16vF/6QdZe0X1h2csQJmwrpQsrA+fLkWPO5+jIZfV
fSjs+syhBUFyfj+UoV+P2AOlIcFrwf/N2QVwTuUfXlCg0jULzLk1G9JyhtnM
4VaoSFO37SoFDEHcCRCM7Dnxsn5VvQU+fdyr7AZxIKjZI4eMr799vroGSQRJ
9ZOepAm+tTGO9nfaBxnod8KHe5CBIk4x/sbRhbcxTr5KhmrBYFdnr0WjneBn
8jiUMyDdHXQY0kSHMYHx3xTKlYMOuu+PTII6J7WjAlM+rqc0GcTqZyYm9ieo
CxaAIdlZ6C8KpgWWf96FlNH86fqgQPsun7hNxsBLflRJuwDMPPoZUyeAYWvI
gAhzwRYdIjDxg3k1YCbhsouwc3d3qiDKM3kZSYzCi0HCvAbmOykjEQGlt1i+
vP+hug6hbMDkYRl5L+6AWf4pfuMG25gXFQEj0PGn6MpoewrzbDxA8UppDPC/
nNSXUR8OTLQa4610O9RVTraDFjMgZUwbIi6oy216STyUt+2OtWA1k7G2q/KH
nWH+zc85e5RDiG8fubUkrNU+elTY7DnOZpH9H30OUvOpqBfL9L/qmjMZffkf
6kjbaVZQUmvZNLZTaSRw0Saem1FW5RdkvEj5dlzQhZ5FwdnMJfoiWTTjBfhJ
9+SM/Vr2/ORzx4gp8Wsa0VMGMZ0t0AUjvlRcKOh965t4kiLN3DTHLFru738S
81/hAQhY0kU8VH615QQ3QtJ0HNSAOsa9mPtVTxSsaai/3wQ4xukEFweM6cTa
yjcKAiVMP+LcIWoD0EZ5aiUIsP2ImFrSs7jAwQ+4QLAEkAmLfIslPUN5p6NZ
DakXUH3MeTccsIv+2S3M4su0DFtKrzf0MYav/2ai16Ynya4CibI58VHyZIua
6E18+CVLYz2L3BlQIqivSuBSGKL6Pmox1/LXNq+mudpMKs5txlL3uxpvLJl9
1sT2gssYOCa5RssMBfdb61L7Rat9sdwO6LQ9IeftpRE6+TPTYYKzBUMO8O8v
4g35wH+POiAylUlUJhY53KGO6pUQuLXa1UlG1Cp2Q3bCEbhk8QhHbhsGfBr/
l/i5K1J/nQZeR4ZlqUKerStrOAc5lqSDsxIG4N7+bLgD4IaJ3rfWLGxqGCnC
22hOVRRJETkXtqiWzighQ0akYCwbWDJppulK5xqLW22EciDl1+MyPSzQJ7jF
pLp7vkLUjaTirNLnebEekfKUv0k5jHLgci9cDB1lqiUmBraZ5h6tB5c/3W88
an4sUvpdHESZcSuE5DNp//7h/s8RGc7YrJOgWl/pri9iVr1sVDNSiFhEDF8c
51nrobz+x/3sKSy+R2/XVgO/KGGu/1F8W2+16L6K39QWYjQgzkW7zEFWsoZY
OaKzoDMaPZ3300tqAfDv0ab4SH8V1hfo0Wi/dQ1b9Xv3S6W08TWOWKEUb/l9
CtzF5zLHCqawTPx+PlT+y9JYxLoFMaXx5w3z093/7pYwbt+Z1dKuKWOr3Q3C
CYg5CUPx0hlQQpvZrlXitfGYx9vOEqRA/zU9MFpVH+OwADgBRdTKYrSkzX+L
ReSMQ/DqUEeWjRCxaBq2vfVESvTWCKi2fu9I+uGEanRBHqFZ/SwLyrfHFaT/
/0UDCkCpU9AGgTvZsnxHrUuws3ElhxEvqGyw7RiLNm8n3BJmFXK4DUkISsaI
acyq3exBPNUNCNkkl76oKJGVLqWasmoc4JyjeWBmAbSGLKi709WQ7lOoYY2K
YLTvfRAgA+OocXwhkVQDFm5SuaHj7h7IqMTNnLWcY/HiZGikb40hUSrZQBc9
rRoaXDjCmhJE/eERl/l+vpTaEu8UqNb28R129GQT86QjwNom6KqPERq/wFui
JTGWOeTBjNHu75mJACRKtdcsLiC7lY77bQd7T5ARNw9zy3dIOII/pYHVKD6H
2ErNI5N8n5dOY0oE+gIuA/unr+gMc40ZPwvDbAP25XMOj7TmUsnHzTo66vY8
QG/hZ8RC+xTy9RQFrbUboxuR/APy8hM4qSek//iGdc9l1HtNg7gjpTJbr4v6
m2FhYXAkhO3rJYkc+MMzLc4pJJ/Q4S241ykzai1FzvQYedm+SOuO80J4BtoO
CnNxgfwWjd8lEKKjNbYPegTy8DYsgtcpHDAsnnKxCxitLoymKqthOAaBnCi1
tj9zCY3KJl1x32QxK+zcJWyNrcC+nhShOJp9hkI9x603I7Yua2W8KBpUQYr2
b1AoDF6IK2eSY0dJYZMmAe/Ft+OKtGN4wdPyHihY8K8sDZi6HVdPwgXCrQDX
5rsQ0v4dLjvfo9HMaAeIj8jiINnayHiY3xWI6qSJivQgoAhCgYTGuaEAB/RJ
ttXlCqIZfOFfSJqrOhW6K2tMWgxR1CIMKr2qmIxxD9fdKmjv+piNC3TEfqKd
2qbYfjutZpRT/WUO4tbPilNf0oukLkpupUogjKgHEHLt6nxkUeCMSuVquZ7U
q/So8e4IcTA0amts4e6MdgzjfwM2XZcCjuos7S0/nHNPacUBoFz1ApD6lSto
AsNPzOslRjvWE7FxaiPPd4puPFICFEXWtcHYAGDt/nUe1ykvFxkNXda/mtfX
C4meC60dZwTh9Ir5L/2P7ifC/nEEV0vJ5M0SuSi6zKEF/iWhWiCDKvwGkgRo
/ys7As2dS7juodUdEPCtjs37HrBlOthBpMxpaeVzewnUA3UhgBMzhybcy1P8
JPbNZ5wEh1NYejB93cOdZRoR8e7RiCpvkjzNRSCQOyMU2EoX2snhnDtsWSf4
hhV9w1ZPcHzQC58RUP0O9MR07lV7VW0II8G4TFYdzs2KELi0PG+6SmKoZip5
0WUMl2wTJrai0tdSXaFUPIZG906bUTMngMcSLOPbjoircO8XGgz5vZlb8W6q
A3JtXgAvnhQv8CZgvNpBFUaiwcIUmoB/NIdCd4Qkuvy8aFbguYzfjFp9aMS0
zPABi7rbLWPgpv7KvQH0Dod+TSWHmxnhwm/bKr4cxgtrL+f2kE+K2LIR+mTG
VVTEvQMW3hxI9ZlFcdRjvDfhALDg7DgdtSoidixyypB6DmAEzr10+WajJhR4
wfLr2fcbZsLXcf8IDxymxVM7wO20Uv/h2LAU5c7NPdAWlY/gMZ2POV9FHp/3
Hl4hCJe43GpzyFDxxQA50nZaV4GYtDqkasFYRJ4hkEryZ5np0nuBZNznscMS
tz6iHl2o4iomd+2OONtti75PzPcqLHrhlEC24/gEbNUeu9+KfAcxiGYc5Uyq
J0ypvCUEcX4j41t40tQaVjHrOEy/OgO0nltF0Lf/SnV7Oohcc+1k/UpV1if7
dx5uOkIj9hDLnoeZY4zcVVFZgpH3MhMxjH/4H5z8qMJd3XxsyDiWjA5lYYAs
agGENUMi2PBeUecoIQyQN+9187PehB7VUcbkbezsy1DoCXdEG+lwGIfUik9h
2QNzSnZqw1Gx44ahkZ9y+bxDEeow3IQlsLlPzoD1RKFZtKXrcvt0kkOwhLDk
7njdhiy7A4oG6SM01K0/mzXkAvD6G1ON7r9s1fxYTlO0ulW+lcZ5eqVMQObN
rrTWiEdIGeqwmcre2TCyX/4TUUE7YNLDV8NriX+VWqoD8cE1HS2/TUiUIBr+
v2wBz0+NC20kRRz3rkBeQqzu5VPWzi5k1wOpNFAoBGliGpp2ABfx3tIEMJOP
KnJUuvEom24RkZhhCuV8oqgdI6gN8tA21fjzzUqyRdEB1+Dws8+3rRoiQWGK
vTkhADNmfz0+/74edkHEXYMSXNnX4stCcooy3JAK+6hS8rign8NZBYQwpFrR
3lOzDP7bVVjTySTCaCaFaS6Q5nQgMy44v1HWg8sOJS5T0Xe/9ZQUL1C7iVoO
5/mYX97Ra6kvOE8SBeb48P6bqzTW57Wg8TRJds22ZeelWl7d+FyX2oEFXzS6
7UZU5AMCT/VYdyXu/KxwUBO6qOf8833JcaM8hYa+gUFmTTum0O9NXhcmaQFm
PrrdktWvhg6ERLUwU0x8vMsTLNe3Ky8HXJyFhLri1sIydgw1+Rnsdf09ZlFb
+XrYj0k6PtowVIWbQ6cXK1UfXnU3/KFYQrrm5SM+bN95L0BPVp3uInzE5LXK
HZ1ph8nLb4qAFn06JTtqQIEgPZOgJtyqwh4mAXyBHt7e5mxwzGPxbqox5u9X
k3onfWktNwVLOU1npynWMmwcFlafVKWEpluaVt6BquJeJGVhBhKuPxLlEMxf
Ne+Pf3ak+sTvmCLpyncmnqAq4byCReXmZw2j5ReCe40US/MgKMPC1YtiXRGJ
tqceDUME16rJR3gpvydoWKFuTuGptyDb5js/GdLcP4u5SU2u1spRWeoABMyv
MwhVBxL+RXHDcj2QAj9mQCAyW/qS5txpkXdjd6XBuEolLMoVqL99E2VId2T+
G0cwr9G+K7SgP3tXMfu9280WTUDs7anhvsxu+cHysc4yyzNYIEpEX++wg91O
vx5KRXmXER78FUTNEyHhNZ5YIC9OjXoKZaisG7DtffLQyAEPbfe2hB1Z8NBI
T4L5jbmydP8hY5JghW1hAtsMXZhURfK8XE76WIG8CqioTBVAdAsR2IZJ6Htt
XL+6+yFH46HnF32T4z5h+zLc4AXFLy65Rj1HQ3JaXIsezMTPiGTOYcB1zNqG
QsZx3HTjNmvbLfeKoV3IQem3woplNxubf9+stEIVAXuzb+C40vz0It5242Wo
sIfYiVwr79n1NGURnfeBzxevPMvywqr0TL0F7Cm+Sx5ay/cycMUepYrMaY3l
LXERTbEu7+xvWahsLlfLIZ2Qtl3ugEeqolNvW/E+9TFh9HAwbaECAybASLKf
a6ap2SesJkscD5SOGTMslslnNWuEIrsJp/nBGFQpZ7M7Y0+g7QF98ZRcEH8G
ede9dz0YOrjiddEEDvjLWb/CEV37s7UddIFZq+uYSwQ4UcYbKkqzSguJO7UL
50HCRm8AYMfICUOtA3+hQXbhzBTRGr+rnjDsjDvnYMsiPRoe3/KFiZI6aj41
skxD3ilYak/FMNoIQnoolf5L4/F7XnV8ZHiNXx43IqjNZiaIHDWngZtwBFGo
LU+sO6ZlVvuumfvBwwtx5QLEKZuaOpoIL1snJw/oAttuEavLSwBzd/XiM1CW
k5/GpnlcgkGtTrRJf5SsTDyxyW2S2GgvF7xbIkB1zXPOn/tWEeWOLO0buKLS
W+3pDPCDrsR2qqTBg0wfHvFdeeOe4ADxFEGllqudtz5n1D0X4nEhWeRtWItM
akzHaswIgkes5cYnLjhSPfBfCpOoTa39YujrS54VCBmmAgGzbjzg5Wt9ls4N
5iQ1LFWjrrtgpmSUqt6AGoh9HLVX5QU7rFPAIaWCpm5mVQTvNv/l95tFZdR3
Bs7mLw17lCTDU8D34BTA1qNVGVE8/xjreVimRIXNEH8Xvvh6udxuBEP3vxaf
EYr2vq8i3kwB975UdB7e8v3QFmAaBaU9PgCTMbwfPArLqSikrOxL/LBr/MIQ
VPoBvmprnjl628e3HhXFTwnDdC8OxQYAcaDkF48Uy69O8YMFKhnFOTu9ziI/
K+f12Hg62jO2dQ6r93U1guD60qOGa9uqnGBUImSmVIdIdz2Gc6Ak8Inf4mGU
HhnWuVJqWJb9nfP+VGmqBepZoDx6igKguShWqC0G1HFbZjadGpmi+UG67N9I
kkXU9jIKqQzW9vx3nrNH4CeOk/AlP/aPqVWDnwRLDwyUFI+b7bfGO+RpK0L1
5qqtdEIsTLOOY159OwuBXKgqmmfpelSn9X4s9mq2nKktK+8z+P8lP0gUnr7u
Ro53AYmrWPj9znik16227Myb6OQ45Vflzd1ZooYjPwn+tilylDn+4VcYVbRs
Fe2d9FhUw1e+9fMcQP44SNCe2KTUKu7fn3pzp98EaHURM2FqsnmEhj86D8YL
RGC3X0Xr3s4dLoYFbi1rtrhLA/H9/yjXJsMYSFetHJeK2UjoK2CyglNEb0IE
8KKmZxnK+JVnBI99IXEuvjkNeCMml6Ry1Vh7sqm4mG2NQJUVJwPxVl8RdVbd
oh+TcJXGGWEaWNeow1GVV7QlpaMb0/JlL7ccPOoc8x5lTd4+YhE8sob0Sp4k
3muNWpX75EQLqNhQveL52PeRDaqtGBg19NHPy1mCqzf3AkrDizMl29BNHCOz
Ndv59eaVQjV3lkJXXHNODm+cujb1tcHbf3RnWIsu6MsoeERN1qMH/1Cu+yZE
TFrkAivYkDr3inkMVyiy0HJbTN0Uno8S9v+AQBwsq3ZvCVsm80jDurWc3ThH
Al2E9fZzmuHcVTB2ec1lK7dHW0CLf45gGnq5dsYfYXXwOosjl/AbF6OQo5DP
1+Dyua/rwei+c2tV2kyxy+uN1ThUmu9P1eu/QRxs75jKzJ+ict7LKk1fWsTl
JGMz0FGyll7MpWT4ZoTm+roK9YHiTmPdpwci+z4gLcSIr6S8rhTdSu8Teseb
XiFUgEbZnbob3VisyIAnXlajLLnammaBoJ3UK71fk+Zg4JyQzgSDaHI9irc3
VllUaf7fShBwr8S1XIaDMFgK9lpqkUp0nNqd4sFvDDTEd9dJ69zhQe9VBy+R
aqJ7EczPrR9iyNiKQQ2NtcHVq1gZx2ua7k482gq0RO3Uw3qtrV9sclxCYIgN
TMvCYD6bOK3iyJlueyvJ0EK+M9bxGbYF1cX9bWLbFf2KXKHtuIK5dF4cp3Pm
O7IModqEBgKBjNQ95oLfvroQeQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+lUm9sP+oaRfloTeYTqt4oDZ8d89FzEhmO9j8Nf9j8xOs5VkV1ZUEM0amMyDiHAn0u8qY6GFaHZWNYEqIhD1LrsIZ3uI2XyT36nMOKwkQZUwZeqQJc4BzahCAHHtruEWecJykuQb+Wm2iRIkm7UYIKd4ClWYgkrQIGTnc7LeC2cgw2v1y9fYVVd/1lH6PIM6YGB4W89FtSmGw0H0t4a3Ro+6g7ehoF+tKIku94KlInY/QmSOF+uI3efThbvnc+HrwWbyP2EQXCZLcyqD2EKlcq+gZzuTMVMvIV3BVavuXrXBLpt20h/0pHGicHw1mINu7aD0EvRjHcMQRfcRajTBi3QE0eRJMP2N8vvcyIYfHf8e52PEeCK4sfx0+NNjx4vmbML7QRymqW11Y/JXhGM7f9wI446AUk2KLojXQ/nfIqkDlLghm6WieichVGuscTVrgWi8YQU0wTAFQhiZ3A8F59dndq7maRYTBQlwbY5sWOnEFxJuBhAX6yPcn54n2N9uQD6+iP3feF2STo5I1UdEHy16g48HRWV+vSBcmW1ZfAyyMUH18ZUQANRZIm+nAhancMsUErg+ORfcs6Srs28R1U6FA/sW36sdpYv3AgUHl1NurcGnKquCJzzb6IkXJv3Ohn9uk1+gZWUYQ3pB/CR4CJGa46pAXh6/A0C3HCvAUKKSzC65cswjxIRiCzohOO5MoioNA0A9MhQpVq5cMjI36mRalfZ6K9+TMjqWIiS6tOhQrBCcjfMnAtL/1JrPN/4ba/vxKL3ojdiENB7QOJXkC0x"
`endif