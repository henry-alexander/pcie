// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NIMEse6pnKC/09xxlDkdExVIJ2fZ9jFUJsQxiha/JrYHMSYycp0C5GpCoUzO
JRdHAMrf+lEhK+WT8+2S5Ep8DpzUvq/yxOpOqM/RQRH9wOUs0/Vd0FMbtnvs
WksqBgR5hIHpcANwo7ZvxdtPlm9XWp9I0EViOCZAdwuzoUM+MTRZ3MO3mgJg
lzoo9cBYiHXtZOmD0NVB2EZx0cXoynJCU7bYqcz6FlapRi8urcIKjdL82v11
kjIIvfpyNVdBrIbQARiEYKff0v4enYJiVgsDStTdSYNifrMzteKhrMMUzb+H
ZgcQL5mzpD/JlyIoRE/+9ZhPjL/ALVj/6mPc0Wdp1Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
K1YNSWIpICZpj7eNH7e0uXuV8PnIeLHdm8HN5VrWCXwRtg3i1vjyuBWg1PF1
Z0tDLuC9f6oCeUEnyu5uMzA8D0NILub7oRDSEhJmyFuAnPe8Jp0kBIYHsXtO
k0hMu2TM9/khaiklwDiWy4vNMlhl3k2V+pPj7V/psCFgdl2zFvA/yhf72hyM
fTDrZoPWJJDKtQtatTiHx3/H7BsRmcDCRUjm6CRxqMbD6N9sHSf6BlfdDozJ
LGSdsyG5uu7D54E1J8ejrIRHSniqFbiRvdG/2cBkFKetN11/mlCbA71XLjsU
A9qGe7J9VIY9u7XKvvzDnJNiC8FIpD0BnGGIfLoLRw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iguzfUZqMNckmYDRD3kQzaooyhdky1ZV1C+OFjOWxBnl56/NKKI82XMtSp4/
9zptriUGgXLh91nz3kVmxnVRBcRu0UfLSFf0NDoVaW2U0dv5+2b67QwU/I8Q
exp4buxYlSYu2mP9eG/mg60MjzYdNf8pGbg8+oWx5l2PQ33EUX5H1dxh6q6W
llh67609NXxcS2xHQmrnB5polFMGLpbbUxKenN3q+KP1sZqQa+11PCNNrt8I
DnL152BfoKtizb8S0GD2yxH3bFPDTqLmmdZSYnL8bIprF9eOXXWDv45bNGAq
2MOwTSXa9G75sD6P/Uex2wO0Q2MoST905NDrjlA8bg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GeWz1xvbXQYL0YUZcK/HPN6xpzIChur9PZSf7xWqRhdrmNO7I7NibTCTtGrg
Ay5CJlusyRrEYC84+LHY3qmC0Sh61+jUyl5QjdHH7PjJl6sayzsrUq9T0aem
X8HcqZxq4ZpqOA3USHvrcoBNqI2q2KYC3jcWCSFG+4EHbDRaqyU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uOscrJGs/YKU+Om+RA6syuwQCQvTagTSAKx2zCJjupqpNqJIt/AZYROP0cg2
Rh0bcvLpL5Ysh02T1FbYCqXyz/b2/YyKAQD3uD4itsICqvJd1q+VZzc3w4dT
YUWwWwfSe6p5hbVYIwsu3VFW4kDgYF8AfeGTUtsnWPlfxOd/pnamgYxKnRCA
hU3a/q4n+CGpa1Rc10GwIuA/Pb7O0rLOPBbNzYRQSgQp43vJl8hWX2qyQqvB
u1ym6JGe9/hUGcyNyRsw8ZmsDGCKRtWCH7oZxULziQmRM2SD4OZDCz++XmCG
E4WEjrlZcKuD7yQE56hzlc1KkChTgzjjKCd2q/Z2H6bu8VTB/Tx26IqaNMMF
LbeOd4es64+bUEgVTdEvuhgGuEmmB8w5FdtN6DXH73h3fzku4GfF4CaTA2Yw
hV4RgiQ8ywqijDFHKdCXHkiWmYuUMUGe4KZDKTSby4omPeAod5Pw1ucWR29A
QGztik3/JfAsPsBENkMGhmMYs6II9w0x


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LInJkuP83yS0PdGwHUKGbjhom5OYxsG2fMw1Id1+yzsKM34FLRMhNxFwcRAd
HGKPL6V65MSkwgZo7dJXVaS4eDVDzuyGWLLNxjkcUg0susju7+y42UbnptkZ
MewdMwfkhGmWQ1d0BGTnEo1da74LFYo2icPE+riP4LG4+H58gWM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L0upM0pLYUPo1mWhaHgzGO/jpuVnkfRX5rHXhxi4krMzwizJ7mf3wEWsR04d
gCaK7Wq8uEMcHKkWZ0W43dIqWqbpjdN+Hn1HuJAEMb0iro57S9HGfJtSMmnf
rOackkD1LOUSSB3LgJLh4enzSZgLofgd6oqRupnvfF2OzggCLWQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 37040)
`pragma protect data_block
MQlVRDjk5XTtb5mkF+8aKJhRqxv6sNHNQ5OX19WyfchOQ8VCjO8UWNYekAX0
KjMiiOjYOyXlFmmwhgL8Ow2Em0gzv3rjOxWrhGdSPet+0lx39Z9h9mwhWOpG
V7LP8zcv6SRYqPB46oGkuhRRy9bQenAHkpFpaC40HvpqIYH4OLdSR8wNn8yz
9B7gc7dev0R2+BY0qskDklnQB2oe41avbiHH8MPBAM8BG2ns5UeWZDm+X3cK
uT/mXFt2EMzPwUjKZY3PTHPAYwQMA4cL8QZRw1WwTPAW6djX9x6iQ/IavzT9
SL5U/LiONlNT+mv6EdkGdEnCKMJgquddcI4Kq+1O2qVROtO+ABV3VjKaFJR8
EfkwMr5PezQPHexzhI8ocNyBrIhqR3ZF+1skkr5AGUqfB77jVyNvZV2p+3kX
6qCitqWueo7HWU/vj4FFiV1/VFn65Ai3bChfad4ShJu9uQxPym8DWd20be3f
EP+RwcVB0hTXJ/tV9w9SSJmsaKkyYvs35hGjM03o2bQd70X/NuEXrALoVG4M
V+Pul55aOJSffk3LteEKXU5l/UBZx7q9g1pEQrPGAqIkYjBhjZwFo1X+tkFo
H3QtQ55pZSlKWBTXs2RCH3gJkW/hvfp70SHrhCPUS/3Nxtyrb00JtX/FcB29
ntVDIRhcexzorJmDyeRK+qArkr6f8xUGVhCXpl29+OeMWZPVLkn/aoMR/5gG
6BZW0RUlGUNEDHx57cXEtlLjM/L6L3eRNpa5jexTTDA2SmowiobbFkOo9PlK
UgKrySaJo/ucgYLmXWqe1RjzIlwU1lHDEsiGt2uWzVsYUpjZuBl1P1Gv335v
VhuJHoYi/PgbWJ9L5/qgngJu1iadtT02KwRXcmQNaRiiOpihv4O9qbCO9JDH
ZjedsG2DW9o2lk3hUw+QdimkgcwhdUqFqVS2DS02BS2chHtWGsMEcbvQt+sU
VwGEkvxL+oos20U22aq0BmG3g5IdetJtXslSeTh7gCuGKSj+Kpp1r7M3lPz6
oFtzSNqkWTXO9C15c1CGcKs9WvukcwDMA3SJ/xZRpNyjXt+Y8bbI39YeCA2s
8oDthp9zRw/a0JwdK8ZogTdY92l4hm96SYVsL5u1gGccxzSFZ1JhhsbAfxQp
xIuejjpeZMB561qxuYxrwt2ojWXqrjjRli7K+2bZgBoBghvxD5uWHfd/nwkN
bmY4Vhy/ansI7jX6rxIhVSLhXO5r0YX6Pfy0N0ydXTNpkaoBFW0hLTZh//6Z
9GV3wbZKPlapYV8jm6lO482saOOWdgOwnqakzyJprrkzF0BuTqgHwtfYPJvd
VmiZPpmjV78Y2uafVjocoa173XUOrFsX8OoG4P8iIxz2SMmnLKWxWg1nAggf
Mg1QOs0OpadBHwdWlQdCbh5bf8HcnReJPXtbeVDRox8XSkmn8EgNyMDnSKvj
Oc7CUfgNzF+hfA6uNLjFnfBNTEW3X98PGSHPVleRmTKS3KP07fr19mm1REAB
viymqCcaI4IV7hQExHNfmLCqv7U/N8WPFyqefzk0VaFHQXYMgwymqMJgbqP9
Tp7SgD3mrEZsewRXHXyLtmW9NieHASryXDBnYrUJjoYzKu0puKIy1OeDjnNI
vBwFBiZtAur7Gq+neieh5zKl/OgF/dqAF0cWQp2jweGkli40cWjxFYU9m/6A
FgO3UfphpxqRIifKkY2yAoplD6Q0TDK0Wx4w0Z88dHL1XdQQujuOHTvxBcd/
b36ItkoxYg2mpPv3AGSBynnkHbcOJut9KcV44maPWuAFi29n3UsPPWcsrXZp
aDgv19jUJd9oItuIrGLV+qPeCUbfCn+SqvpEdlYFd/Nvz20zn/NuSsktZ8NU
+Iui4fgPy6ei/vIgbdGhycmzM02wvOmeH+5zK7vSgtM+M56XPSeo/ZMYJS09
VdWKNs/RDX5RYl0a9J+HXLsNpgYrDPKLatUJbWdrkusvfeTYzkgux0oMALzT
0Djg8EIvJOgX7boFBMenE2foVwCJL3xuRyHEA92ppONhTWl5IxZAyCUXw446
DzH7AOA9YC6LYb2sSsYpYg7zVGDTwHvRGM2Q37ImeaTTSmprV5bG9CpzyWJ8
cq/FNfIQbMdWGQ6wQU52RQ+bO6YoyCC55JA1HrQO7LrLEqXCAfpLGYY9wZS1
WOI+jxq9k8tc6SjrAW4plbRL5k1jsjynSSCIK4vLMlaS6Npwmn9lzpo8Zd1C
OO2kk0U0iri5Dt+NTcf2H7Pxk/o4hkoIaU6M9nmGqvY9izFa/WkKFCarKY8q
WVE55xGQgIPdfcHyWGQ7BlqCiSOHkAZNzr58Y/ysSnbprZ2KjfzSmMTrElJE
xRJaIZHppnKY9rPHGdN3mWGyQAugqZ129ldTXqxqekmHFTfzZK6sIXNv8RcI
fhKN39l7sGGbQpNXDqe+xgx8wqSnRK5Bx3vgIO8oWJ5mS9CMDT5yImsxaW2s
0PsT6MsBK/hMDK+1B4Zj6bYVluu7NbtLjgwIVPwmfoZ+W8R6TfS9vIRI5MZc
tNaZtbD0y33BObECtP2sLV0w+VtmgwVWjPWloLtlLD2NgaPKx4VE6ChGjgYD
6JiAuSprTPfsGDINHZr0ofTFiuxLZXQWAkuKuXJ2W1wsecYU129v+/DNAcL6
tyoThz2KQOWqrJROsJTiPU27r0iTSWPyhU7WFHwDsUBEUJOm1bn2coVP+3Yw
aTb4BbZdPeF7cXqHVX1GsHb8Dz26PADPUZvExq2rSjGqeqQtJ2KdvKFCR48k
Pf7vdbiXylMmqDl8GFRlkoWpxQDqp/XpbrL3TK1TkVnePnnmdR1E+BTJGu0A
NDY9DF9QY03tevw0jk6HQYZhJ9CX4MB4ga6793XvM5rHUQ5k0kFjoIPuXS8n
Lib30o6def2Z620pPMdVs8ZiWZSTNdcBk3Acj7tj1/79fhkl9UXhd+r81ndb
A91VFeYfiib9jP94fIIkmAfbOpbV7iGJtEO9JGfhvA7ap1DPhfaMDze3Lg0K
hMBVLJCnSZErrw0tuUTUGh/b/bB26XfZB1ySENqG2rnTYwrCbSJIS0wISLGN
Grq49VcOHFBHJjyCgYxHEHqxqGxDbIYZ3UEh7EoFIp7I/MQLvzHX9RvHapxr
gE2TG0wqJ5SEl5RFwN4+FFYVwjUsgB4YXbXPu/PXOeph+vhUSLuEAvZFs/40
SG/GxvgOjcULPCOdyNAzhdWidj9vL8uHzUtzzVZ19AAVY2NnpUyuxJ3AXryY
DStEcioWep3IRyB9QlcN6cnjw0bDngl+th7h/WyAqMD5Yf/6Qn3JTCQw8DNu
NawjELPW1dcIw4ey4qmiWic6ZqAmMxRRMUKeT/nE0rRODhHFG84KAB+haV52
KC8cWeFjNVRgpb1thkzWikJ9G5M9ofaT17V/76BpueLFH9H2cU8C1Dzx1gHD
vqa2VXiDgoKcKG1mm6YIM/q/NC9oSL1zeQ/R7slRjoNtTTy/uzEMxQUpSnev
IPEt4oBgyukBPReJ+Ds6RcyvlSaur9Cumb+Vw+1Zk3imZAdmBscvMxH7olkw
sE4gJUn3A6Gf2Qm7l2/CsffbUrJgOUXbQe7OQAk+24pPqUZCAb2z+hQuK1ZO
wUSyKSqCmRE0riuaF3DCzz8KBPBwUzhKKe3n6nKxET3ehZezNUKaQo/RPMSs
E36HWTlvBUu1Eb4E0C7/YU4rUMtI7tLkFxQ7K4zRehtufprlGsMCWuRduqwb
D7v2CFxhPPmY6RoQDxyelrzq8bbaz7ZJBnPGp6ls+XK+4rDliA31AJ6eiaz0
SSdD6IDxFxpQUD0YvEgZb//02k4v9/zJBtqKIoAjsjWVtjR8m5Nqnl8aNwzm
cDC20jmOl83UjmTCrTsdmQ4tht0cJgHBrV2XSl5NqBFca6IZaLaly5uCxGUQ
+lAaPxb3VPO5IFyfH7CnV6Rhb9RAX881idxgk/JGpDPxemUhCAO80gx/X/QI
lv9FITYNKUoKNZbjNGHEy5+HdRgrredg8XZdY0AoymGYge+KRdF99KqcLNuE
ObeLgMvpIz/v+9kYE3HgtMsMUTUZNJ/bbjhptrSdYjGy31RYjWXPepQW1LxE
vdP8IElU6Go2z0/f7/kBRCo9bL0btUup12oEmQQX3Fz7iNKZ/NQcOw0A5VS1
TaeUia9bas3+2HoRXzCGCNQMH8/vc0Ge/iY1QLO+g67AoLcBTZPrMzYrky7a
RdFW+1ltQBISaPtHocxtZSxkM1di2NZ20Pm19wBXC/QSYnG5icQQMw0W77Au
+cF+CFjW1Xm4ATKT/MVgj4ZwEBai7ml9S3l4ib0T9Yao3jPVLS1jtVoHlyYp
4/mdg3cm9XuVvN17CUJnLxrz9xvXtYKWNjfPomMP6FEAswXAjvKN/6XCBL1C
2yv2zNejC0QmqEnud2CE7/xiEPI0MZ4hG3RCnEurUCrCEK/ELZGZMnourne2
npjpQWyFaQa2X7OVkPjmM3fcCYa1I4uZeCf/M/saIPqrq8Xne2CcYIlgyWUm
GA9FU4BOxgEljh8la9OAEEQr3hCDjKLKGOVreF2RxhQ3dBepeaDMPW82yLWT
F/g4aFtgGyyp20Mt8BgC9KG6uG6LZ2dWERmjwwifOvt17OqJ5NLHajPhKB66
vNmSsCjMIooqD0qOZmocMXk7veFy7+qd9nqQTg9I6OzqiWq/uXhiLRAsJM2r
EXSFLwULgAYOXwfeAlmTOezZeOmAcyGxpbl7TPs5m7Vrajzb6kZftXMHVxUw
/IvENmxdXq3E3uApw5b1KTlEp4BePAciID2O6tY5Ibki9dxd6/zhSeGs67Lw
fj3Nn2Q9eijNv6gOwVu1ugGbOv5z/dTiJGg0tOgDWmtiUumy+HPJ6VthpuAM
1iQx2eXKfRXQ3L457ZLcwkqI9AL/D0OPMb3s5P0Us1YAYB7X2t3GTsWFE0SN
IfHaOOcmhhNPSI9hq0W0qFGwVbq4uK4I8qu//Owsy8GYJv+QZYCdfG/VoL4J
hbF8R7f0md9IysTpX5m2E46yVqI9u02Tt5HacvL4a9o/4gQHz3P+F55iZ6X3
E9ICXc1NB7oS1APtEA+kfr5h6S6rx/dC8diVYlmhbHGoiSY7Lqk8uf/ey21Z
zNKms9Kn0+8fTib/teZUUOQtjcG6GW5ymMd+NEjoa2yXm90P3QtcFzHMuoNT
c3O6rxatEUgVUyUtcfy6o1eOzPXFHbHHCA2Opa9bIxS07zYlrgm1uqpyTG5v
69SoiDul/sa6rzoCWWZLnjFnXOEIIZ+qKhigR2wDYiYbErR2ZotUpMzTEir3
U1F9Zpt2CIT2wnN0ehHH0JJzCYfedXzptn1UdYfSz77d7rDclyJcH0htGaIJ
NB6sXQbUUIMwDZcz0VBM/lqRFV+UQff2Z4+WtHMOIqUa2D80MlS0qO2zC2kX
nIqBSuR4CVytMQTfWFV5oFm3+4wgkJJ/ciljAmoFTQOTLtavweFs/QSwbV8R
tn3J5eS+6nwG04cULCknQUKpjRROGa/9wwspcRRFkOLtRK4sXT0S4wbLldYM
eMcyURaQt6FaSGBOMFKWlouZQ9E5tPq8Ofm4i0XLoj4uL8+4tZQsxBmhHIvl
AEWBWkuo6iV3z99Q3OAifkap2VZAMAIjem74iHFAJ+CpsiPPY/wpSFee67oM
I3EtCFW61l9yzUVYpL3TG7+YdIsoEp1sMA/bU3jKEx6EsmNa6O/7L42k8/Es
dz7a8QbBCfVN7C8o3+hvIx+hIdLD3VMuLuj9LR5MfXhE1AYpAUeCN1covE6v
kLo53QyYH0yDuM3kCgTmPjvuLSqlEmbCtbee/w+3GwEtbkUUSf8do7mic73P
j2FmQW+XHgbS4QSKH5PAi5oOzsrPU60GvCxd4BFxzY8dI6Nv2oFP61G7bIZQ
M8I6TKS3yXl1J9G2TLuCcFSJr5YJX/JFBGRWPZmoEHTsAOzcWLUB5pNxQSIW
avnLJ77hRTyzuSQ6yWuGLuYq3z21IbzOb1DQh3zWyG0yrx7CwL2iebxRl+TF
8n0PJEe/XH+DFl8ruaKl2ROK357H+w5GZiq1ZyySrBS9UktqKXPsjOUd0BN6
9b/wz9hN33sLiDRsitu+TkAy4qg29bhX1JR1snc1bts96uk/xmjItWWkEX1O
4zRwoLaLh0i3IxlF96ooHg21veN8CG6PbgJxx6bnwjJKusXU7/UN6g8IMvMu
v5JhoPpfZa+MY+StS4kRiFqVBeSZrMe9UwpxbAgV82VMoHUe6Ay3Yn8bGiSH
ac82F39SSIju6XOISGf6yBOKRO3NX04k6mu9h1/rtM6q37xoW0u0sfCt43Jl
tboMkJzXLkkwd6VOeRHF0Rps2kgkeXAZi0WnzngCjcYzLj60a+yKMKMp60HY
iKwAv2H8NI+QbdgDwtW2XlYDja8btfETmAr6Zh2VFmM/uNdcLC5MGfMS6ZEs
d6OPj9qd5bMXjhMy5Xxx9EYsteSk1VHBRG2Isdxbr7FaowI6xdjJ2z5CC/hw
xNjmsqikXch+QGmwIsnFiMWuRnvYUcnbgVH/q0/9SdkxY10l0KewbG9JYR1X
xV6wtdPWEgcPd3R2KtRaoS8Ga9wjh+duxWbRZ6CWxJfapSpRJOAD8HjDC4wN
Tv61YUcayUban+dfQxig1OOwn7asHOW/l4tjknoiOtJlrRFDeztBiNwUBrRy
CXdVxha0DNNsvykdHxNu6N797By07GBmBanOwX349mFl+HAjBzZme/O9X/9+
Cjq7C1oHmPIp7o6GJ8ZecIjJpClxRlm5noJgYtdDVyc/pOFiiqtxblofOdAS
liVRbNu0QhKMqY8IKauLu0PyLrKeDfYrRaz3OsCTs/qQ2QVPJQ8bAIdBR0Sv
DEr49mXv86PIzfXbXGyYfP0BGIx+VKyuxoj3QshhafK6vBCdb4WeSnA/jUqP
/abrskbP5IJ2W0O8w/4SY3yM9dAdl/hZGp8rh9BvS6qTZgiLkriL+tcblC3x
FvvW8OXUoTB0kI8pMAeupfQ3rGEo80RxHp64B7K9pmnBkSrfxGdwfGaEjXC3
D7PnjINjSdd7talvjZiNCnvUS+9MPDqJKB3y+zNPk496LZRhjJ9ZQuZD1lgE
d3cNIwHVVuvG0tRxR6lZ2m6KzOh9voEKu/wPSOfRhesowPfZpBHcVuIBsdBQ
YCrDypmofjHqUZ+bPbGTjelqXYQZO7BJ74xqVHWyJd3pwJsk20SCZQGMBtV2
HphrQXFU1E7EIWg10p4wTbTIKd6oUTBHo7iBh/GEYhhOvbZl6w+/Et4yilVp
NEt3kq/AGoq/3eyttTNgmo9Rg4yodoYxua15kEtcl8E3E5SRoln0Lf+CISZJ
pMiUFE/TRAPYJ4F6PsHhZm7uSG5dMwltnpEUVzLeSXrpzqIWhFxUHxgmxhGI
gaHditRFSB+O5uoqyIGUAmIFLXPwe8Ie92iQkj+LMQ7IFhzrqmrvUqFMRNuj
RjIE4MARj9exq8/87Di7VnfWuGPUOOKPIxpVgQykwvXTGP2J2duIBfGXNAOw
nezLh5LC63iHRpDMDRureht1BrCwc1DYS91uGMcb6ZKSLH6WD+wIFeOFhcHo
cy8UOobTXuZ2LsXQuH1sCDrfQL+W7g6d60yJZK2tOjKIq/w4+LVmBPeuPVkv
of5F6Szjq42L+yVrc09hf2SkMeExyEbhGrWgptR9wxTUvuRjhWiytU+HgaAE
9DgnVgQUwfgZ1MDpt3GS5pS4UIrmkEfs8f0phFqYMgBUSPAt5Z+GAtU4Is9e
knRmBLh5oK42LY+Eeucdv2LMrAdQYIVUGaXFTJ1hekKQglzdkSKR4fquVj1w
ufZOywPFWonJIvsUoRo99xoACSefwO7s8Fcyn0v7rT2Vri9PY7lBWBwk8s5s
aNgjDpf+vsoPESc0/rj3RDRse6WO+9CYm9ahVTovx8JMWCyGqLON9r/KAlXH
MAczVY4yyWmEd7jvIB6/1fPzCCjAsH/4fVPVahMTGP8oGw5B8p/wAi4YSojy
RFVU6+DEaSt//BqvPd9LIzEvZZaXLoZJIyH+q6OnooFivJGPUZry4YCAk+Lk
fJgokzxaGNvB4Q74us6ICdWBYuwH/QiV4PYNFkGkKNBdNZMU5a0F+3wEXWPW
wFMPTu50o8PYFU/YRiKBEEZjdASb3ApgeJJLay7ed/x5BHvDcYwQlK9A651f
utPBh+gA/snixMDthXdqpJY42Q5+LZ5CXYrD/BXbZ5/7330i0XN0tUiQAhe/
1R6K+Jh8qVcoFOcSzO/pJ6rcw9i9Qydx1ii8fupMwHxx9IYxJ9fOy1ATLLdQ
5oYjpd0vpXR6ByNr4P/rRUH/dGZNXleFRm1myraI32QQdqLyZRaa+CWWL4vJ
b69sjDlTORrZUKCkAuGMrkfCocXx2clFmGOAb+J+6HC3olbyx2l4bnLjchQB
GIi0NT+UfjLc9rVMfvnjzy8FL4VQTM5rUqiKuYcejvrNoY/KerPf1Lpc4/a/
Hkujr791voB68cP3MSiPMZsC2UDHWNAiwW5sg/P/6VcD8XbMthZ8GVvQO3ZK
Ka5FN4anhcSXACSnOkIYC2Eunte93N2xUV73UJ3jDOlJTds4qV/6PpcI2SyC
26h274hyyNp5mVZ/FiaT9Z3eU6Ql29bG43Kf+ClpV7VXR7H7ouAGDZ6gkRQR
4ODppr4TJs4JIeCbCerMbI2Jm5gR2ysFMrZ7MGnNdSF/omRdXvB9+FyIEOEH
/2GK7dLgmorretWUUPTt/Fe63QyvaHiRfaCehtfVBWfIOJnBpzC9byZrb5l7
QovDRCX+hNouoh46vdSzUJmgTM2iHlDo6epPts/bcIXZYVwNl1xGksNR4+hN
ynQskqLI0m/LTh5bANGQ4DqeDGbRHFfr2bi/EX6u1vt/fVZQgn6cawMs9FMB
hYaGPntCYJZiTvrdthgCjUc22UeF0qVqrO8EKN3zBz+6zt5wiE4dMbcaiyKa
7NGp9KF88Kx4bpvgZj6lA9O/tzyU5vVnJfRQc09Q/YgfH6ACtPnMJvAy5jLl
RzPeEtttIJ4BID+ylHhR0MRZdRtdXyjJDOHe9khVU6/Rch6WJA17aZqM9Hw9
junhtoiOmaiR5g22BfDfdQpl29Klw9uwv3uNTbR0r2SZvUeM+0Z30tNBBVwH
ES/zCoPp6YfW3S1h8quStrZM7r6Y1rSUohoiXFX8hgp3JVUAqOe0pNfODggj
VgrMqoeQUxn+5QG3jm+eTxi+epjKq4dc1oKvKOiF81oHGUW8MbqcbnCkvpSn
/izX+AinmqH+YWmIa+IsAz6Xd2wyF6q4/YaOH7CEPiGuJC/zE7LDK6tU8mN+
JTvLfcH80KMy86VALeFLWajZj20mlHkSeoxqd+iztl9sQwiPD7TBk+aOYCz1
4gNMvCET6fzZ2TEqPiFoD1uYcGf+q6txdviRKAnkWeETeXuQe5QllmjOTZSY
qMMiC8DDi2ULE9/uftxGSkuY/sBGFl8GVyheYqyVBPui8mkte4ZWxKe/Te3k
AVmzZA4A3WUjpVYh3TWu0xMgpzLhuyiaVV0se0uUQQEJ7ScgeesoljA4GioS
EuFHTWCYZ52VHPqAJcirNsjd74/SUZSI7PEX0G5uuv44ausxsc7+bLusep/S
YL0xLbz/b9rvm3hBdkvNJhgqiW533yGZhBgTUcQdgBgs07HUae6hLzu8Tmfg
9VpVzO0/9728um3IUKBWNcAY2LPnAe0VS/pHhhVIBCb4M6BCrPgtoaPx8cpn
paI3adks72XiIG5rOO/ZCyD/a/Ii+j4vxFUNgtmpckogxujZxrJaJGEg5OaQ
JzO5D4mQRH7dDjEOy9gv76PoLlllQd9vgo738HYnaLPtGS2fmOhnPPE3wCca
7r0Zr3b0eshWhnntrg3Uc+1P+uomiwj8nTPv2jnD7D9zRxZhTIzaxOb9dhip
aZMWF3f17PCBHCylTjBhfeGCCXonNKkQMdTVzarBBVh3gXmSAQ6A0UF9Z28k
BXMhfp1AqFMsbvFO6tKlq78YzFFp2m2Xcsey/duG6zo9HTFtguQE1D9RKcUZ
EHGzd7mZBgKnWpWMSBsXGWjK1cKYVtM6+k4cZUzebW4LUKTZuQipa0tC0wpj
Z1JSo2DqppBKlnARFsZNrVRuOxaTz5tQgkl3pox1/eTTUWRDVeraxZy9APon
udmatbj55ejQk78/ngJLTFNL6wdAHW3/ojy70IxfFbbE3Su4uvCmsmNC7iuX
J1a22BxVk2+227PSI/HJwo1uB9beGs9prMy3BTqDT6RTVXkVEzTqzAd/IWpE
mJHAUo+OxDgDzijJyFwhmTlS97T5voGOVtzxG1MpC3J7FXsqadmg/0ujdhy8
8lyhY+z+G8ZnS0E6LAT8truHcAgD6TOxXrVjrA3JGp1hgi/OzxB5/zV5TSo6
/eZVcKBkpl9b0WfjPFduS0qxmccmRbwwa2xy2QAqr9agGpdBr9/RIbWj+rsc
tRR7aingyp8PMNiDX8zDBThbHvLrSFmWE6NPgFO6ZU7XFZM5bsGav3PSXs48
fsm8BbWvUKuXQ0NMLypvRVJKDvFKsWPf1nAMPyYE0d9Y06MAKhKTSQ+hPM2N
Y+aa2Vj9bCH6CaFUZb7+YUYPO6S6rGJrEQCgHey7Dl8JTsxDZfhVw1u49Eke
NnVo9gSnpOOaA9VlFcgQ76XbdB6JZnZHSmDVVNKIB89OLQ7GyCmLGUOvhdsX
JD6AYyaG9inwTPLrdUYp8EmDH3Fd8GgJEZUWXmRAz1TlT1dKYL7UNjt6wmHT
MZlhWXvYTyxxH4RMwdyJ+CqjN63CpyxEJqAnZuLaL9xkIB8BoaxrslT8Wqx3
4bgH5PxVWh7tQUzjs2H0ikRB3eA0rqxFcCqqbnYgzcHZxAv2B6rqCt//0siV
isrpK0NTNurybgy0nYmnHa0wM8/6wx3luQkvqryHp0uhSyctnSEpR7O6WhAz
tEWKByduOFbFOkA76+xNREebfFx+dt17drsZeZI0KOSV+EPZWCznogzhXo0y
FIAT03/LEumatoOlylTzQpZgyYHXsaB96hhFjiyhihLBeTgunmhqh+u5eQkJ
J8oDxJzEvX4HFRnIMETxIl8+EtLuTMJDb6gteatYxkpx47e3YqCy0WUhYlD0
6JafDfMk/ZtEO1aNEcYnxaUY42KSpHgKP5dn9u1XbvQ1MSJFKrGHHMrotV2+
tgYL8t8i1j7z+etyQM6Xj11JBYDLaAsSxpx8jD6DwoP2R5SftlY7Qt7LRv5a
ujYn93dx8MSmEA12NQn6LHsx6ncr0MVtrsbjcKX9jt/Ld4e8mJXi2Ny9OGAK
jGhNrj0RF3m2sKvp0psbyff1Heex4xRQIQDCxuoEVMQOzoQh1RoApw1rEyJc
fWLad2VM40mwQQCZ/pdbdIZyzCm4xv/0aQZZ0Jik1WbVdKRGES+eM4+HFFid
kcKgbbIat+xc5ovAinIpqnjW0+t33hjIo/UefeyfjcyZkL39l2hCVYGdyO3y
Ad6IhvEY9pR30CEreVpUsCDtgJXTGinmcz8ZlTt8x+B5MOJclu9ER788SsPd
jPClCKIqLg8qzddi8gtMZ9/iViFnTM/ALLcvy+33bmXEktsaBc8c4aJ8ZvjZ
9V5f9qix6s8/BDpF91oaJKnRu74BKSryZSr6x8fpoWsDyrJprlJ2JA6/i9Hv
2Ugzag8qk62GiSE+Z02wLN+NfNEiGgFCFijI9hfjgsYfE2NErvELeYtkASVJ
zPUr/V/arClNUfySmR4VX8Ncrq1Q/Xr7XU+I+1ic7auBJRXRwFU/zIVirrha
htjV06jYt6yhRcGQD1cN/MhYNVAfBWS+asviV9Z4fw5PEnheUx0Ezfy2rWpM
VzSUe0TWn/RY7h3iKtCTVGNAuFGE2MboCwyHAEJ6nDCeTNdRLbmab0KO6IBh
gNGX6RiswV3922/1yxgzCPTwJMuFUycjt9dwNLYV7OHkRfJMkjAs+Zn249RG
4LiiZ+F8ZfMKnbSf/lr7ArDrU/onZ4XY2fwpJkw33BKoM8gqOY7ZF9A0mr/O
Azkw1Q95PPfSEjev2eg3d6UEBJy+0YCN/xirWjjJiqBHVvq939j9n3pQVcwU
ZxbTpVDNzoAC4Pi/2Ri97B347upRXafMThAFi69DunTHqMtqDik4uMgapzI/
JKMpQ2hfQgxVif+iirDAg+BethAy7s+Ao03YFf1hiC+I4BdIIHx3M0yp5wmI
3nBg2q/IeVMRkt9QxopgAcfLnw5Jalrcri0/1JWEt5FYc1+ujoXBJpVXZKkn
NsCo1ZB70aiX030SVrYnwtG/H2t4ObUhG6Vjr50vta+b7cNHv0RAiLcb5MU0
ZzzGFoyS3B6j36XU4ndCE/jeFlXQ/7WaxUNRSe6G+U4PO7AkW0iBXdUzKu6r
ugpyturrR53KPSpZKNvjhHsQz3VMZQ6VNKtyjmeTgEQMtV+KUdYjIxR14AZo
8vtLrHhJuJEFzBedVq39UPVjbO7j3ecUPKVdxx+8j5m1dpALNaL/Ev6cmKuJ
CbrlBShQt16uK0Tu/NjbNwg9/D20vtPUWvgo8LZJjc+N3Qk+0bb48lhYATRG
qDMQr4ZhdvvXpHkONvUHsrI5A8mVdnz+eriJjw2tUfMc4Ss8pJGY9zDBACmv
Gh6m1rsog8U3xqxlKdlFQ6BCTeeGQ5vnWtuTrdSESHXVntgJVy2YYXiYvvsv
nUCDmVMifdNPPeG4eW3PoVbQ5QSYji1+3q2t1Mz8aXYyDQCnnmvTUCKoMJP/
dYFrIZ/CGyCsr+3RXeDSn+DYTMbqSseOHrc3XiIInSM6Htx+S5b7akqBgZOp
KNKu8ZvtK5pxp3/j2hksrDCM7q92pRvLQX1rCO/mfFcExJKMI0/iXHwArg+E
3smENbqhvRHe9MlsMBO8meaDdG0qNKKIFRTwhtWK4TCHbnVHaA9yUADW/pSK
lUMScjDc6K775rn5nnfG6povwbNbWfXD6ULyhy1I/bs6JCqr/0m8xggfm/ws
225vQCkMsluRjaA4evnydYBYISMslHY99RUydTd12csyzLf2TuuwinkRqXUW
pOcFXpSIJdn472BskRbXY0HqhZ92MhTC3d3ZKaJYJ4HQyzidU16iwbpfU7ko
NJPLdEnBcWV1qRz8Sl0eAJrCi8tU2w9La62TRoIA4BrZywGCr4TQO1hpU7CP
a6G18n2Vx4vDjhFLlKPCtl4qdrOAI7za0dfSeeds3++LS3FMTdqNGao5F/Y6
gAwEta+myYzT9laeG0ufMqWWDsRGYkUvdP5WXEAB4CWUO8fNk1qawAwJ5Niq
e6p4D2G+gS4mQ/5enMJ10e1O7Y3aGvE+7ykhSeB1Vrr4FjhDBXfH8MOyoNq/
I95netp3UX7E6+RByR7QEqcJVSuV7XV5umYLgOd2F0OKtT5Ybdrft94irb2z
IfaLq32tUYg/buGFZnqtpl/HR25xpyt9LjQ2OoVHQl5xJ/xzKnoJ+0c18Cda
VMcXCV0q16XHPfIX8vTVpyrPm+eBoJ0TV3iKQdjCV37I0X2K/e5EfDplg0v7
NGk0uBqjNbVY0jc/mlMT6IxDLPB28m9QQ0j+gEXzRmTdUyYqjR0nFgI3BIsV
wfA+rZ/xsgMygTbDoRJom1PP3DQZ+7gXKZrKIKb6qCY4x+uZK7/FgwlqVkNp
3vBkAhKL3tBv9SbMIDk20/A8b3jDzXdxzoL3UejwKjBlzfzezCZ9A9eUdxgi
Kks4dYXkuiGzRMb2MAF0g5XbRRnEUmu+ovVCNprpbabO1g2blIcFfNQVPB2J
1AfnchJ5LfNa9ysrJYFy2g1BGSy3RurWjeuwh7HaTPtBBgKrUaXaF4mkmcXI
Sugh4PtJsUea/rUeA9sN4UOZI01/5QeG2GMXbPEggm+efPdiTBldY8+HSO68
+eurGJZD+udUbrbl92qmg+rKipbib+DQ19Xbphaclkd9O9eg4CEqPTAo1gUj
0xtTMjYlWucnLyTJRXTNl2aPOX14gR4+L985ySjsnYkOlmomCds1rf4Bo4+2
XqlS1GiWZns6IwzeSGyrmUbzrFh9WTH/iBc5lFrkrYI3A+vvkHjGr9vBIxu6
j0s0EayIfPTjnYB2pHsCILTwJaQ9rXQYdvqvVv9GWREoBZ0P0PvGO7QmF3K2
Ocv65VnRCrQ74nduaHAMqJI2TakaSUYyM28C/hUgv1CBOkXCiF7Aufygp0QF
p3pygU9NV5BEwr4rUFLl9c/NSSwNwEm9VzvnunVX1J810uzzUEauhjN5+BWD
9LolG1+rHTQGaves/VDhf60M1pq+w4PLEbO6d5qi9gr9u503W7cw0oF0cXyy
8YKlRMfiLwyXge/yEkljT/CoVD/Ahi8AdqwStvdgRPR5/0abezrjugkj9iUj
1DJV0fGKVkUHicRhJ+WuZqkYLecvixxfiddS9CvLov52X3HOXNvWvNmg62Yg
P6pr1K4NUPcYlXN6lui98FITaNWyiETuoAjfI4UUFFnsqTUjcyNv7fobC+7K
ECaY6B7xvgmf4m1e/BPXVhEBF9WvM3WiIXpgvlfxPPXvelmS8im9Wmqhkebf
Yn52wlQvbKgufhtScmye1xFn/93P4cgTuQjYnU3dboMc7l45Z4wFjbk3BiPN
X+bNmKiLld/3sL+JRsT1sRIlCoARQLNBiw3CrwhH+N35oOjmmpfTuoeZzjUI
26nHrPK23k2Ag409buZm1SQianAo53/NpGtys7VAoTCSA+wMnU7GwUCbyBho
Z5t5L63D8CCfaoR948RB4+YNqXu5QPiiUdYldnOcNtvBaI8VHu57z/ZdyqDJ
Pjp3yuEw4neCZ9kKXCnfMMLi2l23PEYoX8S5V10+Di4QIgH9R3NBWb6ZMZkO
7TK1UjLur5lSLW4ISvbqgqR1YlAjQD9YHFqCIHnbSRStPIClUAg9svKK3o26
emwCqz4e+Vo2L15Rvunkhdskk964Q40c4CFPXKja9Zxmb6OMUeTriucVY1eg
R5r5xh5y9nAgM63+7dm1BDnD0rsshsLJ6f0pszuWlEM+iH9g0DAI8wYdGM2P
l71quFPo5aIJ56ocbvOdw5F6EQFjiMWerO+JtpBLmYwIMQ5+HbLclAAo0n/z
JmbZiSUsSOrfQs/i8o/CwZon7UUVtgCUr42sRbCLr4A6my8J0kw2tVn10Yjf
LGx8TJ+HKBrDZvk3WmxdDtDZjieVW9IpUrQDfmq49lwpzxjE7w4f3K8Vjoks
ebbDtT8fT3QBaNkPc8o0CXwg9HDlX/XXaT/IpXyDBJuBK5na5I5cZuDb6Zf7
Buv6ZaVaIJ7Pe1Y58/+c/Drlod7piys29NOohaopfK4R+7hECSktubEVrR68
z0S+HAvv8NeY+gxpKE4veRVZCzDS5Z6/lqs0Ri1pvHxnSyjLVquXnVVExKxk
jimPh5VRX/UHt+fJ5Ri4VlLwIOF0R5zOL2EaZfTwx8EhkjmwK/f5s+02rUmh
NFN3cimznklzNXOw1Apps7NMMlPEtQB3A6GQHAfvVKE91YwBTPHI6EsewD6f
EOv6ORNYS2G+RUksEJVyjIO0pDnBr2Mwfp49hFyH1vRFCTK+cU1fO4WpPiA0
KXp9Nmdz+G6HZdnaILN7ri5II1fmMAbzy5Mr7V+IT1YtoWVX5f5przTZWX2d
EoC9n+13C8puj2HScxKhGAckg6GriCfdSQYHyLwdmEAgKJCkSsGVGuGP/p68
hQ+j7UIshI1UFGByAwaHrRGJbykqY19+2biBo6g+UPV+Pt1DPgq5LF9gV/bY
o1V5ZFv4d9vMpu4fgEvm06E+mgkEjtdWxngtWYNs6QkpTCrichYDgMO/eEuv
kcuuU4Iq1FIvf6ucim4nZx+/KeZcj5jjS17c5PXST7ARqpCDobCpWec24kVI
kx2uY0ev7EpHQZ/uPOwdgF2dawkzjdGA5WiLyVY4M6di5gW93b/rkt+JyK4V
asFa/sPGvP0UxNdk8JRG2dpnJOj4m1JCkJFZma1NhY1Cg/w8AN9PpOSdsQoJ
z5SqTs5qiISVHwVTk1tEcwVieg+IV3m93cPuxuf3K5pb5ibcbCIhWi4C2Lny
zIT52Pcu4L+4utHl8bCkI9ImfvoaO2ItQZCSmt4FJr9QHEv+8rFBA0/aLC+e
Qo/x6Ng4c/yNJuUS6ahMYsNhBo8dDPNwzhuVfs5CWNG+HLOKLCvf6UHgb1PY
Vy5N9llkS/eur+J9uVDGEyE1whMOa2EeYJ01sXYDxG7OF0PBYOnSNe43DS1H
kqB6Sn4qyhcavoVbaJr/xQWiKbNQyHYO+tNyWVFr7Tw+xjPyspE5mm9Px4Oe
/yb0Ib2GGQ3buSvEkVBDo+9LgAadNs2/vTzM8js5psEhxT/HuaYqEI5Py3Aw
YF98oX1C6Pv8gahKS+dcUYwEADqMchhHf04fQpfHMqoGPfaYcfyZCgSgCkMr
HeHvXkPqsbOOe59XzVuEdOSf2YNv8/yVc+D56GI71OQSJPbJpA89JbHSmsOs
SGrvtWyTs6YHHrbyWWqTbH7Om4BuDPq4UFt2GwjH7W9WssJwftfCzL4p/kSu
roDByGoyYEnC2RGFeWmGLbbSDjsl+cAPLceppzB0bqIgQd4DyOuX8QOKXS/m
nUkIXq+EKYNjlFAY2JcQf2glj2AoJle+QpSJrV+bjhc7w4sxqI1iATzQ0YDN
eDdRZugMQnsf2s24ukiM3kYdjxjboKIIucdk097crL9+Vrc4ISQ/rlNzZD+M
rTHC3n5Zyl7X81Vmrb9e/EftUIzX2kRkT2119BRKjec7WCBmae0CZbJ6AhAt
3NO1LL81S1lYozZ+aIRIcHXiBYR15Z9xWu6QUS/14Yqrigjz+pUunna/WxMP
zBZmf3b+4wtEBlXOMcEaKHzjcSUAaFaqDhGSkI8jRPpSVG+SnmGTu+lNc0jD
vcxv/UJP9abrgjj8akbM8FVJXd0ZrQdVF4Beu6AdTV79YfI+nYRzGwP0Sg6x
sruVRK/JwgGayfZZ0y/Rs350NSrEqCR8UhlXmLJ4ucP0abMUwxa2ZD0+X3Qh
LzE9TW0HWT2e6tNNqt1IvAsCRe5SVJwLMW/mqGa6SHiPM9ci2+0pm9mb45YE
I1kHbOAU0lJpu31Ole6vCHrv1FXfO47v+JLSVpVP6eyWcuwX7kTgZOPG8q9R
Jf7KCg/5GBf0XfjSWXbhvtziXdZ0rK9Uh3+GYzP6Erj1fXRzu+dl5OGMn9WW
apctanBpDI/Op/thh4U7Qh9ZtrjnJ6WW+SUghvJ8EzkCX950eHjew8ycucWt
0mA/wBjvYfznm8Sf+Jhlzj1NPqso6inMjwgbF9mtqkVpBcmMwQYyH+/+Ww0u
c92pQ+xfuDus1IC8i9gDNQYKg6FMgsYosg+pVlK+/M5hqHAl5e+jusM/1Wf0
+ID0j2lVmt+YEZwIlGKhntPmPOcWwo5lmCmN2sFBkM6ojZO5KZ4N5MiDz+Fk
6rx7/eFDCMZ57MI75ykc9a8wyL2oFFFEhdNLeNB8F1AiEXVDh3cI6jiGL0lu
04w2B6E3rU1I1m3zkHfQeZF3y3JctkLLf3UBurvzXasaXSEMtOPKgnqbDR85
uFo9sYBMNRkj7wIwZzp67vG9rIIhlTgfYAt5eV2peUBUfD91VV1nFLiX/S5w
fp7lKG6wTu02LeRYAoMoDYah6GvkwjgxAL7+rUmMF8ihdVJgn0VSyBuz15DK
qM7CUMpZwJ2031+oRaUw4SS43OOcbjXo5UHMm3+6zIpd9ay3BZWwUPIblk2S
0VAcneaGkaTsW6zBB10BchHzHT4UsH86ogn6ewyx41nepILJeNeMtapVv3s0
pF8mnz2FxLJsi1wlNdyqUS24gu1PEjrZhYMEycwl9iwCEpfsLR/Y2moVOkfE
1WFmV6opA9Nt247jNe+r4n3kRlpozYxGSs8Wa2rjBwArFKxPcY+OGpA45DdG
RSYa4min9DEaWCLi2nxCWzbUXje0hbhDfyYTaW4+Ri9uK5Q6XrcvCuWtt98E
7Lth7Efa/jkywxhSW4c4f3ybrXN5Z2udMY8YV9+TrvTyrEF0k8PFzP4oFVPK
CSQpopj21wZqQFShOEhsWOpipAwPrKDC+Ab8R2eajNuU0FO1eCvzAnELnDvX
BEAuC5pHLh0ivHdiruJ0wxYt1KB5cqfEAO8jCHUwPK2bwmiMmw4ALRvBh8m+
Q4yQEgzYVMFWh9PCrD7K/lrt6RurjVSSh6btSaiuzjc+K3WPSproRKzRd/s+
Jcm328du5Lx3xys0wBJ2FjSIIu2qaRUMOjfwo9shKrWijZAY2NjMtfG0JHZT
Nei8S4a3GJQ8AENEFR3h35obePDyddztlx0Zm3F580PpzuLBNyMI8gwOpi5E
StH2jWdKa9gjUWQvtGcMlaf6mC2q4W8ds4GfxAPiRR19wXr67hgeydXWE2/w
zqubkpHMzxGmwa5/iJhFYfHgmnUi5D61jwohz9DsFVqYWQhxxqgg4wQHGxcz
y7QTBRlNdPOzxHiw8pgC5jxq4YB3dQLi9BcI/FWLAfYctiAB7JY8nLdLENmx
3A6/geFBxu2NMMFG0Fh7YatEQqOCdvnNMg4JQuniVGyHWIAmA2jDNoU+71Kh
k6yZ7LjHtQuWzVZxd99e9sDvB5PGZiaukLFaFw+qBbuZO/uEkMg2/+Ca8ZDr
X1ACm8JCF6iJFF9OdY3iCNhwvRaoLfLT0R8AJgWPGXWvISZ8sbLXz6E5qrAq
V6gypTbzU4T/cyGrxghdJxJW5Ftvh6Zt/t6mujRwjgkyli9vuVRqiVMCJgfh
AJXWgCA03+eCA3LAZrCF42e8oGrtAE+HcozqzGpfyXkwoCCmdv4/3yx/rxtw
sNmUZfetGmytGZGq103XpytsaUACpRFt7Ja8i2euKDYf03/LuqeanEUERWK2
JWjHQPVeAINEUstqGog9bHbdROrCO36rgWkWdX9G25/yVrnLWpL4FMdxBTLz
wwszihhpTcLEVsLWWBM24/6eZDhuUB2VvldmUzUUM/5zYigo1hezxlBwcLjq
jpGNbXTvVp2L5h2xGYAII1pKgpGakmlyD/HdjNTzqvnEaYupEOs1pSQSvpYx
9vwo4I8jovdWvZ0IoDyF43/E14z1z70hjJAwmJdG5iohbyZDnOAyaiZMbW4N
5pjovQ6h+6HcSHYzncZBv/nnTQ8JxhUcfCL+mBGfkUD4bFtWrjvSWj4VkTiE
Ie+mlaRmeddg0dcHmlgR9lKXisIH4KmwMXSQO/US/LOSRRYVYt87JpPcDGmd
pJd0lDhEW4x1sAF2l8ARBJRLwTrAf2HlgIZ+Lvm91je9dQ+JfhHsKFARWruH
QD+scyVjTF2I77XuOKBiYqTBbXaB88GN2GBVjZNM/VWQXc5E+G5ZtGqc5ctX
W9Bzua9vva5CprijZ0aLQ5V5Wa6ZqRlTpDvKsM6ip/kGCkTHu8lHqt9SRGkL
YTxXI8crYJLsEKYKqPoc+g4NqrCI7tzxR9d1a7GgelV29TIoPZ+12xuX2AfS
vH5jGqI0aPWO8T2OCy+VxXMSQnmtbrwjRCLLfICrPb+TRJctkt+wAGINWbTq
yGEB8uCaybfyVvcyKd6kjx0FEXpCM3vq2GSvSqibbQroGDDOZWTzD7/cXjTZ
4XTj/031gn59j/RYyP61i27x+H2i0yx2ODT5U0XmCC7ougVN1Irtsr+HAgR4
5GaKU0mv7LvK5FQIKoeVyX+1llslCAuOvunhWwdUWPXHpoJzaxtd3TIzAwzQ
TfUIJe6RSomL/Pe7wb78tZmdrzQYjBDJdECgXmTc5YDF+Qd5V+VvJ4190SrZ
KGuQDGgCzZ5FpfM4JPYuXXbdHHTmC56qWYFXuPtVl75YBo7F2xgKEBXhqitO
hEtQ/ZWhufCF1QJoJ6EtdyLMnd4DYPjnB7pBRiZB/aeLH39z54++OY+BSCz6
y1ewohwZahysYqQ/8Ns10ZNMJ3hRMTV2CrN8gLP+WjB+4sjZ1ETAP5sgT8kV
aRKW978j0B+cRaBX5OUpfqQ8fx5MDYztRhFKZMP396hbaBkY5LPjxkxN+9ad
5UcVRcWHs4RH6WAscTjavWTSnJeA+vHHUrdmC9G+Eu+jDOAIb8zk3i7j3I+l
YkwkGa0P3Mea7hV3r8a4NKZGq4nEOuKe+7GmBIUDVnDvPTMFkmzW5BJEu6BU
Gqg0E9kUz2KRJ1Oy40eoca95EAhz7Ad90/XspLdvnZrvLh73fE3hUSmvOVxO
C86QNRXuis1SmzUFzyuwN1NHs/OmCKxnL6eQPFUBwFMYWHWU4XK92P9jDtJR
DQZ1aCsqaUWyO0yrL0rSdZbkpBLN3VIBdNdpPNFK9xZ6evUYOdqGG5/UMEbe
FBiVDnA8y/ZjpEu4qSbsnxce2bue5PxUhwaxOahnVQIR+/26mZvsBHvdPLtF
VN9ErgHOIJDfvsRmZK7yiguUBheBD5zzVYsQvlioYNjeqH8f2cDOnpBIzgeM
Nx71donvNEYYJfY1pnDhWWKO9aTlnfF8pqjep2cetgwdueA1N5FEHNd19T7M
k7NDriFGOrDpmmXO7TZTmZropxJdAquPL4LIV+M748Dxw9NLy5tI/Rsma7sy
T846aXTUKYlVmTBVZkXFj30lMAAwefoF8AYNfJ9+EWnwR6ZWE+RSO8ImCdAu
j8U2P36cKpL3ObFe+AvfW+jTl+cqhMsD0lms20zU5BQbNBUY58Z0Kd9c7wfI
y786I/FYbv5L5Fy84Cq7iBeovxPe5qv+mtmdNliInBsPrNv7liFeSwfBz/1/
oQ+JDjjd3+FJ29metHD3Im26unGPFAypDrztoX2xgG/bF1HzySLnEfNV8m87
6jNxRJn4/HiSXfFo787Zr3e1SgbVOsDG8lOFQJkdE57Wuk/CQgjRb/6q9cB5
lornMMW48ZgqXpOUOPvFZl9fvNu/1Xd4sCou4HwJlP16zkxmVvGvHMPmLgeq
oSrLIhs8DyhWELMSBSp4FYvIbrJpZXzvei9ycFRYDLpLeVkmTZs9EGdtCUHi
XfzqW4hEaQWhz9YZs0MDF8rj9y5rjO24XTjFSM5fuNl3vX4dtuw+mWlYUXXG
FoFCm2e2l/pA0fIehEn1mKAMXXCd1y/6BjCHYLSA4OlPdyL/MA8sx/xwVSvZ
E1Aa828qxk+dhyLkAHOAjy6f/CHxBYuNr7TmwvWD7pmzlgrjeBBnJwhooMEM
JGGlldUon0xnOsNbXdYAEtDH3F6F5MiH3KcriroobdruGwRCdLfSpEHi6HwO
WmRO7THGgcHtV+Y2OOJsFz6eqCFR4lPnMs9YU29XKBTFAEIkSoMFoRPeRQq2
1zVErRU6tHlXzmBGxiObfoJgNJ4s0oayeIiodz3m8AQgtdMs1b0X+mEcIuyv
PNqbvtO9Jhpir/ydFfKs9wsVH+qfU/KoOfWYVqffIeqC4kWu/v9Cil2PJRzF
Wvv/W0lsVBnVgL2ozlUD8GOqjoZzwp6kR2PwqGlsdseENNg9QIOluuNfsg+M
lxwdN5U2jG/ojrMBWIp2jdNDQRWXsm+2kHYIF0Cl3h9A9vcfvtyUVKgdOaGR
MsOUp2x59q+RuE44+03VQ05vW/Lx9qiS2/vC+Ok5TNKzlxdOxk4OfjJtl55W
Z/YjbTPcbgaSSFnHGp+/JS9UhJU2QaUqJG1V26zU2nJzVF5TXTnlv22A6rJL
rgzqwyzJtIw9WeLKFr8IldoohVQy+aUHqoqjna87R6Td0z7yodurbLQIaTZI
RK+CeMrRFBI45CqQMWvTmpJnyjxrc/mcQTQZct4xN7oKI+gRQjzQwamHi1ev
qyQ96qdNBLRV3WrZjdze1xQO8I4zAulaUeSjMQtk0jYl1aeJymtg2FKx0/f6
Y8c+R+q7kH1niVsezq2eRo0af9LvXjHI94ALBVzINsUKIGiZMDoX4d0ZN2qe
Ri8CBa8HmE5j10JBptChrkK6Nqy0IKfS72Nm+53qdUopc4Qb715RguGK7vcL
B0IXdL2OtJJSzLV+VRrkqkjbU+ROb3Me1JY/CGymdffYeGEIdIDebsTSZss7
nMG01d3lo7QOTlVTxa5nNd+I3yfUfiEoyv1tRAo1gp2mHijvO3WRmprca38K
XfnLKATsiDYJ+oHvvDW3x4hpaRhu55AIl4NLTAMRExaXy7Ho1wqTJFikzYyt
y/oapuLBhM6LfFQSdpgJ9MYkNpLcRWmFCVvuGdmmAl8XNKfCZUsE6Z4mSs77
NN+POHpul64HbG+beXYMNx2LAj+YCVHMSMscPFcLKyxOj9iPzFTQv2A7HNIf
Ss42j2DPFYW7B3fK6UkvZjqeV2sC0ihFo/dKKfUVd24Vi5EqU4bCUuOQNtVp
nTfgPiE9CRfY4hZP44pmk4Jux2AuE7fLfs/9y/zlgXW4IkNpuxMDZWBtzGur
gc5xukTqDiTGS5tNrn1QrpDVBKpEkXQQADDTN+5r6k2JF/f1YqmEEFSZ5xXm
CH/7O96DjxdKt9oHiz0uHal2Gumj1Tec1MWm/CoKVg6Q2iCWwSX1z2LaRsUm
xl/HM23lhcOxWcgF8YHqRFU2ogpsO/s8xxtPoIK3fDZXO1Ky9z2lrJY2S515
/mgTBQHbrXuvFWmF5hW1L26skGw++p9DEmianf/ZzDqY5bh2Pl4R0kIg7RSW
6v4UV8Jk7pyWx7eWopZTJQyNC13ZB7m09cvo0y2GW5z/Qta/e5c/7ECZx8kZ
HIGEfZuzb0QJcOmwD3lohSFT9FFoCtC7NZbYcop0NEZbgD2QHXK7B2bFhjw1
Px2KKwp4m5lSgJLOAniZeKPg9S8ykAdbYmYDqPTt7O1V3eFcpo5xJZMqQsFx
l4KIbyNfC+2+W7rKZa8UXoY2UQr8YRNRW2WunluuSuFK/GOiV8FmF3qT89AW
xMnogEt5Hgf3JQzf40vcPdR3flWU1UwXo+Ftdt04OcLeCO6td03kMo7zFjlJ
agR6NUC0w6OpMTohqiRkSw2/y4RbBqaT+deGrU8CnjyliHuOFCrcC8hioB5v
aPwt/h0ZypxqwmY1sUyKyGqiMxZsSLxT/tCKswHPGqOVPYeeFCQLQhZwnGg7
zpA9WwSi+MwrPsagygw/B0bsr2Lu1VnFU6LV6IDIiIdS02bPQ4H30gRWKyWp
nO+37lZvTWjt6hfYXM5+B59GcXGfU0A/ljbooL+usomnOW6KJx7QbJkevb5m
lcduyK4CwK8kwyFjNWH1TsNm4efaBQfovwn7MGE/RrFR++nt3xFNenIE3gnY
CObd7QzPNrU5ioQbjnD32M34hMWPRToQ/oMhsPOUOzhvYIAyAZJzDOId/W3n
uoW2f2jRvpbl63j3qeI643A5JTF8sOvEPzb7o7qRJ2NHQoIm+RMtgB8MqIGl
BB9QrvzbiS59GdSVR+YdyoaJaDavx5F8lskAlX110EIsVJlhGmRze2ys2B/R
dgXZGYnEAcxUHOlU54+wlYKR4C2G/rXOpbf5aI8by2Ol2Bwl7ubdxYS5/oe7
YX+JAygrAtToJZRNOBZw33B/jhN0VT3/9quRfhC5KUz+QmjSnrS/wFa/QGJG
Vj5gUmTLp/DYrdX0UZY4/2JJpVEd8dtlih1CU6TjGVuolTNp6rRCZQgTsLpM
9D0WGdweCaTJm6vVAVNGTcFTdSYEr9fUgwcn9nVUBqkWIALLMVbvdJUD7smd
x0cRGQk/IGrGfnx6nsTjEe5F9vLf4n13bf7Lk5r2wtY1vwtwbWBS30v7b171
isLbinx3VcoCWmQMCUvjUB/RvWsC6daXs/FnJGwtjn9zNgtZiIp7yMvb0+iU
DYt6HxzOBHi4rdc5yV2K1rQtfj/ebJW8ah8D047TPR6WzkiYjKW/DDnLZr1X
GPRGmFW+Sd6W4MQ2G0pfMn0njdtLkVCaHrMTHUbwmI5HXtiIYIY2fz373sei
csaZwKJG4+6Leo0l8QypbdsiGcGLxnrqDMMPZRuH6avdGk9E7YJj4cC+Qz+Y
QA7C48BKGZvfleGXcPe4ZWm/1uIdFTcvzH7gVgDHQxmn4amzgMFCg34uR+K1
nzwl1R6/NsZipRoFJJ+waZHq6TfCmE04IJexEw3aIV4v/FiN8EtvOnE+sSZr
vUjDs8VPpBGDOargpGUtcPziUUEb1t6Ucv3qeipXEIk8AnPtGSBHpOj/KwLo
i//1QNG0Pq1y9eYcH0lnsvfvQt8k3HQLUkYifbHKxs139wMbx66uJs3viSdT
5RVL03fb39JKSPBaN6fqkP4bgV+fwp81r307+F6csZ6atH4IOCDCHTRsa187
6icqCewNC0PB6GsDhJjMwUms6MxaGG9sb5pDtILPd0FfahiRXG12olA7V1lw
bj3wXKBuLXI7ZrnNfDMO9jpaPnY1OFl6nsvHo2roVIXpebkhG2d4DsnzoywX
MEowE1Mvr8ftstRqKAFBZ0wQZW0SfpQo8vOskqE2RMfrTK8X7F6W7wTkHLG2
s6GYgAowra/E4qsOMgCjDI8oUKkA0BMgsb1UcGWSRLZ5a9AN+G7aWqjgpz+I
ZJsoPb6Z6ZZDPMweJWteLVKXHaKb8bdKNt7BarP7QU9hM9yF2Ae6f6AlulyJ
YSwmPvtw6YeXvorY3t+M62elBK/xRg153cBJKSmSs4Zf6lE1wVuhkaWOAFSq
hfpq8IyhFk0KJ35AaxCCEqvLpcXrGV24MYdg6OrP/h4hQw2BHPDHa6+ybvAC
7l1crnW8ZB+SedikCkvlSut0SbjPZCBVYpODEXXbjA6KEvE4oSjXnNkJ6loc
llPFB7rSmY8I+q5CDlyCDwh6jfX22PLnVcEn9Wp1VXeDMmQJwmsj3q93iH2u
s2SRgv3ZasO6HOqfLOIAnbzMp136e/W++oOIi/+/B8nwK7K5QkFQQQViUu3L
olN8hxVXNI2oLfb3PnLtW6mh6c29hutJ5aUcGFGLw08vOJHEt239SHvKJLNG
g4nbkGmD6q0wU2O37f+X0qF9SIUrUQHyqSOgCkVbZbPZ07x+sL7wKi4NwG7p
EEnkUlvO/00X4KM+UvyYFn3w5oub8x96pd/DCmc2iAyYagThWDLKEHQsCB+W
7Afm137wNAYFc5ry2PQCaERMucsDPwv7aFn5fW14YC1/eOIa5l84Mdx30Rah
SReidjJEmx/xKgAizR3iRjtwe6pi+EmkYYaUr7+cuI6s4hhyEJNBhtFY7f2M
Wj7kGdsy8OaMYvS8zrAeKHYpKo9TejLV6k6ehnowHF1pbCTxeYCJhS4J1pXN
Du5cDAS6p0vck9ZknGNhx1jiOtoVVWCXDuc8vmoymQpR5QZTcFZVlUfnBLz3
tOwqDH54C60HCM4WBAZFTHN8gc6Oyn83wDNdhPDEtFBh+5gdSi4zwU8S7QfU
vGA/7+J2IFnSy4pzV8CmbvMqQhLrFURhCKpeZ5VXNgt1teGtoTqzwutSv5CA
4r12Erop68vHOe4dxm/gbeMtU5Wp6V/BjRAAmk79jXg0QspAVFp0iUKMReb4
heUHbeDpRTiPDefMqwspJkui7VGalckS21icDkrPEeejwK3VswyJrmuGI4he
5scAUIGlThtfsso9TvA7QQ+AK67R7Nvl0b/2s28q+UFelX9SXJB415FPsNNl
R9jNbWYCVNnUFDFPq0yDjidxeKGjswPefLxUHcoHZm+vQ19QbjQvY02z6SY0
6o3AFlfB8ao1rUREqOGyUV6DohKJJtjNKPzylJzhKwqMS6LbdFE5j/y9pglj
PGtaAy70SDKcB1j6HkAl09n28eNJpDBAnayDuvZK4qHm0UfpyRgZafUYgBzc
8QQsnJXs7fTuyca7inY8YOQVsGQCBCvskTn7ks4jmocLgQXaPcQsoHYMmqaV
8ObIOjWOBgUWo/nFdwJiTbUmrYeMMtShtJkHvn4Uoi2uQcEnz+NppgpeZALw
uMohRbXkH4kyAz0qFrzPBuchqnqzMy5Jj2p5K1k/AUdBYD1zqhLp6USrRAqI
4NQF/m9bhD7f2WgD9pUbyh4+eVzRvqZWf5jG3kN3W2DPbMlR+PjBhelDnBe/
E5YcehGm1W7vAUR+XVulcTgfBOvV0zSI4gdr5l+olx/1ZCjxz4RO6/srHEjm
Pp+iQfCbGfXMkNu+0gzlxNNHuDDk5yWxv6cKW/hidsff/Eue95EY+yoLeUVr
utaJ4Iqd4esSH/pvC+GN0RKAOMFWte85swgFICRYaQkPhD/1+3jM/2F+1H5r
jgHWI8y4gO0BiVQQQ1mRYRXgzbQX1H8ouwKGAgTPLrBS20TtFnPnnc+WhwlD
6DFbbf0m7hqw9chQDfw0H6ydrFx3Vz+vDPQkyXUFO9QN/Cx4OIk9rpBAKXal
d7IM4pc4j3HXM3f2LhMRHRfEBOmokCNKyju9gJfcBIsrPh/FZ5fwI4H9Dj3W
0l5/+dQkAIGGNg+jTRSALayX7Ppvb5lAdZVHHYoQiRjCysJTgY+qHrxFqQfG
hbPt3dy9qKzHcyqjCMh0lQoVkSl8fxy1eUiPENl+txgP7C2ANXAP2Np9/y+D
phhiYKo+kvKa1A5QN7goNqFsn85JmB+MHU4SWV6FMp92pvIiIItBAVRzAPZJ
mBds7pjd2Oj6Rf90E6n9+F3T1dplp8FUqrppeyQBEx/HopTVAMkHnn4vovrM
UDDLwUrE9vZTFgLkl5MOODxoM+R7YsMLRgA1qZ9RRJWndHaXlazdVF2NXaG4
z9Cm7rKFMuJnUFTaOawB1/nkb76u6psjfMEz/4nRVRV++WIWyabESShhsjo0
mSsCt/R4CMRZpiZfDKmSD2R2s4L/aVkOrdWB+hd7ZpsLDP3xde8pQDsPf9Bx
ya49N62SHM/OgHYpLStu6CBy9wKrXzTjfBVef8dhTQ5SzRbMWNwdRyRvTxYO
buQc/J5+0NiuS4q93m6BIAOwpUI+ALz5KoTtbb2LcDvu9SCFb2tFGmYRj7+4
stRLZ19BDMpyPXhTH2/5Vg6gRhmGQ6Q8qrHJljzLQEPhZzFSY4dEhMZx60uM
KlshDiS1vb7HvBD9TqrSJfN99IZnJSv9Oqw5EYm4exoJBpQF1FbWDgv+ElcX
tBOi1dL2E9nBq1I84TcTe7gS6ppcb8Ofzec8vw6evtNXsO1MzqvT1/NmxsPO
yWD7dR26pXR6Wg8Zc/OZtnLk3Uu+miu0JprbqWnKw+fEy0uIGr3pxLaqaNSI
r7FtRlIT2m19E9LhWK0QtVNfwup7hfil6cMNoYm6VgiPmH/bii3ZC6/H5/Fc
VDcT99xxmhUYlw0zzjGI7nBf989VVetz/qlGdIHd0qVtmaffyGlcBdbzRAdD
hCLpK7FNmRYd1AmmGSzuNaFakDcqWI4d2W3Jnjic/+eUhaiAA9jo5AbXZgA7
eAKNBB/+Hsy/acxD2xhXvNYbc6PeFJuaYS9RndLi9wNETwdkYoVgp7MQZ1s4
OX0r0toPisR5ts0Pr37ltcNLkERNjmzDJKz+o3lwFqqiOk3zY+8jzWsXeLoj
gG01aU1vHBiC8fHexsQhVq3e0N5RdUC0PwAc4LDkhpLGYCp6zlrwpIDXIYN7
1J95JeeXMBOXDKhvazdK0wileflTW/Yl4zLGaFzWpor8OATN/sWPWZhhWmAZ
2i1L+PH3VyBR7psRT6dgC3yCEBJpiqYFZMaLbzdQ+jbW9KsqY63ngS15hAWU
CxolTKWpfAbx42cQ3vlCLq5RmOG6Sq+0m0AwJlLNqOtQJ/P9zBBJIfHTJvD9
q2LFeCihl4+tigtpO5s4wzj02dHYzWZAgK2eT99RnKeMtuQKfcGL4z1lbPVR
/9IKY2RS/sC2sYfrOdKw05RDEuq+jtIZTPCU2ReOtN07zxbo8Lg9R30Vyd68
8mS5r2VRM92vgKicph2LDYtnX+PIxyrpgHt681w66EteNgergO7PMdYvAFyd
hu/8s77kBkM6kThkTlQoLWWFE0YVMrGhAMB3lHJ9tGOu70NvUUjtl7nSginU
WJm/bwzSoep0tw83yELvbOlJgNCZ/Oc8VpxVdfKGftxdjQYBuJ0IKhx4Qnlc
ug0RawW1+Z4zvRJ2VpewJb1UnJp5bxsLbmQAqkY1/0n+MLYSIebi7sPIlEKS
KJfyhoe34t4sOa9F6lAvKqMQHhWhlFRh6Kg8Gh1FfnC5Jt0uLkSLam2S6pcB
/eP6nMgMDmH53zE/Kh7jE045WrMtLV1YDs0fA8jGR4KBGmNQE3h+yiq+d5UK
iJNCY3KLuD5jgxFvFFaDIhJjs6BzkprsUPSA2600VE4LR+7eQUBmAu/2PUHM
tr8t2/e9wEf6Sb2akuHBvbYW9ry3LdSnXu28S41YMAF0ee3kdfTluXVvY6D/
5KsIZWJb+m3ME74mkvhZW8FrKaBXXOEPmc6od1/JgCl5ULAIO78D8powKPjb
sq9nY/ea8p+y0v/rbq0eVOegmcQ/L2PqFOiJcBKWGALAd7FS+PDAyYv4n4BS
XQQSR0bBzfqzRrnY6MZR+AY6mypdqg/Jx2tQj4U6WX5al2bJbVjvYiSZcqCX
PEdXrUS/A6dXMe4exlPS5kZEH8qbbHcTGorEXPsa40H4OJAXySafLAdxSO6r
mSHI8s2d1XJk4a2+3tLz+4wuLFmSMp1TdZAIReKBtOLab2XGxsfDe2PaY9ot
OlyvHDTpi9XnlU+ghgMyUkVeMpN9YPpm33XngLmp0Bvs3dpQr2cK8HGi9mSi
/Rwh9c2j592JkOp1+tssz1T2LqenG5ls/1VS/iHYVgb5S+UmqtkkdCdb//9z
y2wwqmPEUm7VEgFolh/6iSg0Y5IY8A34E84Ec/rwrQRQ6mb8iTg9BfpwGDN9
ux24ELHMVAoFSLFl0DaiWOxTow1XaCpLjcx1rgix9c8ScPkeeQlv4ETr5q2Q
GHoOTY5Z2fwuYBaf4Z4TlkM5DVO9br4CcwvA688ILcPZ71EIx9Bzwk3HesTo
mlq7myjCZhf6CWu5RynGFIIps47WCfuEWojuw4RxkyNVVJLmw+/7iwU+vBYn
lV1ZcmHoxJK0XDBTg3DUcYbF+Z+Y+YHTnyzFtIfYDeeio3NoTmZVYMWculho
YSF3/7u4eDweIGKHpBBbrtoDTP+xQeJbBrzMg8eYBsHkserNlJ18AsLARfTT
rhwXsBPiB2ew8qVHIFViq6QVt+fS7OxMBSWTwf6IL05GH/X+gAw2+sVg6qWj
joXujKHDTS6aqV9XKrpJxpLtPitqyToEQ9eol8hWML4X/HzJTQUbUlM5+kAV
z8fABk4JJjKF4yRSMKMfuySFZYZ6KlP3+kd5U+LuV958afZyngyIFvprB0sf
R2RoWkFwBegUBjf0KherGaNt/4PPgaNEpF2duM68bteKcSHxhrAsQ5EYI8Q4
qaa0S/es3p9uYTFHgSdp32fu0crPJNg61no7a9nRvgmHJzh644f4IK1BgIFl
sMKSIxwElHgkQBthxwolu2JMEE6bS6V8oEO0yU7n1dRq0YXVQPZYjryy+Kx6
Cl/M8GuiLHue/VkyWAVXC79DWDwZxh5cxFiEWYk4bnWpGyPd3ThHlbrnAcld
9Y6PCZZwx01yxkhgdKaekuFL7mQ+UPsIerP0bmyoAOolCF6A8xvjR07ZhmH8
vsIATu+mW2gy2nh4zeuBd6lz9Fl+bHFP96qT7A1jctLG6uIrK5ndoEYg11AP
6i3uAGeoZK9oct7HyJmt34s4G7q5Csc6tsFT+H4BkWzgQrAG9z4AhNwX2dRf
798jMYSz0Nm3raxbmHJYybRi7JSgiAB0SB4s6F+f1Uzs+cxXIk5lBFeYsBSi
9gUVhe9XgFuNH9wP25rrG1dgSevOhFIpZYvcExYIH3X3hy6c9SjPuCR0TvWX
JUrIJCs0hN0ZP7tAiQdIQoqujpzFdIfGvMMElgOUxajGgs0ottor+Ny6JlSW
Rp44XhQw1yy22+E4JEt5JfZp1x0qB5lMJKWpXT3AzoBRxiGAgI518WjTbzBt
olcNpdRTJz/KhatrDXxWmcLfHcKAyVAldTwLseZ2JNBVLwdZK9G+L6yg5E8f
ifCy4PpZiI3n8iBFVdN3dnb9ayN76L6RIf0vUJKsG5Bkiask28fS6aTASaq2
JAigvd9Wl9WAMCzQnG5GqwZWGN3fJ59Z9euhdm5BIW4uvlM1fkxzXBEF2Qiu
WbwMfJZp5TaxUuyUV3eKLzZRF+QI2b0kzM7ebFKghwcbEwGTCPcwsCp8OC55
RcDlj5e9EC6H9PHff9MHMvVH9YuqomfnQ55lSHMQMENf+PqlmWlQm1RkLs9A
VDAxcxkKPxggT2vuhDrdKg6n4l+Ns+GLIYUZiWllrmi8ZrZkqA/wORrTQViC
/GE7hHai7rrXVi6EeGN0BW4V+jp4Yuh+pUl8eYpo0YfIsxe9d7DFnLA+/fme
jSgqP4uPdyBxKWK8pxrjl+dTkEboYUzmBEQEPzad/n74LubVq3qAzMY4QMVp
PNP/TYpPYsr5v7Uct4cozbYBZJzjloHTrIuXacAFteaSaC8f0E1wefu+VYtE
7hx2N99xAAO65YXBBKsAWi/FeYSSCJUXsccH5UL0ZDa18aCVH4bhoDHTauaP
AMuRHNBGA3LLC5XViPbcIXiu9GUGaFAZCT6NpiBwS4AJX790f7gLpLEGoLa3
KLZMh1asbkkSp4axnf140T+G+Yfsfhi61ZGX9qDW1sK3B8KLtr2cChrJ6N4t
SlR5ZnNkJRWnpsUD+8hBI8zSSPBS9Efee4mKC5iHB7s5kegcTSwdG4ouM6V7
DWiGcprzw1Mp6lzIhLf+y7FKaDTpqY/jK9M79nHPizBFcNftZcgU3MyIX5XH
Xzk3u0yu57BBXJsIbx1pTvne49drZP83+6F7EZScla7cMJ6bSQtHwer4loU9
yQvdGA4ROe44NLNp3rz4xyvZWeM5xQ4KvY4DvydHrNJ0S2sTLanwWzwPlEcd
/5ia0Gyjqo87yMyR7eXorZLYRz8T+UcF8tbG1iD0MFdj49LTtzw0WB7MkLUC
jVOrkEzzF53yV8U/NU0Yf/5N6np2MCH0s/92+zvm5TNMbpEd5u6T3mJ6zFLo
KFflE6hQ6NzqGoHcaASNW2i9wN/6519es20M0ppKUsFy4Evsz9JKm8oDUxC9
F9RhjIX1w5qhoA6g0Zgb56YIk3O11+eD6xS64YyOhnBGrdh2QaRjqVt7kWDC
/qPz59xJbqk+0/pHtO2t3Bxg9IWQEE6T4rMERL1mqj1A7bf/biMaYG+Pq3MH
M+kbzBzpmZPjwgmLL9yRnDFFaaJScFG4eh6M+oqV3R41MUXFIEfIx+FSBv74
fIm0B1iQfD78GEDs5x2dGq6LgVPDGMrfJpBdxFHQM4bfOX/2UxOAUvK4K43j
7/oNsDOmBse6Hrh2ejxyQ7eyCydztbJRPV+yNCHh0pMLJ5pKhztFCr49WvYN
ZvV781xtKSaRe6oQVp6gm+Ulc2PlPanVLMFmatviEASsC3POMJSEa4rzpQZq
/IB95fbrz52FId8Lp979xs+JbOiQhaRg8ZtzR9zbfSFEPzv62fGKkC5wuap0
z9OhbhFkj4cAuUciRlHuh+bzwlQqA+6N9wWxB+ak0L8nFfveqSJaFAZg5fSf
1Lu6P0OLqGwN56nRa+ZVgCEBNWoAWb+1FbBma72OAuOJS2Sq8AiZMH5+I5dW
70V7vNcwdAplSB6UBg2PqIQ/GGZRUwHKC3g1IatRUy4sHOJlypAeOusJdFUU
BjXTVaSg6Jtt2sXzpDXO6CCH2nrGLe2UNqlOGMlT0TREtAf2RnXQyNJVhF/r
Y9onaOvjqkKsbRblC/wQ2sWibDrSfOTz1+wbUpWRLlyO9PW+KfFMZoHsYlZU
z6VpmG25U+0LR9B6RUPdcQ5oyFlPipA7WCq5me4dWHLlCYbiUZkrO3fhMLO1
WPfa9FfWUE8ewfJnWZM5CgCoOEFwiJKIe/GAcSVD6M3jUESPMJwuAWwgZO8Z
gG3IcP6l2tSpDyunjRuj01xx7oaKAMYBRsiDcajNKD6tEkDaENalkZdBSXeo
X6k4Ym5i/TSZMO1JNAFFKR5uDKxpbDLddoka+voJaMFn+K5kW70Kl19g66cK
2lYZKSI6na/0R99fdlE+0wQ+RSyUxDPqauB8l0tCSIB4uGz3mVA/SY0J7O9h
7iMCXAJDknRwaejSuQP8d7+1L7V01b0tXzLbjHiDzSAYt48LgKjcoJ5/sTzW
KGQjPfk2+G+rZt6fAV9zs/xRC+Dgx/Tn55PWyiImfzYjazxGJ5YTvDZ5Jc07
rTK8NLanNUlxoHC0cR1Z410RdYVrDSCzlHj/ysnU+Nn9hLRp8Fafw9/INjoJ
9U0riMtaDf+jcqbl9nTeAPpRgw7IrnrFGrbWdtWIUpqlSG3nqEJBYNCWVKSx
4FqepsvzxNA4M3+BIcjQN02SRboY5+fLVW0+T/2VfWTPlekPPfoT2J7Jt/FG
yXybabahrGSmNRm/h/JNlqa2rQTFUp7IGj92PZguAofGYDhdKbtiilxmm9yq
VSt+Z6VHtcI8PPZaXpzj8sfOCzv6fRDLDDHCq1Md8AuFmzPfKIQ4CJ16j/sI
Qkiomma3q9N0i021DhFfAyBB+KpGOlYM5mBvOnO7u4QCTph+aNv9301XFcRS
HKMxXYWzTN9f9iwAkqTtA5k05D3DNB7ttNI+LN89g/WCQmJWrnycy200DRMM
l3MxkJaE6nIIFuuISm5Jy+SmSDuL/jYZt9VQY493JB6JFElVE365iG5QQgwD
aHSX3iiL+JzkuYkUA1Qbs5dtGiCUIO8FpHLqmLmN0GvFD6jcig49T4plmZDa
6mQys8A4Y9WK4E2nu8+yN9an6Cs2B3iQbwnBWMVUBmbqR6fVD1ZfLnE3eYHM
OODGVGupOnhFyvwbuKK841NPbPw6vKQT8Z07wQDmd7dOuQ2b922+1gquBFMd
soMjdsWpUbTWXyH4P33DRFECUgxJK41CQC3EwITfWalbuPU8V7qVrPEKgITN
2G5bou572w07f4IPfZwSbpIkJBq2FTK95pr8jietJ07lkaYM8QWjuQGIPbku
hCLq+Qzd6vrnOwtWfP+yR5s6hMtop5qjm3av2N9D8OTfqmDT0Hjf1+AghMUg
Jidwh4EF6JxxlGTirMQ/RU3SU93ou85io+kOAeiJd3L5lmQ+CqtENjlYjcYj
Q8LmkiXkRrYZeTFyswnz6EXdp+pmt008/KgXkF7qE90Am0qNNC2+uJTiIWfh
gSXVuSO/L6J/HqcSaYjfdb3x0iwbeTtYA4BVnhocOw/WrnRwY4VVy4IH7Eex
L69R1Ra9HSr1uIGTCAKYdjSEYa/AgQwnFDMHYjnRgJ9NZs7AdBbiC9mkx3aq
TIxoYg8uvCF5CeLhBAZM6ttbv2ojBPB5WZE9vIVE5cHwul6NBScV5NWWFatG
NyAMc4GmWH7ZcB68a+SYXdNnJT05qIsZn133zprXLW7Kk22TDjimmry5QKRj
n+n2WfCjR9tdwreLRz6Hyb8VPcgZxa/dp2zKZ86yfwCLdB+JdPDhrWw3YyIx
L6WKUyvpxTJ+Bm+hA2AVMPzG4/qU7raVZWKWr4+fuHD28NRcKARMMcSqxL9S
OBIObLMDOecx0PAW6Y3NG/nqwJabB7lD7rxxOga3uGf5ZSGDZEfrHB699DRE
gfjiK0MmNR53jVLkQ+jaBNhEvSp661MpN3E0cx+h1fwUFohzcxjaN759eslA
x7eSu9ceuxrSaDkvghSBP2Kx1lpxtLTZhsrgQ20115SQCZ2yc7KVSQkJc8ge
CwwXix2jTMkNYKqxS+76Sljm7C1hTL17QQV3YDWYV7hLPWoGlOwJsGftsdGf
tHy99+qDqfPlmrdxoJGCCbQhW24Tx5nTyD4RcNTWm6z4kF+qZ7TtL1zQWGYs
UQWGcwKnfEBhEu3k9FOajDgfbf+dbz7rpr5LIL5CTnt7K48zJoopTfl+F/gf
BtfkBNOHT+rOxHmWjD9+rctJUoPy1ehZdfGuA0+Xgy70TCvC7SpyXrQ0Zx7Q
etCt4NI9663FCjhwuLFd1yg7rt0gXaaUu4Mt4K8DyYL40hT6MhnuRoT6ObTQ
j+mMBMIIPEOKAzhcjCelu9VPxGuXkXaeE7KPG/HR8YArEfYIlb67ZaMy80JA
q1C+bEB1HkqKcXAplqZQLii0IJW3gHhJhTaQb58YlpwS6qUn71AGixvHANrr
xuEOa8Lsr5OIMJiVWhRiuxbvGMmMLAEC58PtXtc3KfRgaiJSyme8mCQVNMfF
A9Jm79r1YZCNziTk6EnMtaOzIPqEcbAG3HxBwcgDqmflrYYQHrwrp1MVhl9j
jHSjdeEWsFY+CVEq77FQp2G6oACNHXMXxxkJQs0bK8ME0bMSGUuAlbInWZNU
p0MSVe1lxLrU4ZNrq3NhuHK9zmaQts5/ArnGI5R+tS3CB4ae1bfisylpfcXW
HHgMhzf9TrrQ9X3dLievzt7DCH9IZXPAAAMZVu8Il7EDseBQnh6yJ1qDYyQV
ClGa6sBfOc7VeTTmqTDGVpnDmLV5JSWHnYEDN2WYsJXU5LvZSn0WH6SBUUiz
sFhEejhGC0lr+c/hLQgQx6+Glb+UOGfD/97RDUBC5KpwHSAurPDW3DlCOhPk
C8qKFN+C6oeCDHoDHpEdgKDBSs6gf9B8ySqkTep/RQgjwI2BrjLL21fsgxx5
72XlIIx283B2gLujPfJgNGlBwfJjUGtkq/Umwa2xDhdce9uZKDWYvgur/nxP
l57KmoycB4xeBpge01i4TOvKttvc/ONSRawRXNw8g4LNaZEXDewpObIdU31L
X4GETi70JqyB21iiJVBUBgrkaGu9IslQalNyOudPPtBsC/Rif2YmKIpUSHpL
Q+lXMV7sctPkOEI4NWl4ta6TXJdGWiaRKrEMbwSnSIqCnUvl2cJu4oSSpEkh
05miFzgu67c/ctR+Nym+m8Mkv9yfZoNCMW5IRJSrI8Hwh06t2f6d1ercDKXl
Z0JuE5NvWrH39O5MAsK9VtWNR+VmJ69y8dkI0IRdT8z1KvBCfJtm6mdmwykV
axdNHkhABSj/nqmUadK2+hVpHWq79PQD+sSHV+htGZfT3wASvWMH1O+VoRrQ
nUkTiT6QbADEsdRway2zDKnP38uPkYo7gcp4B3h+qPivPCF+sA95CCLNeZok
iE+MAAyMK9/soVAzengRehMtAPEXB8ViqYo8CKPcTOVaXgygYRHq5nfIal39
a/GCJbmzuNWVwb8+GFw2LGoZMb+RvU2qRlJZeTIq/I/6tpeZ1PbQHIaibgjF
FNz8zsfiuTimN76kLR9S3pmmyKW3cnTqL1og8cpO4ejhQRt14f7AjMwPCqmI
NTWbfqHT2eW5WVCOqqYiW0s3GZSEiGnopwlbGyXTTjedi+1Oglqa2z9pRXEy
iv9eohMnI67oriyrmyAOSTswcMfK1wov6wrrvCaOFdgYnaBbCKBoJZVGyLrj
/5IGiE2Q77znMsQ2S45cmTw22govwA0Hrbo/H0X5ba6nylW5D+RQpcv//Mm8
rToXB5nooK6rIGWOOI0/YKhV7EMskNOUDLJc9Z+NCgmqZZflffUYy8QC2ocS
0AZY2sRx2nt0xy3sBOAimptgBBHLIVzsikwypOScKMY/A5E2wkTO0tm6fIi/
z4rlLpT+DulDdLQm6D6VdJZKGchkkZ+aE8ATeWbbcv1xC03UZ614qyqCJfA3
k3LZ3DvLItRtk1YQ73cpnD4yHnriChUG/aUKMMxJ4GhHXQ77e3fEEzGI1ffC
77bphH+mVnwrvKn5QQRgW7T+JHFp+l4ynCeWezcOihQuffgA10VlJ+qt3rrh
V+WFcJhkdB4PDsLbET0EFcLxJcLQxoySg+8wC6xLK2nhl0Syfwh4Yo7sMBLb
vGkKXawTNVcFZBRey0wiimB8kMA7BL052pdOqdK59aqwyQBTSvZNSe1hk8CC
KMZVFz+4c5uuPT9WfoCiT3SwTHBJF5gSxYclX7iYPSuZbeSKjr3tB3PF/PPx
BfiY1qaTkqT/ZxRATD0+bHmcJZXiTmkP70eCa9NQ7M/H2L3/ZMD9fuQJPjBJ
vdd0lkgUPxLTQCQ1uZ0Eoc8fjl531FT0XBMAIv0ko64dMvDdWep2UpD8kmez
u1dVpjkhRo2JdDz3R6RaCygGMJWkGrAkUkCXgkhiTapZ+pSdwX4KbK+OWpQP
N76Ar72C2/EfhG7H3WZQM0ZXQze1wW0n8nbcJ6ro8VB9dRpvvU3XHV/mHRUa
zvCzzKlLGU/DQ7plBXbxPSqQOnCIbTqiYlGtWuR5JSsEDLEwPpPIOGj8W2an
kgyIKvaKgR6Bbifu2TeE4+T5iShgZ5jXR8pNPBnZT18wbsCM5WBOfvyqv1TR
3Tc1zvHrvCTgcSaee93SWtqAHMtaR9x9iOwPs3jp3deVhEUGw4UgWahD0odr
n22u5miIF27hP0QsVJhzeZU1WDDYRNj7ppDDLECja9BFEc4+hendjRCPC36j
rwx9k6DBLOtMchZjGq6uVD/cfutsFlH7gJo7BZ5e8fbl93zAqEeUYgvDo765
LXDpBNb6y2KppK/1nPyQAp9JEXTjRgEVB+gZV5M8U5OAtaPBHajNR/LRj2lX
Vj1mArHLAol1Wzan67kpp8AJLwnZYDL1maVyUlqZ1m85WSE7ANxw9jY3RpKT
1cl2RUFcTgO8gJ/F7/0di5PN+0sRaUmr/o36K/dQ8e2I4sBgPm8VthmyMy3y
sUN+0PvE5qVFWepj1CjrUnaD0j2sI7eSnYKhNRE5xvkMKyOFpTjERY41NjBp
bWF9S2g/LEzZ281lyivnlC020xwHE1FoHTeDMslDQPm08Yx6HseeYhIiK1tb
SclxwM190Z4iYIafau8PdgKoTrRnHwp51PWUB63BdoAt1VTR4Z/UmsTvXx7n
QK+fDe5meGvsE1Inxp9zbk1DTjWp2D4GAHBz0H5raN5MEK0HF9tiPP5mYjvK
CYsETgPDitccrHivTTHX/TPk41dvRxpQPDQ1qrEV2VkJhWshKGYfU3o+Nz71
fDrRa1sloPBjDOXxSAFwb3yMpSE3v7hYjgA72ci1xvKh3fqtMiOtomS81Ew9
QzrNjU15KhmvYZXSQJQBj4bIwBRa2fDG9B5sP45Vy3cd2GLz3r9egg65zB4T
hh1aMuSMLh+HWk+NsDgMHMeO5uRFOmcxl7CEz8yVSTQd2dHDhPXmWMzMP6yy
9MzPd7K0c5aRzbRx7T4Ct18Z053uOvalkHFqK0OQNzLLbrVtt3lH4cE0jeJ8
kvRu4H90F+yP2kI0BSM3HJnuldN72PHXiNwsWP0Ypu9PmHGjwD/CZ55+6h1z
JM6iZPccereJ6y0L5UMbXrZaL9gjR/Q8kwoaDulhweHOaPezW6NcepKfs8fv
hgCIkdwre72bbEk0LaF90ff3cKEY6iebNNcmfDpiZr/l8KjALDqoQuc9bQ0O
sIwskR+2hMZLYG8qBlXU0OHdIoxVccIAWYQ/LPxF7DdvneZ9fDL5WxLOCw0/
Snj904dokAiKVRGkczNuhu0H6kGJmi3I8FLXQM/X3yqGFAwRsfv5RDslZzlL
1MzJnnrPmV6W5hlrB21PEdRfyOLKF8ySWkfG6ZMwEJsGp4uZhmc5cEmmjJCn
i6YXpVAtKiP5hjC0QpFLkYQP/cXuuNty2H4IXhpqe8imCNEc2vCQ3gNpfKuk
qp98pLhFMPGld/VsnDKdbH0APmF1vPj8Pje0bZ07t0BDMSFJh/Ae12fUGjyy
bH0NJcm+GJAMtrHOMjlHQ1DlE9xDeBeUEH8kNoEfPu0ntjWDYFalHZyZIH6N
K3CYeXkiswe0trqRMu+ly95ezJ5q8ELu2DRvOO9VtJy6aNILG9dbkUM+vvGc
c3pRMwk3ybAej1mMpQ14rATbeeC3JctBdVipCiNpf5aq9Lye4ZuzSdCX8hGd
RbZPpDJrB4BVahUrcsi5g77BTCoUbqCDIzX0dbg1qsH2i8FAGH0Y6pda0rD/
ejaCTl0mDyIqJcyoFaUD96p+a2wldVJSVkWLRXs06+qT7KWYqZ9FJ+E87LZk
PC3aPCQHhfcda/yA6r62fZLJq45ftpbh9ONNyYfugCu8m25kTW39z6yucQu0
D7NjRTKj/Np8N1WDdnszZ+xEHZ2dhrMXcTJViy2MToKQfFfval/fahn5af04
DCd9KyW+CarqqyDO6atY6w76vvnoo6tKaeKc8D5tB7Jppurq5XcZN1dHQL/y
snRsCU6itFj5FqSUl2sIwt3XE6O4nytaqbb89W9LY6iVpAeLx8GPL7Hhr7YG
vBxtImmBBEUPFKzGvlGaEiFKPsabQMU+0kcw6mKg39zoSCE3UIx3XTl1shU2
knlCFFpnhqtN+qk1LJ5NZAiz2Xg8g0vo/enocg7tvO11J+vf4SC/G8wMKHpd
OEBitFrJmKv2OCYckhTzgVLsip5TaJxY3IBU63gSupBlOQXyDGcI6OcSRex2
hx8cxGjaidTGZDcj1vY07G7749dFYx3C5Wxq2q0fgqFZ1QXiSzVbQo7DDSfG
QcqO7UHcgMFQZRnLM3kpuKytrANBl4ZDBVC0uPg+xKmUYDmG4LpIekEWJ4vt
rxiIp3zSjf0nq5Be6/fJlVXoDEAiHvpaQZEh2vcq7jMK/M1GeVUjIH0Luv9Q
ejeUOpElaVhjHZnjUELcUoh6jjYuHGNw4O194gHQYZxmPMfmgJqPPURb9Rzf
RVidhsVr2EygurukBnHOSQX+SJsk8eqW+VullZ7xvZoMe/N1UFEY6y463ca0
TQUBdxZZwO1sBFadxohOBk9lmQLCfNaQBXjZ/usfPVW4TRngqCU8trYE7jEd
TooKWhr734wEZeiQsYhXREgN+jw31fLrMHZQbHMcIXiO6RD3PVZudCMXGvTS
/SDa4peF2eLcPlDz7qs2Dvcu4EPN5zJ1Sc4t0/GG4MKX6TN43AslEoj8zeYS
59ce5XkB9CnRvluSlHDHxngMaR3VmlduiS7p8Dbf38PJAERfVfVWjjbif/JC
zDgtU/9THZ9xOJkRAlFgKe3XPbf5s+6NL7xzFUpVFZlpK9mLheSyY0r7FkX1
Tbj/3sa1PnxZnISOKrf3aF+bs1gV4MOf3RanCIUi/n/y83IOUGPsq0ASkjd7
TIEkD+I3YQ8qbLYKZGiUWRxg5jUKgtp1sXWwPFCGt4WSUGjz5ol5t8Zzm5cy
JAEPRv5wGow6oUfPbE1xpx8dvFmcEKLRf/xFirSuPJBOA7U8vnzO3b3i6sJ/
ggw4X2EiBUw6ZpAhxIfuHfzdP87vaQ8XbQYl2h5Wx0gEDfJN+Pzwa8NyTxVm
hQ42yoTNOxEsEDKopNnM7N0BPalfYXd1DBi44lgJsKQoU+sH9b111uS7deI+
hHSmtHbjKLXDawa88F9rp673BHwkVvjN46TnvTSqj/Hojb1U8PuxObkq3xYc
FXK5EOO7efeVTbkNkDOBkdmJ+CMDnT4IB984lDKJKL3rxZYUxCOEjFUrw0qf
kzLay15Rb4aU5pcj/mL6Fj2sh1USaecCu5LPvSFH1P3qB1IKhiL+9JlysKv/
luxydrdas3m0mpYyw2NpNaaT1CJnDUtPVbB071okLmh/BP6uZaNLVaVlFzJL
E/u93OBo7IJf7JNvNEB9hKUf4G+H8gwPe7B4RhpcgDZsIIlGM1rjqJaTS3TW
Lw1z0ZeDbeHGYbiKkdXht/vOPAiowbrEC4FGUJrFoKrC+GBj9l0Tnrpki9gi
hnLkyGjMY+7YG7TjUCANiVgqu2dXv2KJoUy7yGdunjMoR00tLoqzcbTc+xt9
x7Eg1KRntLT5YatFTheSWHXUqNRKLD6OIIXjNy9uC992zhtdYgmYUWH0v7mQ
zzv5qX0T+szcuAP81Rzj3wsR29HPI/UOlkBxm7C+M0sV8GOIkwSJZ5vPE9B9
mID+KLhKFbdOiTlLKYPcLSixgRRXBmTX2vcNike2rMs9vc31vXdWEOKdCFfT
ZUSahHY3JNGHEhvmwhNBuKA4NrMLMezGz1QbiSJGrsYv3ycKuFwx1dbpwE4Y
JVILa5cz7I+AA2dnmuQasp2fvKtrSMNFo864QQGLGpyVTB84xshKxnBqETGs
6rep2BibJdBH+j2Gvm/wgAS5dM8wd4Mlees5fdrxwRcxnO+bmoW6pGgKvF6x
zu3DvuCBh+XKKZH7YcRVfO+vrIexq+BZEgi2OPTpLJnqO6nElkfEgNv34JBw
FLGIfrLppaW/LPmb1lhZeOJn1ppvzdT5Aai4R58eaLBe7GC1z+2wJONQYAXq
YSOIA832YC/menQDxSjfyTVfQvhK6KTAwBeHAXra1oScPkxe9B4GXoONiXgI
iabokyexEr8EHHJ98AyWiu1xxJNMNg/kVOy0+B/KLZcmeon1aeaohn/UFly1
UbfvklxsY3zLLvkdgomyqwT0jJ1vmgJX8E41L+ci0TJkzrlfSWx9Stycj5ft
JG1D7Si2m5SYiYZUqFvP5pohucegyqYTp4Z7Ie1RuCjeIkd8UJfkTuoZXFV9
nQQa5gEFrPeGqq09G1VfbSx2lh4A/VBCBMeVpL/LsLQaHJRVXE8gisoAlibj
9O64bKAdNspXzYNUpCm78Ki0esBt7RrDyD6V2djtN7mD6MFcfSmZe0LkEo9d
B34nHBl+L6umMYDC/O0XKeIAf//KsVhuo2J7LYAV0c54GGsbMs+UqxWbzRVi
nLq8xb6s6ECCLIWP5wEBsS2K/Ur6+HZZWX1T3ETB0M1CioJsrfkQKtJYQSPs
g5nNgXJOtbdPtXq3DuPNndvz7jjIPDbkYWoSaD69qy/IxG6/xnAs+J/mRlYQ
Dm0Zr94HmCnh5jhV6033XLNRLlkMGHBGXKiNWzcTw6wfRoLIGvqo5cWyNkqh
zxA1jal4zBrQcQuTz9pxDakXbF+NGZq6VINn5BWqMZk27RV+b6oVZ2BtL+VL
uhenAcYiDeLIYnKT3D/8y5ZyzDl5TKHovRDS+iSkBGHUHu8CkW4Gv3MaJ8NX
FuidwR7G7bVBOqnqD4JKc/6SoA1Iz6Ul88HiZPkK0nDIM6amXGq7R76E67BW
EU/ukNW2NxZJlbCQdRH9bn7Znv/CyV7W2ShHR3kZZPB0BsGJtMGBMEU9Pv3J
wn86PaS/YyycUw5086Y9ew4GGph2j9J+2/IjxZeCaR7X/PInQc88l0j0ZmeL
lrV5pHHlkZLut2EYgx6Vi7wGn+Ua8/sBoJ8aCzJofdbFhJOBbL/ldHMAIqvZ
evjnn39gnzmK2/Gw7eh54XzxGbyAwO915UejGccqqHTzCHVlHgSlwWBlNv4J
XiaXXRkRVOA9AvjDL/GjpSYYzxux7iprxLEy5CPljFsMsLk0kZH26/KVxMr1
SqRxso3xoOgH8dLydBs7jyOfVgpdBfSYlQdlzhase96z7l2tp66OnAeabsr1
+XjSe5rg1ux3a23+EHiYDMgG/JISkZzX4tzc5dUJvMlNBYjr3TbTO9O5EjjP
++LXLUhtqerQmklOalO+48wEXIwy8Nlh//zFh81Kqaa/l0VUrNUyuzpe971A
bjeLxXad8o9Q+PvoIeasbD5XyNxzLTd8NPU4721Rni6YYMj5WdxsLIGJ5z5D
SC1vwEn1VPObFyjZZQZi7zNJ1xTC/rlLDuCAMt31xip8dSIo22sJtDnxEX4k
Q57ef1BTUt+x0LmAqjDmjlgG5/IWQDQ4qMGv2j3JJn+7ysXEkV//aRi6kg1t
IG4niII68SQITM62kibNOvSgrzBcljC2ksZm6pzxs2ABWKyOWdpS929qPlHJ
TxF4RC+l+wcU+PaNuzO7dzpRET35D6muJ2vD8k7GQ+OIRKV6ELnuFY0m7oeJ
qizunqSZFBVKjVQCVw5+PqqcKWGTAmPpk9dr2bukWxKC7JUgY/dUnY08ItgU
sQQEVEusmztBTzhlMC4Lf7XLPfuBY3JYuAZqJ5vfmc5dkW3tEOGjgUMemH3X
9ohPK+VtmaUTKdAtdF9/FGv6RsjHE6O3QUBtZA99wPxVZP0OqP5pDQg4M/ZY
1LpGsMbu+v7olIGavFAE33GJl7dgvU5+buh820zt4g8UkmCI2F5bIiOtlB0+
v2Rn+7Ls+THkWOT2A2eIkeYmeA+gDTDpiUFx0U4USklBGigssxPacr+OSFgo
Y/qr49F+A87oWwqgCZC6vxgo4sRJ9DYtT9+iuK/AP/V5o9YpM4EHTf04u0hi
bPN3gIqK73tvSjqRYrmqh5iuJNqrbEU9upF++hRrOCP0EGYhD8U+wATAX+6m
jwKCBh7NiPnZh4IV7NrhQuOw+Ir76TCM1qZ39PVFEG6FjvkPx2IoSVMsF3nU
7JfQZrFs19n/tWCiVUMD1KpBeMffBlP0atUejTRaHybfHn113D5vmMDpygk9
KDS6qLphOZoRbMAkhTGilguK3ezBJaV4Qh+VUAwLxk4nurMxwkXM8eWhQ1Nv
70Qv4D28OaLEhApQqsk9T2abRHT5cFRD3n+cQu/9umKPNoca3AjlkRRVLj84
/b6ASL8oSe2U1CSMqPwDIqlUF2XCYJSsIBStpYmhF6DzBwP7ZanChvChZzZr
/7Yg29mEsS/Yo3bMs0J6JUrBdFKm/1ErUziS2PpNOxfrXngogY+twyWPizwk
EeWNfCqM0hJyVC3vY3AzvjK/UI41cmQA+Wnj6AHB2FXHf5sWF40A9lJMor68
K2GXBBCdEfj9YbG8CSlGEU/WqvYB0EEpTjoU67XQr32XuGpATQ9JZ/ErXBCn
e93NUdwaTWv6Tu2AiBuk+79R2DjhD69SzWdXb8evf9XPYR/4FJ1RoiXuBAj0
xp39foV1GQLzWFbyYp2busL3xzS02EktREzQ7Z7lp/VOP8ZPbEPzHHdf/Zrt
MD6ch4+xvaGcrh4/ut7jebBtzpwfx2Y13n4RhAGb4a24ZwV+i2vUs6t9Wgcl
YpD6quqd12tMJZ0wGw0NTxjhBTyjO+tKMrCA8fSYdCEuPyVLMCKXse/KKvN2
Zo/LktCWa7Rtp/Is/mMriCKwlhoyer7+bg3KlEDE0AtUcYzaZvXv3Rvbww+2
qVq88LreAmQntxFO6ugf40eMYzOOTX2PCbQlnR1bNIU/tJXTn6BwNsR86x1M
x6dHq85nm2iS6YcQ+FerclCLFoeYcMukO30t1IeT8v2wnBNEvn+kUNnTHn32
AOOc3cP8VGPEe+c979f3zRRWsId6Jre/oJ4FaN2OyZjkFBnh3+XKobZDJCeE
Z8uJH7qJDz7PZ8wNDhEKegeBWB2hHUUNa5gwsosio/9v3aciHIPYdUH+OAah
Y/jjrcM76/ByJipAeJHPDq4Kndzi/6oEIIVQYF5iqay+5sTt5lVwJgCOUmt6
r0LCRfP7iFbUnHiZeuAljjUXBFyQH+eDrFIhF7+KGIJDnYbITqwzm3j4sNti
NERaZrohzDO3D383Y++AtCsbsy8LnN4vgxnpWp3EIyMkcz78V6fSVHqsC+Ml
6PIggf0Kw+00lM5Y+i0/xvXI5YElPp3v+GErfaEqh2Vd5F+7PJ9BvFsQEV57
c52JrC25gAgRsEAFkxy5T7JsrA+c8EBLmnkObwM68GOlgltQsX6nPyleN51o
9+gObCVegp2Gn34ebgQSD/2VqFIoiw8KC4WEyXO4AtMdwwCz0y7TvTuVIlT2
kgcQR4k3EjJ64MWWa1gGzObHHH21SRICQkAY9h6AEugsfmA+HaC3VkQMwehr
JqhVoErBV5g2RetpadXGsVU3DyfkGzWO48qzmiU88W4MgXYRL7QkTs5vatf0
6VNBqcHRtaBN3rlkIxvcEQ4Ovv6/hEFlosybquVtK+1RhBXNHNWD5vwyklE4
ATOHtoLxz3xrsApHvaNpiX7agRmOonH8+BDtWPvkNFCfTNMSCmuNNzJ6afQQ
BKwyevax29lQScLdDh6rPqQmjQHu2NF6PpsmtBEgStJfO6mmGYoeDV0IwEMl
IU/jzPQTzY58dEilyQnoJNLk8aQviP8tiv8ueJPCzzfV9N26dwI3pU4sgsGD
NYH4vjth3qfPJAtxIPHWKNBz5pVL4pHk9bEQTPrPf1T6qlw4CP9K86eYH5tc
yRDRGI14oH3jAojp0kzSl4KwC1GWvokRks9QUXJyQUvmLxexB25+XX65mzUy
o6Oa332FRgm5w3ILpDCewF6/jxBdiSJAYgAipwHugvOxL7ayS4ZlGd+JpPiQ
jdAY6M1NKQNefLfrNaCtrCKwqVnw6j8Euh6tbK5xDE0X+KJstsHQm473souk
k/6Dho+IXIwq8oO7YtIonHf9kdnpU9Al79wyTI6I1oRC/bjKWQOLLv7VKmZ+
qmVKc6jCXQK5nxrcM1gwogyUq7gThQA7EHaldMStsfyOPDj9mSzsPvTgjyk3
OD1WJSCTKvBaEAHZ9b7axNm+vaDsHjnmaeoAWRPS0uG7WpnaID35s5iYpDkP
d+fxef7SPVECVpifYi6G7VCNJgovw/KoCqsZEamoXxXcpvsbCoBMJlpKwGS7
nRbrPCwSYXi8dNNJWWQc+hu8vZ2BcvDXp4vTCy9cvjCDEZEvy4GvtDuvH3pz
dDHpsOxAJcZmrZftIKaB+gkbYY3r9z7TIxPEOh/cAVICBzM4tlpBdRpVQZt0
h6n9e1fy3O3cFkUppbExzdixfD+cXhcg1b+LGz7ZZGIIKqEBh3gKhTRU3pCB
7020/hBn7CoR8X2+a/b8drVxGv+hRmfE4m8rmbzz6GP6PGAKLMD0KuA4z5gM
hXHNp10AYQo5VztQ+5qzpFuv9sHkyN9Txd7MgeUHPlW0y8fWtqdMU5pJWThT
s2mBrVWsGW1C5V2Ha8fEKzcsTb8VJmWveSqFH+s56Vsl0WNkJXzpfQ3SApIE
oKsfD1AvB4xtToQ/aoMGI6NMUWVoUvF+n4TvzGeQxeKOrGcTXwPExMrHwjp+
MPVlwSe1fY+pCy/Ea1kFJU3mhFGJcQO9WoXSZLpx5S3wl+cHsX7/kdJ7aMcp
A+9xxT/cAYD4jgSKAOYfKvd2uYOGR6XD45ucwyJwg7AMFEkrs668Jj0QroNF
p2anmWlvGF9nLLBM4lAzhIjAniNYOIsQw5oiNexN3QmZVdvCmOT3SDWAWIjl
XvnnSVREiM9s7wGTDVU2nc/Mu1kajZvqgv+KsHKNU+fjJYpor5K2fOr29YGs
mp2DhHgtlhwdUGKdV3Z14amoMhXBwBjX0tmcYtp9qEdNUQMzlE4AHMJNCc1i
ik/I1wtDMxxg/zfqMZQFgItwe/K4rEkNeYhwxezd9PtD/PEDktGRS2OY3T4x
V89Vg/w3+/eLiOnoeiONcvOJWfnyqHl1xQgn1zncEJV9IdQRfhw/7nWVlXPi
kVnwejkIdVJ1hnmy7+JkBLwWi898Js99ehGbrSK2rBGE9u3dMUfDxTY+UarH
+b6dMEW4xgJsXoyKymePeyf/Mjxm4f9PkgEeVcrE8Tm+6TbncHzGode616xM
RXEyuRHQy3ouLCJ1As5qjILWAvtFDfPEeRSHCHEnY4Sa38fVFZ+LLPvTHN37
XrMJqDjo9n97DLa5n+kkfLxcFDkvWLQrobIb49D9Xm/+ib9fsYovqFrCVRib
RHnfka7tRKc4BvjwdvQoPzqPSY7Whv7K25XaTpXet/pAq3z91ZWLSGAcWnA8
zqQzAKbTmzd31mX4Gxs5Q9TFpALSJqdSfoKQJ94D/JajM25aLkZmW1E4R9ng
CSnZdc+oioZU1ThGVwCx3U5l9kMSp4fupJzqstZjlG82lvJn8s0oi4fP1Gp2
BbSLBNWlU6aBcbwYTAdie8D0m3m3xzEJpn5NaGTawUP7ScZHA0pzT3mN5IBH
tL/8+C2d+fJSrDyVCSx/DaAn+SbXEGv9YneWfrch6mvpAXgZSnvfnhIJG6np
tO+/hZqEFoqCTSXjXHwwtuuro3IQ/P4w66QY67w91fLjm8dRlxpOFfgIPseV
DDSBHv2zZCUKUFzu29KiKrNZpEEyzwxAr4OrktORiXqccLQDvD1Aoipcljof
B43F30AgHgQa3iJiQp8B0KLiTuPWkeutLEDbDbTj27FNNAz2mo0YilqTt0vX
gYAz7GkYO+lc84lXsRwAOuZHTJdRfsIk1Aqaer0e0Wi7HURjDu0URx+QmBHS
eCPARGIBjtwwmxtEDcyF9P3klXG4tgOKOBOA+BFU7xQkR0zusxtnT9JECydh
grRnUp1flk1kTOwjRqAlnhb+C8dYlfXCNf0El9rNhwdXD2XoR38pAzewWBWI
EnvWYjen7opPydJuoI0hp/PHJod64Bz69lVzPF6zcwz5PD3gOEat2iXd17xr
CAlO3Xp3uHM4sTrv4sCGH3X//rHS+zIG6EeDhWCFhRDa60AWeHq7UPWyGUbb
E0D4buusztZhQ8gZhYm0Uaylb/n7qzNNuSS8qcF50jtpZSerx6w+0AvKpJ3N
q+sxNeQjJTLs3ksh/Lsk9GolqmzKr3SWes4geytjzkE/92WGcKBH9sLwD4qt
xdBWEz0SX8JQqSf+UcBVXz5tHU1hvKxvIDf/LO61iGS5oEH9ACXeVpLMNxPk
DFi2VssCyCS1E83KlL0mAxHJ34RwqFhfYSt9RvZrCMnhZle1vw5h6qApVZP9
iXssVinhCafWQycM3w3KlxkeSkXDmglO9j2bEYAFnznP92+edsSrL1GrEsun
yZJ2+f2yHm895gfRtYd9tui2xQ3SRXhsOT/U0YtT5o9k9RXQbzFC0kUsTWr+
cryvKXWK/NvjzxjXzjPy6AXJ8tg5e+xhkjecbtZrnhG56ANzqdLX8zTsn8I2
JwfPCMYEdL4vJQdOqSLHYy4PrkAlS5A7vwzGnCWfp/pokIAHrmK64imrOGbW
HjrnNimBwZuQuwM2mWMT9+4YRLayaa9gschSuxxDYNl64j7jRgHJHxapppMY
6bIeiI3KCnS/l9FPM1S+sAyhZMEbGnV2ZtI9JJn6xmU8p1Vkc1MvAhf0iUUw
th8eKz1ltqromHPEXX+ezzjoS7SFdYBptOpSZZMHTIsASvmto1BeJhq4Jw0q
zk8LYm++bddRmlXnnVIP9nFixfxAvIdO8/wxej381GILu78cXCrm5CZ0R0zK
MyHuBJM1NHoExslz+IBta50mZamNiizM/9CwDcH59wwhUOmZwN1ZKpHS6JNw
WwK+MTjrluOgaIVGmn18pgrv9crrA0q7IqI+UBcgX5s61A/s4g1cCfa7tfx5
xCcW3+gU27gpwEBSngdzfAI+QEH97I/EzgINMXDRm4PGoVHFP53M/xmPMrkV
/NLd/wLTYkN0BhvxHgfLLYLyHtfNLqVuwDwEnt3ByrYbWK07DkqX+ez31EcO
y55iyNpXta/GTmfbv5CSApyNaNlz+RzjPHcnCTfchm5PvdUY/K/FyetLf/5S
0SZJ7k3o1PbtOxbd1XaCafP3jhvl+Nl5F+6F96MrM2i3F1VhTAT3UD0RTzhn
qKX2uWw27BDDvmeusnHXnF7g2v6Ub6CdmShnGp2S8MNZp5IeRwtcdQQCOS2C
EJ6EfgCO1tewbj0vc0Aowmelx2kg+d2A28gZL2gexIgpVBcEixrYMvU4+Gq+
wcGM8FLrgtbEJ9i/fNHCXraMLJrM9G3lSlvPYIZo2I9bifQSg1jpFHTsZMRw
htjyRLZjdoJWMZwK9H3Bq5yUiTmMVIgpj4nphXMbRZQoa+7AvOpwf88zUz2y
lQBJVtr/o38V8/p4ElhEbTYOfz9da9AJXEi94I032T8ORGzpAeU7J7hafSEO
23C5itGzjBACzHHWonKpH2WcmlBhXWW80v5DQJsZckDjvsMNHWa+5gQdEdgJ
rFJvYB9vV+iuJk49ezEO6Ni2Wq9yr/1P8Qj4hth8/AxfalsPAri68tc7uB6I
3KtJ94LsSMv9/1hXzr8kf23YcAFwGX5EKP3gAG0xMFu9Zk9iIzCU89uagCRA
c2PDuq/YhoYGsb6maYEV+116sIBoPAjXrMk2YdsJOqcHW7SkbLX9JWYT/4/z
KP/TMfAW6NrB8tyqw/FjJlh6IVFKOgq4vm29iPmBnfj5NN+1m/CnfF/e+1X2
tV50nJGaJfbpPXTWcmdRiZlqX7TJGpGUYlgqdK9aY5FucxALgloe+95JOc2w
kd+KznZz/Gr1HoL1T016rV4tVnUZAEIWFnWQ4VPQs5or9oJnXUzEJmXAtZKK
1J4b4bdsKC1oK/R3IjDLXjmB5ZNwgci5sg+Nrd97UmGUL9RPgBdWTyt8Md91
sQRGG/2ReAzhefShMfH2BbThzstCiIarc+tkBWTW+yTVZwNQOXYGRvww80i2
Eo+OOL7K7A7GiJCSHBzpcWiJ36mYYdTLbGLdesfloBBdW1UbUmXMPZgAKCwj
y5WsU/8zr3b/uIa1NCOPObcUHgh9F2PqerjYGEHleQ90nAnrPl2ZHdglYo+8
AQa1QSBnl8AFeGpxOgI+hvTN3ghLF0ZJjCuavCGRmx8Ls86Z8zF2I6+rIE9u
eeQWEPwx+slScolPL74RY7prDaOC3eml3hXs2tAWSByYLY0t/3Cq6Wktq56a
9hrPzZEvQyY+NCcejeUqpJoDZbHLpsEYAt1mHMhCItqZyvO3EVLE2FILzd4Y
CQlY9dhynXm5JZ26JlyWnTYXNv/QeAc9gpVF36nf0iaN8W/gRbD5/4O/VSUQ
fOGbpHjK72WE7vRygIU0HGjXOj/4sjUF1NuVZSA1TrhRjKXMJDyG4BtwbwBZ
+yccSB9bPS5D8RAAxiu/cEvVlqbHv/maDZ8aIM+CMvp7bBh4MrIrPVqQW/Ly
8NV5C28hLDs3PYEWQWVYDcmkUDXvWROgwvMTo3/IxyX0V1AiaimqA5peIi8j
8FxKRQGXo4CVG8rhNloTpkTL+O0K0nWIYabWmkCE4LRL7+0S2MWWjTlw7/21
ESVYF9Pom6MafhEVRVF7Xe60OifO94m2HRT8rP9HuiiUmbtS0ljiN3FeD49K
qIZI7HHYAhUYGeA/fDzBfiSR7goo5G+cqyzobai3gzmFKFEuOziOXXKj4d90
7zDhQRKobecVD3j2MfcwDHh8jfj3t5gCQ4WFlcF6nWCpD2/ynVLb/MImTGyT
uDEx8Yy4CaMtp1fPlRGgPSlwz3VTm17oMNtOSlkjbH3oRuF+u/vWAA+JVMuX
4SdfoSNs3xd1+w21BcOzT6elz3vf0xN9ZNTDy4SzuIEp12QaLzQF/JKtjl0m
WHRZb8Tg2y+0s8ofq9PDtrH6FKseF0+jGjOrV4cgDxGsAhLOrWXT0s7+IZ4q
JfjHQ3/BdgD44R+VbWPilPIR7eVhP0zsx88Tb44quv6AVantZRgZHCesDfZr
tNrMLD1SiGWa/mOO48d4k1s8DnM/Ouz7iB+4F+11RVRkujOm999TRwY4EEbL
GayUJat7/cPOZzhaKqNCiPMf9yzecEktl5AjPvrNY+gkMG34uRyliCIG4o+e
d7G3SqvnsQhI2f3R78tffdIjGzPrLbnpO14BpsebKsNvZVz6r/5Yz3SArrNC
XS1yqWxsohVREdc836F/ELtc7AvLKNf9Gv9p9hCB2lkGtGfmUjry0OI5jsUB
XvRlCXFUHlNwCe55frgfMvHBo88mK/4mfV9kBSnd1mfo4Q6k0Ps9O+Ua7vn3
sudljM0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3EHmKIt0PZptwcr4wisDP0XhWbOeWKrbRRA/lWRkpGZdvUEqozaeoI6nxm0Dr3zEISVNNwArMnswldJRFTeTq7kiZMBztQz0zeFi6OG2DyT4Vf+O9+nhQjiDpfCJRdYad3gjla88DgI2QN6phXdAu8vmK4KHWzeosrjygwUAsWDihIN1DMAWgKJO5YJ/l2AdZ7XUrw1nRbtIRot1xKmiRhqVe5V3hcv2H/OYWxSEnaJJ+s7oQ8YhG6y6r9hM6XFbAqdLnJsk7m+nzDBDnyzWofSVv0FdGnqGxbfTjjL/w7VtCT8j/Z9w83N/FT4QvMgzS6s/stTIihaOmRoTWJJgkfGG35uQINlJNBU0JrgD9z8EP+VREBPxQX3hKquGS9DVLRJjMip2mjQGZEtFWJn4eXhv6nR9ZEeURXm+wmmKQJiKYhBU5aZuu1dUEDzCfLnqf7EpAbebFin9Qbm7LUh0jjHc/R+o0rZUcReSJZPVhk2IGLXqDODs99NDWIh5Ps33rO9ULPTWAc9iUsm/GfWpPT20OTgtsU6Jej33rv5NnQBhLIQByFUfUxDlj2B50f4f4X3umUG/JTzaEBxqslAY26IHAesKThamMXqFZ69EmXBGITvDlw8+FR5ZUSWOAi+tAKY/s6hk8/A/jAor52ad3NV9R3we6tu710XrirMEjzxwN+U4lFW52yWddTh8HpYt/nihBlUZ2JmlOgzMKZ77eTSdWp8fe+B0Xd/IX7a60hK0CuXAMoaPh72FRbwUnmHgkr7LEiJpywrV/qOS0/Iu/yV"
`endif