//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
y5ogQqwSvUnOr1lj/TMgeNoLkjlg7107UWRGUEY0g+kVyW2cgR2qBXN4Vrau
LjLDIGU4MMNiR2IkOA/VwYKCBUC1qnN/9umwMqC6xIikB0NhNYfdtJDCtyts
TqzyT/fT/QRa6tjeSo4p85rTHi0QtgkoUF7MeDsWZ2GWRdK6xYSSrv5jWRuQ
dhX4uPwA12GisLQO1NDeiBg3WSbKUWoSTFEx+1PTT5y5mUEoNubSJTAkIQeg
udyVTNXuzDZ4oigAz8xqj0rAtHHhjmKxGtNaUxfzU1ObSTkmZXj+dba/n8K8
jCeOJR1eMjLidHb0wUejjlzMWLwtTH8PpjKZKrhPIA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HkQGjKfPGwW9MMnxi/6xzVy9QHj/c5oUIFmkfPm0fpGzlhmpuwmF0/xhxcJU
0WiAjopoeMLETriGFbzmK0lucNZP3y07ohbjSMottWnp/2tVzIeRq7I3yKO2
zlqtNn6azD6N4WKF+AusRLmXQFmSi5BzEUeSJ3jfj35Psc6znYyUXCIeiCND
X5+1+P/Bzbip5sAb8U2dKOeNtWb5c3CSv+gW5CX9/Nfu52ty+r5CJj8aMzUn
+McaX7W7VxjU8b+2HnC6X9m/t4C02LEoZ7nf0l7azxW0+FqMSM5hIud9xa0v
g4sJD9wosgftfMzdu1jzCItX7C+/MqD9b8CPQouVQg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q7o3k3vbKbKvBENmhcSTU+20tvahP0fyNv2Rq2rcq0TQNgI7wZbBktPMjNtM
tK78+R5t2rH+ZGa4eTd76/emmJ0Rrti7hxoRf7vPYl/l3bQ7RBUixYvNr9Pm
hiUI+ZC5tdJv7dkmJ4llVkDkOGaBXBte2OoT49PIeeizaIvrCE8akQ4s2zp7
xFu/LSa74tQrUE6HNmUVQ10oK+gi0CQzU43JFbQt6hf7udG8+LTMRLmgegAz
rhJTFkE895+Lazzrx4a8Nm3J4dTiIaH8HSVgQTOj615gRFbMcwJ344GKAVGM
Cnai5RiTYyvR9SuCo236pIhLhWgZJImiWGLmLtw7cA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fXUOHtfRHN7Ll2X42Ezd5k+dLHRKPp0ye7UgRxZTO2NX08mA6eJ3I8nDeaGC
u4JapBXexW2jeuOoO5pvbZeNtbKWSTIfDy0NEHIiot0dQNiRE3s0r2Ra1/aW
ol8m1c8yHiDNYBy+TVT8dNAqwJaQJZ9kMpgJhYm/vQ5ekwaNZJk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B0dLW77OAUULJ2bPA95PXC3RdL0kg0RGbk/HzMh66VE3+D+FIA8Ryt3gA+FA
lplXu5jAKdSd4qw5/K42R7y7Qx3Q/sLoslk6hWPkQPRXMtZnMimE+YC5AzhU
epXyxVKTFPDBOYwuRGTkF/dO/t7WTRFy8quxw3wIcmjevqstitYv93k/feXy
F6Uveyd6Fg9gdzI47rSoxMn9TNV+WGgbquSaIh0YLB2nPpiywRASpsbTNxki
ikgR6/vKYV7wTtZn7JF3EaZWbk8yh9qGB6mwIwpvYChnTVPaTH6un0LJ78gN
uUuyER1NQT45oT27hYjUg17jZesdWjlyy5R6PCyHHdTs2fRFDAinpFr6wqMo
Kns1vodaaY44gZpMyxoI1GMYBrLfVc9r8ZsTMlKjGcYZXr8cc8EFyny2YMH1
sW2TPd5I7mhBZZP94NSGYfIEPY7vwSnjITE5R+C/PQ6B6AAXchjfv98CFpvo
3/qiSdx9LZ3pUwVUzhmh7Xt4HgmTNeJ4


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
tIJOS4qZf2imm8uG3+1cDWHeBMlBza0uutXVhbCR9+7NMb7QZnDWIzvmWx+c
90CK7L+PyFNh2/fTApjmPsvz+fPRsSPsm3zVpC3P6o86GEj4N+A348tnWVEx
ZzkcxDpqzQWRRaY4Y69ZepDRs2UbS95Y/fpB+De5qB6JdG1GbFo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YDGEYkWof9TcEQ46mlPEEs74bOQlRBvGQcrlDiAqqZoEmADF3VdvqJKHIXJQ
vzQEpJfqAt4wzb+DPLk2l5MknE8remE4Y7EX8Iulxy/hxRjbdbnZ4JidrhBt
IuzVTJa/nEbPNda9Z9fi+Fb6gD+ZQM0PbfjSfVBSEdeGMK01aSQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2880)
`pragma protect data_block
ForAAUbPSH5uZXk+s94VIu9mghp7SvPWUWAjbFjaB6CEFPvErfONKUzZtH0W
geVrNerQ8q2dOTsd1q01AiFQ6HVyEoL9vQu8ZFiMa4bPZlgtzUv6vBN/J1dN
EpTRF9n5SNQVVXbt3Xn9YTFpOeY5GlD0qPTSJbg4+rUkClXpRklcRSKX/gGC
wVY2hKEsIbZZ5bM8FT7qlHUqJ5EaMgUQUvk6HlKqRBdi+Eb2u9cmUnyR1f9R
nbfKAAVlmzMsjyd686JzsCZnpl1L7y915cNYU+pcBL2kEVR4RbpXimlS96nf
/vJQxp9kKmNCqlLcTv2i9ZdIomTqgEfc8PotHiIXddDA9ZOcaPlQnjzAGPC0
d2c6U28u1qEi0staNb1svoX7pBd/7ueCVyyKKbZphObJcnJ/blVefXZ2PGPg
mpVQQQqrW0rN03WpT0HLV2Nizs1gb4Oep4433DqjRIQJV1bNCm+DE+y2XGJ0
6n3B3NmEV1ZbCo7jk1bcePIDnTk1TRp3D0xViy44AylRki+OdUuLPK8ifvY6
YDRC+EJKbWCgbMBwTa4RrRiy8Myf1S8seU08kF4BkthymQs+elPywQrXXAB2
frhhbCaQuMHPN26JzQuDZgKR7Ha0zKlyvluHzv6MzIIDihup8p4xcIHUuqwO
MznSgtT3NyZJU3FLQiBvgHA0vHhMvn6Qo7tCxbmk80dsIjhrl7Oly50/Jys+
ti2S53tjM1ERYMtUjsgIrpZQVrH3sxMAKMUjlTXjdJ9UKOB/8ZK4uGbGIE1i
Vv0TRPizWH3B9yXWKrOOMt1XGj5L9CYNprFpXEzGHjOx5cx35JXTV03Pssi7
7evs1yO09wEz/tqdAAn8sg7hVi16NKl4/Wt32j/fYq+k4nRAtXBDWlawsPmU
4RpXcb73nrMF8cR5H1zv1hQWn9RqPB4nlEeosR3fTNwEefnh6x4czKdHZ6bu
7QTOcHJPIJr8Gz2grbJXsjRXYGUvUtThBv7v20bm52LrPByhsn6dh2low4E2
lPGOaMY2T+gjrS5eoA9pI+Eln3raynI9mbFZjL9kjwrGkWXHq+NHXITH/PK8
NJp1Dg3bv4LTTD7RZ9dzjdCmI7Nb2V4IcEgdctc/FuIffco8DCY13RVYmSjG
Hu1B3ffePjikYWqiXE65+nQSaOsIwM3t83L8XQx/8ijDGK3hgqfYEIQlxE9w
QRFvbruHD5uGqngRrN1ED2z+kw+hUiBfpNQrA011Vo2xSdXqXzbKs2mt/ThS
+97gmVjR9dLSFxmRGHWvCrkN5CEQ0scL/K07Rz1twcfmOf304iBoZwStJLFo
YzFLbtN4khLOpbiWeYbMdKWPuzEUk550boqWi7C9KhxxCuEnsR+PG9I1P6Cg
qY6ttG9bvTpqDfrKIf1I0yH1S+gDOweJT7uc/ZM2I8EWQRFOcxPHWS8GNuN4
ongL6MXp2TsuPWRAIovBP6J8cykPsV5WwJVq6Do/0fMG0VnQpDeRXY1LqkRw
oZs3Lm9x0KgKLxdqpNWG3pmiKqfOH/U1vQBp+DPysTLc1lZ3P94v3FGKgezD
PIcltVtx8+4YMqfxThNh57i2WoW6x4aJspyPmgoZeG0gwoG95XQAWI+pi2UG
dtk7xSQkTEKCMVA2dyBkHRiV7eOmIWjbmz9HA+rQC+w4RBWiirHQZOCWswx9
1BgyVhcmolArQH6qTdPsllPpSK4IQnX16aKIVkoz9+RbdB+HDfw2CDp9M9lh
/r1rveON8RX1ZqpB2Q91T072Tzl63Tjz6JTWuABwSoOPgWqNdxNs1VFtCfRJ
QuXSOmHBfjBFyWeMrUVTvwU3f/n15oflc5UBv1UhivT7gSbcWI41YcPY1wgc
2Tkqhe4B57zZXv/+kLK0Dme96omJWsJ62DcoxJC92rZHrw45r5ePGXNsFns0
L1JAeQckSav3HmHJIs1qFhR/v2pv0CrJCIY0Xa2dRp8y76X9/B5VReSalvyA
aTgnrHjdZlkiknFZfZlbqHPLHEXqW/N6bo+o+p9cUs2w16FKdKXa7wHu0BOG
Ta/9LxoUmfy5vc5z8EPGWgOkk+7T58HUVMRHZeT1w2FPyO1Vw/ZCa8HbBf7H
EpZhQtrww9DSFepEXdOIOnnKeW3OlZPd7F/TFBT2P4RiUc4o9iYoz+MPO49r
7oV3v6jwNa60eCdD7ppTAYkZIuB3YXCywYzjQwM3W6cCgK+Oj4qtcl6ZSiYS
3KmfNIh+yn/QIALScr1ybVwBDqpD3syqtn95hdi1DhGnFsb+L2zwON4EidAS
E4xk2au31WxdJIPhYXL+2JqBdNyZQ4IYa6mgUUVTWFiXyzmmy8WB7R5xODy3
/b7aFefwI8t5q4cr2HADmCPkDiEDk251lHXCGcdeJn16vI5ekc32+VBwvcYd
lnV40abaqIFrZLyZzjnVjhMjhxdwlA6p6hF22m7rEzbJr4Vc71CUE1QMFCPD
UtqekAUzrW0J0joytpQfnOtB4rzp6MVCGVkGPxazUyt3m/zXRFFG/7I1lWez
3fx07/BHCENti0+crivZD+FaqyinVemHbTl9Qi6NHIrZil6xNwxGOoR/LTmP
WkbJr4zogSJuFfGjHt0ZzHdfc51zoqUz8sgI1+OwErnYBxia+FkhEqFCYi1Y
3YrPwdUMlIHbjDvNzGR7J1YeXgoRL64Gqw9LYzM3keXmE8ETMizgchnzmpqP
8wAxM3Kt7asbe4bZyOYB0BsOXUqg8WxFRG8gz8Y93XKwGnBjULc3BnzH22KH
+2voAg6PwVa66M4k5qWso3ZbmZxRlAzHcqVAvBEPD0GgM+xiJJRAR9HoGrcw
hF1D84yggMcnHhBP7+s4M60Ei8H0AF+q2xrY5SIzCPnvhpzMRzk9JL3afv8I
KrjkKGHieiJkmb96/tmiCz8WGBmT0dk0I9eyKuVJtwwJU9bktLFHRbNfar0Y
gCy/WzQNvmUIPcD/9QPhbsKJydOLiIQZg36pkzqSRgHRysoQ1P8k980y/DqS
Cw9zmxnOkxJEH5GKKa7D37Ah3/n+fu1ze7ETnxhfuHJPjIqFBrZo87bMSV9v
jPkDTqopJdeAKFrz5Hu5D5n8hRiT9APbUTVL1QXnJM6sqsSpMYGufJh88kb1
62CP+WCsX68bZBFbTxD+uUznTXvgQIuM1ScPVKSBCH4iuPlzei+xTwPPBIPY
ulgmN9slLljZn7hwsQhY6sFtjG5LiNBxtyfXVfe5BjcLCayIpyzSCVMHQ71D
KBnr+69l0iEGvXiM+WpDmZ07foohz7rEQL8bjRqu3QI/y2oR+/QnDK77FtoX
t81pKufz4K3muFmsbo3Ao/cLY/ywDI+ZDWF5B9zvIBL4Fd1R12RPXsTQ6Auv
DpjxTSO2sJdKvJWoS+LMUDa87Tpd1WiYIlaaeGrog1RPunO8CnDnLnW84vEd
/gJHOh/FS7Vfk5q5CtXEYU/tJRNwvf/sE9SQt1gXCaAN0FzpuPZgdHtZZ8qC
9oteuDYeMibPoF020oxLLY5FdOZYXbDtkT0QLfkH8xkMBVsd5WP7PnjT0sHe
JwigWNhhVmED8k1y6S62zaIMmIokt/0184Qj2CUYcokTbDD/D4D2PGsYWWMM
HWwSTnyUX7tO2Y4TlMyKAvxEozkSSt5GOZpVJbcm3NoXVfNRu3bJYKsWW3W1
GquTfgTtIZWukiNoP+IxDwBDvkHs/CM8K2KCjxCZteum4mI3kG6ljaoAnW5j
p1InG+8ZmK489jeFKdpDbxfc6g/aoq4YVsPpAQD3+aA6ubdinPNuvZlnus1+
/5UBsGcCS1M3VBkd9lzhzow3doh0iQUCVoFCeQ6Ur8TUtT98rYKRXsLibn+P

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG2jVeXzh8KOY4qCCu7f2HIjN/w/yVsOVzARx7Hm2+jvrqN6ntL2ozdtUCAdl4tygERw+Qe7vnjjuHhGv75pTyY6avAN/6um0zQIbQLTGgc7wM1c1bsERS76NK2ehyrZqMHWOMGEhL7T4ASHnvWVKau1FvWCfPVF/7g1l+X0hjjrR2pjvun5P8VpNtrBjWB9HbG227dH3rY/szs/lUEYcCwqPfABt2E8tMe7fN34kr0EvRoPvTRSf2skuYDOKb+0xE/0NhJ8xSDqrUWy4rC+Mp3q7kg99a/hJRrOMHdJvtN+WkOHGT9DgNWvAiwBXNv97qJ8WNN3u2XnURihVrPJ/E3/SGfMbxh+i+EhEPh0hCJ0ddJcp2t6j5ItuFQlnYzSjadzUupiDNRrjvc1k+HWvA9s/bxqKe5J91eox5gQBSrDdjWNr5N7i3xxWM6t2aDX6UFCEdayIL2a9TckXVIb9PgBI0422kcqXy+EmTjpQXsR84nv97fjYzViWqggTjtx/uganXVPYS9GAkEssK3+IIfHrRuFAGr2UIdN1lB+cwdIv3gAh8wrfZ5Pz3Y/5fPjzh9GdTDdqaNfgzAgBVm9qpp5qfLIDJPZEYnTGu57BFDN04x0cb1fhFrxlIRZ7CXeCN0ByTmtWZlLiXPJRAqjPRPlFkejJcFfh3wSEVkd03aPauaImcf8gQyRqFPv4Kd2pMy/eVT3adIZtGXVnwFEUePQdkbNuq0qEYzq2iktfVeDTmybAZ7o871l3ED5Z22n+zJGZ6Oaij6q27/UeeQOkfio"
`endif