// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
L/NnwRyFHLQyPv9PcAzvDLQLEiZUP8p6NfzdQCUBLxjEzrcOPlarYWI85uX3
vK4T9LUenXQyBFy30i5Z8XLuZS49vzAK+O6fecrd4gESPh6y9TZefKpZ5zhz
pzLMFk049SmDG82hEe2Yit+HmTzcFdYCjVvmzADTZMpTaDwlOyOyfiyNN7jH
N7u7M6H8C1fHhqLuHJ5cK5RStLKdcDtqgQBXm7HwMiokrN+SA/5gRJ4H9fDL
uWzrpAkK262IJiAIB+ZMaB5Qj3YxxIxNgrAYmLmYYMepjaMi/iwbHXvwR95x
/8fRnB452Q0CklNDL/LifIfHiMJvwf8NdLX/rAPdbw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kouYFmrz0ESPXZ5Y32K6rlK3VWdq/8jWDPdDmScLQSx9U8+GHW3dZMQ1WVYu
WA7JWAwQcfWs+0VDyS3Qh7CzZA6h9ihEeSdShtXxYKki0QXdkGOuOf55PkX3
dJeLvZVHUDS5H/Wa3o71hR6pj1sGikwDGAiZuBIpY44fUc0f6yB/9Y8BtpnM
jB9tNRhKt/g/ReiKIeZ7L+kQW8673PKq6VePUv5fIvWTUqanGqeUVtlKjjwg
Lbfk9xlJqcb0vw45crjJS0xiMKuq7HkUlhdpSOe1UwjQEJYsSQBqQ8JGvgPo
/upQ3ag3BS0fPdL12Q3WFkeIgsrP9hBIY+JBii+N3A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VrOstjzPLQoQtldRLoGD3jlDAs43hXwT9l3iQFEIaMVaTRy89IHXFTZmAoYg
n14UrOzEmiVZoUnu3qQfathaBRi/d4Wd9PfG/RGucXBW4UfdPJLJy5wqGfVX
P0as4TPwwOBZB/L+hqr0cVEUK7pohHP7ipVg5mqkUdcjpYARtc7y3QTpROmP
RJcAlhIvXChoeHFVuAtsl+3Fa2t/gY/KykoANpOS6aEBsNK8rELqDnef1bsz
0iHfUv8gwOlWojpvKg6cD4EYbkjbD13OhHKnPQBnoKJsctvWs8Ll+oirzDFf
89WqhyKRHaOSgibXQpEoeazqAmnAqc+/unOidvZUNw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nzlgZV6+mex+7Mu3W9oU2WzQXSbPxKJu9keiJ+erNnYwFe+37ojDs+1ljdOm
KM7SUQ0zlT2A0QKCx9RILHY+WlwKN3I6xlffZK6bUgG70H86VAeUPFgaHZ6w
BXMSoFmNAK1LEkKA/GDofRjldXyW1lU3t5DVp5dDeS8bKmSZ2us=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
se3wyqjBKPd6hDuA27nL2akbLBQpdEuxrc9tSg+VPev7qYg6LUUymQ4g1oEn
aMJ0uXyvEsMsnSi2IJhLqFKVwoJg1KlCAz+8n9f3SXelbs7rE0GmterHHvxz
Wd4S3aruoxQChAptNRB5rAjTfTp3MUBdo7yrlifbH9TPlksm8c+6/JEW30kt
wsVcRpE7ItGZH3ZQ2Sb+Db2ac+FwlijYOrR2JS9qhYuQYWn6jS8M5cT9lngV
KsvF+UGixUC9xOlslJGur4Y3KVvQbfbgaMx+cEvquY+jFSMMNpgaHwVPsxqM
X0EekDbxyvZ4shrMxQLL+mA6wK1sTNhiYNHtiAlWfrBSas/ROQt2LCvG8CmC
IhoWpUgxGKszfI6AlzjmuNpbOabzM7IdLoojz6iepArh2N0rcnOfsDToag53
HF2XkNi7BScP5nzXsCSNA/05os4K1c5KF32zjnVH7gm02+r/GwKkFhyYmDJr
fn3XxJT0RIllgru/lrvHPrB1onkudj8h


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UrUCjDja4VpSPzTyAzYaCNLsi/3aodWesy6hnw40C/B0Erv3eq6L4pGYlq+z
B8pPeEEGGavDVDi204XqkCltEEXnmm+4/oOovWiqpmqg+hPC6ExsB08E5pIF
gxv6Wa6HVZgv7DkGTpKXf8BXn1pi6iC9vIiDnKOQhub4zOhZpoo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rqY+eOzLMSe0GHqADKC+FZZFYfqwguTVzhdq8SmrgkD0ca0e4gY42KbTumwF
l27KiKc7kPwynsid/SwbLPt8bSnZCdm7WjyNefM7+FHwswE8iccb/hrYlfPD
SY8tOyK7+NSVMofpwIlu7/tCQC5zeh/qMSsUAUwiHGOh2FrR4jk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 42272)
`pragma protect data_block
mNBHcJO8GwZqYWb2xskhB0QNlI7wpgNgZ5c3LubOVD9CPnm/s7WxLLL5HTp1
f5hqzmIuNFVjlVtyZnICZEkuUNcYjYE2tFYnkU2bekgQbztH6LQWaA+rmHHQ
rPJXwqo5aBUqmknfMMjCpzm+PQ/FcgTKm1aJzkgAVzIsL8hUh0lIF4GBaMfi
/cZmTUqzqkJrpAYsKGfqq00lhpupnDd2Nk70wItCNC3T0seM3IqZn7VxX1+e
mdTVfYH41eCTjngE4vRDYF3cJePTWdsHqcpktyHQC5ZyLNx4f/+h3Ep+b9QJ
/UOd/2fPn4/v4TH5Xp3oUMnVvWT6li7Cq+aOfdsWS05qBrLc4vs0LmkB7Pax
1dhASoxoQdD0rP0a2OJc+YBjSI/BvgOrJtGqQDDS7nJrT4NKUjPi3ST8YcUw
bg6DMhxHem1LYR5cEH/Jt73WPDMZGQLJXX6a6Kxqt+Jb7WDkolez7pxSoTWK
b5UqKm58pEXhQIL8RrsLxSeeYAoE3hK/vVEVQTb7LDWz0hDnnzqrJHgyb4XD
k0WrjPblYYuUyA/QRmGVu5r06GC2sKnnCsTTXXFA6v9MNkZ+q3v0hvPegj9x
VWpYnxEBUNZSzEj4cC0fFAo2DbCSFoZJMwZ3J4IJOzAhrhOND8NCJxnfltuW
Ap1i8SWoAIb5REDNA3QYgt7+EGgjpUlc/F6DkmEEkoOVkoxUfvjaysXYiB0n
4l0jSR8XNC0tGiaaFXBD+OuwWFEIpaLcL1a4wXVwRHbQU+NnwgdaIIA86b1a
QoyxYhjauoc8s6xwhK3vkV26o06hRhN0qbw9FrDSTwc4dauuNOffjEWcS4DY
w2/Ls0uju2MtiVrivbTWIJfy4pvSnMiTZJX3IMMSmElEHgX/VgpvSEq9Cm8N
Xelu9PSSX1UfM/eSJwBjr2bMySCqV2sxLSd3P4YXrbuSJ1v/NtwuqooBvgiG
nDDkzANowh7GHOoVF9ZqQWXUmQSy0KBFcPTPQKGyO0xj5/4V1uXDqQdWrXQv
w3rYufZy6TNvxWQVQfqHhus0kVML1+lrAy9XajI2RKUyO3q9zuM49F3mskoZ
e14fMcFYijsBsg10in1YLIzimzHJEVJ81qVmISxaEKTULIeoDrNY1bUjFbOz
SR3MRrOHAEVrt4tYKLUJorPKdA1wmhowQPVBkErp6YrWu64HkGJFYPcqGZlX
cShh9nArySH4oZM58SBTUNCIMindPdr/Bi1pdJUR1T5fR5HiJOQBtA30Vhag
bK9E8xB2tQGfyZLaqauD6aMRnfZ+uDBjdp8U2v+0R9mD/l4vofRIS8mOR/F1
YnBT2U5couNKXSntb/WBI2gLg9zOkCcuOsWEYrNI7CFcpxsDge1D/CoGDUis
vInWy+Y7+eSH9xMJnKBdEqpA8XmkO7+gZjHwtBhgXJ2GCb3bZ8Qci65XylLQ
YZW6ekahBSnFNhK0i9GDxR2xBEI4ZjjspXjRcyWHTEoXcyq1k1L934cJXojb
Pi02HcLOKTm8ho31Y4421rc0gVO39XJleRS3SfVw7iO1egW3eNCNeg4thFTW
ofr9VRA4K7zr130U/OqJ671qWoVAaXQkJaeaveGI+1+0/uB88yjsc3qXS0mf
B9ssaR35pjZN4Sf6u2u4viVAePoEsdOUYDCFPhlYsBiEEtcmomqYXGaTtG/M
QLfBXPNTlLS567rTjwi3C1dPeo6qR+E4fAEevJx7/VSYRTrI1A84rM/TOfNu
LFO/lHJuezfjS/H8UXip4W7oOn8p7rI4IXyK4XJT1k0TfTHlaYWnr3q3BlkQ
8oNsmXRCxuHpKRe50XyY3oKCiCaadShapfyGzFCKaWaG0/CGTN061XoLtMWx
O8zqUj3zOkkfBLnpR0+nl9NAVapvCFGo6Jnlt3qfuVj4kDz02vJJjnXtDYHN
sCOlUjAMTTUt1TDNnpPKFhBHAEUzEdfmSTC/xRONhq6/9pXm9zr49EJSSi6S
jC82vrkIYwkHVzoahbHADmXQR6Uy/0ACgZtnedObfoKdscKWEwd0dSTouN3k
poCrjJTlVLYrPAwwbRe7angwO3+NLeClQU5O+kFh1UjaTrGUAhFK0yD6Eqn/
bsPzXD4JyJVndsMbdoJtYkikJSt00eveIeDXto/68rbCOii6B0AnrIuj9+rQ
27FlwrLtx6hDZe729IaPYM/+o+ehUf7Gc9vCIVZ/MZCnLsSgtwyEqdq1/6WH
qFBdmjpvMheG4ZDgrKymVAl2eLqCp4DqZs9RBrvz2tt5QyysTGwFitk0kMCL
E2Sp0qqwwn3n7YFqawx3R/TbsceL3nwWc2hUnOeY03qXbLU5zZa1UWA7X0lD
qLN6oNQbRmCPGtBlJK82xdJMo4hKOH3ZwHAzUnCACmS6R1UiUT8UOYwovOD4
AxHtSpVQ75ONYOGETT9bHUeVGqhzbCE5ezPdh2DcFxQsRtLXn674URLJdkOU
jrUIZCiWYLUjcm86zi4nWXq9JzMvkYVpAqLPQIKP9t9TyY4N7+DgWlRrD5LU
q9myzTwt0xT67bpTA1ERbtgEzS+gS3+Vkwj8vR9dYER4PsFePI4Cwj0/lT2V
ghgzTV7M3aaBwQAn4tTWshDNP7LDbpLYnYctUm1rlHm2MAuuzlBrcciycgQM
Pw6x1EffMfRgPJjh3W2IgGmmDxzy5em7d2tKOQuVoe1RTjnRmNjbuXnEvZy6
WOWVOceRrw0s854CRCUlsld3yZAkVp5BGoR1rTiqROlpDHHPDkqciq15HoUs
YfphrmVEfVgwcdePgvK+cRMtpQsLGqBI8fV1QTKhHA7UkrzKod3cz9HmqxO+
TaIMSqjslgfvqT+Blw5A0+IsMdtxCNupT5ZnOZqEuF2CCnvhgseJ9WtFPlpc
wIWpj1zDzig90QleaR/T2XMdwVpmYkhKNp2aqjZaUNVd+k2L+wB4bazVfh2K
pvaUco8SnUNNjQinq7DDNUFJdaKrmsNDkYxetDbgLWziVAeBYZ80qP1FNzjc
6shMtlTyVak+4noh4kzTOH3TqtGIXrFUxCJ1X1MSO6OtqIVZUls/sjfZTO2P
E9xYpk+7Y/DBEY6GsFTX2dei5dN0Nv44/xcxEnW3E1U1j3Glqj8sWQw2k/5M
+VBzRb2rs/h5a6kr0EFEVlsm9xdcCeTKmBIZvLqxOSpi/6uHrPTQ8SxPIDSq
IsrPFHmttBDFzGvFjM9JFbQ8pceuHrPxRuaRmcOtlaOTGCZNidqhF3JsXqwl
HXJ6MQLZxmRya89p0kyMH70MD7HyvdKpIA39QXZz268bMxSApgMyAGMfqRmh
vs9FQpdo6QJj3pzXs77jjbUZYY+Vu5pIuiVFGc+stJqKcut6jnNSas9l0nXl
Uvzb9pg5tFYHiTpP6KGuUfAihUTL/LSr1Gh0/6GA5dJpmFAcipyKxWGLF3rO
AKRSMw6joTRow8pR1F8neLmlrjNJ77znKX7HO9xOHxJoUHElhiUqeqF5npHM
h0/KZKOMNNBwPpckrPjvewXYXM1Ui1/8j07w2A8DiymycWUEKQUnS3ZS85AX
esL/NzreMeqPj89Uw58rQseeO0xb1SfKNMoveBbuG3JwCySWUGks944L9nj6
YbkOpb3/Bs2UvGAoOblW4dmiU0jvz7Cigim6zOaIPhiWEvYbpP9keYCEl1Ya
49yD2yVOskewRcRmSVhfdcBzQGaUNvMn3D/0cCRLTLnBFJxdRisHZIPWC+Sn
8j9OOJ0ibQ/XK7s0PYkY8x63W2iEhWmoypHEaQCIalhgDOxuz0KNolJxxqJK
XcRg8i/N3gMIChYInwBS7cypYGlG47/KWxfrKAo+V1nvQelN0DijA3ktdkf3
vgW/PtUQE2X5FNoGzWLPADLsaxXD3wvoW7qU2BnBAuOsagAIyp0rhLZV6KoL
Y3pGtewCCGFPKIIgr0XPtJ1y6BlYYHaxbM6cw0CNUruxJkPOE3c7A6Rv5lcY
74vJKvbdwkvAKGrBAyqU2Oj2v5ragmdEWoja7T8jeMyTQXE+7rZkS8kQiYKF
scCDCGYNcoxz4eS/EJVuJ5AOg1Lxkekrj1Hmi7U30G7ELnbGNzxfk7chkmB1
Z9mbPWIAJFo9fH3SjHV0lqxr5QWIvn4o/O+8RiR4EssJF1SpeMN71qGuBAYA
VT5eXSYm6RJYSAv0r5gt8bx8qzkJS2WEB/KgE2JwyRbAl7IYaa4Mkqbcjwsm
j0ATyss5eZnPGTW/mpUL9LLWSslYNKASIRLGi/0W65ilZVD8hNYSrkndEaP4
x/JCEYyd/ulPbhbbXqPH2j9Izyq8Dzsw+aHahwf4f0KQvmBYwl0uOIPmbzAh
Uywit6r9tbP6MA2uGUehJ+2rjs4eOvKUh2JU4dpRzuC/0MAZeYzA1yulJyib
S1mDw/RmP5sOdHBh3PHaCtfnfuErG9Kh9SidaXSZgIVOyGjRdBYFEBY11r2/
ZJ3b07BWX+WjgVzMrX1xPg4LxEOUjdzIP5xnFz/+1NrDjWG2a6zEmBZ82hWN
Eb6XQzIvbOMsZb7jYOeXctsW0B2mQF6i+dbitT/BDrLF681zbUk6NTQYheLa
gXfr5tqs5vL1Z8jOpLYSi6aCwv/DYWkl409N/c57Q0l9Nx4LAwuUOROsZnsV
dndVY2Q2Ys7yrQ/N+1QvieOPAKfoaBGJHhXkYJaTlW5FE9PMYYpZvbO8p38j
2mA8R+olkYKAduHWxA9lEGoCtVXJG40jWYnT1yEBoWPLDNBqgB3kzfDbrTB2
1y0dynQ9/XzSgi+/lEHlpVxQJYXiCAcG5mIkYfZYt53pCbZLut0WG3u82Vso
kShhjvFl3XMb4GX+ELjSc3yJGfo4Og6zB+tCkEyBUyMJoW9VsTEIHGhuc2B7
gpErWE3eSScUxTC7g1JiVOyGTYfz6expYITo0u+MIZ2MwEmokdSBj15aov5G
l1W7/PcsFuETsg4ydgoc0c8hobT2Yhxuty6P/EugmUW0QbDntqqbfNmy1/or
90ovTc8olAhZrY2+BVVnHsJJvxHxKck35o9b9lOiZUr3f9hBGKeW4osBRMXB
1EJClMf+g3+YOU6KU3khtK5G53JKlCdxJ+pF0ELEaXjLNQxHPIsFm/50AXQP
LFtrbzu0nFHEeT5y59jZBSOJKDzLvxMaNnDpvtxRnAIgNbpsTCDoWF7W0EIY
vLUYT6D/whaa4RsHlpGcv8eFPEe61Z7mXNGTCcouib7yhTm00KFGU48l1r5l
5lnjs7ZZyTZ9Yc2XWrjTGK/d0u44e1zJurpfGeWdhfgPjpanirLX0Qrh7Iui
QCiN8qHM0UeJJ6+gq98qPZLWSJQ7wJdwYQtg4/C87udPkcXY9qzqyaHB0XWZ
j4Uh7ZhMX9v76gqhbPpLQS4QRtpfU0cK2OfitSahUfTXVWk4uMbxUkPVWFwV
MU8yz1BV8nlPNkm5K+n0dVDYyRzwijVMK3pwTWzExJCzU2Ys4T5poPJX9zMy
BpHiPdpZ65DUYOLoCL2hNfXvwIRRyfvOJ4M25llBVfTSQBpV8Gda+ytqw53b
CukgpHlw7cNT6ByVm7rCkSQQPJvKLt/N928bAS8pBA/XkVoqllp3qSuYIUFK
U6VPgrVK5KT0w++fU0GV2dvHX39XhbUNt89E6tvyOxFmxC8TQqTz3Yo+VGnG
BQXyI8bW+NO7IRmyYi5r7mhq1sL26P6OJmoOfAtd2dXCbl0C3+OZ8QOXdziX
oINpTWPbfL/MEOILscKL8ZIrFJd/6ZSvDR9fNB7Cvslid5iawzjgQ1mZj44L
/+cnJZCehl8VqeTWPjGOyGq7pg1paXgtyjvXqWeCCuOUbsExOy2rFf+WZVqi
3s/w5DzbzLYxYV9awq5FsU9iYpDITR/CXU+aNCZk/cGhlnKf8S7kazKZJT/b
aXAknV6ZlO+bt2O8/fk2YpD2T5JjpVR5BV5fpgTQcPsp3iwAMYhHi82agCFP
tNK7/ZZKZ3PMOxfBhPtGfO1a0qdAW0gtTB9wh9qNSzgyQm+lUqmTATBeMj/9
r4U5/2jxo4o21HMJdCMc4Xt2Gq5yBfFQMMTXiI0wjvR6dCETizuY+q1VHSdo
JiyCV+ZpJMEkeMeqJ1Tc4muqhqKiw2UWA6PL7bLKasFe9FU0r8J7YCC8Q3xg
oB5zPUkoySviT08MgFaenFwydkSOHrekpN7eXxS3tgQRB5v2QWzMZFWsE+V+
+eMNbDCcYdvdsgdDESZp6/jFdPUQ8B2uVn8rKYMxLTusFnkFrjIQvh0FWLev
bF0cJTqtsxLJ6e/MQOxbAfTqAKw/CToZS6P4DVoexa9huIaP5c0HA2f62rbp
OUyb7q6mKaPrYOfzbBmOxxmeyuDNd3xWby2dpoWIwXerras2Pxil7bFIRZfP
zM5aYMmFv+0sTspQmfM0LPPTs8MFV8jQbLXIIfib6BECtmnDKh6xftPD6ADZ
dv9JBxphxVQpnrKYJ/iZ7vPwci+h3IzNZ6fqCKwTS2GL8+dfsVBH8crUxy5V
S0SLNtDz6Q3AH8Yg9Z7SzFXIZTKxyFMqTkKDamCQBCGbz0ugX05XM01Ze6xP
Q0A4HcJMKpHK0jwfabI0ZpZlKgMg83GF2mOxJ1ckSX7bNpQHIva/6uXKYoii
K5MYz3c6jP/1/oadyy23FbAxtzjbANPp9xcvs7O3XTLUTkgeTvulmjyHA0Fv
fl7SvljcZW16VLnYzDLZlDJ+f+s4UQssZSZBMeUEt1JIpHM1D3XVfSLSm62Z
iVyB9JUh/QSOnHCxUfpH4L1Q7CzD8c1SWTNCSq1oApxmBsgBOxFnyPF3j5Q0
pUrZ2Gsir/KqffDFc3iihnP0X5vyMsY99RDbbL/zkwOZawLmozNR9WfXuvVY
K8KeyjX2V2p3HNMjK1ImiVSF0w7aNbKywfixCfJgU1oHkeSLzEZIUmLfe6sG
pf+VShf1z2oojzUdxCFuz7hNWtIHFP4ziywqtQxa42E4hiyewHRYX02HNaFM
RksmNhyrwT8rCfSFgg2cCsdeDyGo8m1fWQ5ImzDGqAiGifYiUXiAjp53kF7H
imOAeW5RTuRXe4NTkKdoztciigyD6EJWScuJi93C6xCehHINVQ3n0KH8avcx
RoKxGyHeGFvZ7hHSindLta804iGLJtyesTB6s1r+SX6cBqpfuga0dlFMSmwZ
28kfzViZC12NSzAsKWkBaxZl2Mi91rQ1gkZ5HVf/4H6VnsO7kFY4aJzABBmP
OaLD3/egjylujrbwf1fMem+Z0TxWudj1bBloxjK1CeUxIPn3a1qOvehAG/Hl
cE7/mqqeHv0eeVtQ07BXDLvpuyyS+ARbWOWpifUwVmEgJAV7I+VQzTkpFv8r
yRQNThp1W/DaaeT/YSlSn3EDUAKxryfYYBw3hK3tjaUyiBTP+vGTUqLKfTnh
KnbdwJHMHW8ZsMRc1Ykea1SrK9E9wQho45skeT1augjFy2mG4Q1jslWOCjOE
5pExu9LSINnSpbMV9EJVmHekekcbuJFEHbIvT5rBypVAd7ndLEPNmIdYTERG
QxuitDxcVAtioLMgH7RdGUKE+aXZ8NA1Gq7dMYit5sChp7X4HVCWPUMnwylr
n4kfM6oq2ru4504Kp0Ahho4+Giuhlm2I2lqalrbfKXr8VQUktfot0WCdj4DB
Hhf3UKOaNbhCNQrA0rUjTA25IHkpWSb5XTzADj1qaJZBa9CctSsuAo4tJgF1
T+2lcR3STUGFzYBU9iY76PRJSZ5g3g53HWAEZrCrIvNAWUgbQRMfkAHwMV/f
jqjYLFhUuhLtvdSMarADdPOgPlLr6ri+phU8mjY9yCUb4s1K+bPVIi0Xomlv
a09KVIdIgQMp0/Cx2t45anr5Z77iTYhnxZ0B6KV6NcK1rSkkW0/myLn16D0v
0ZJlRqIwd70nxYcL7n4zX7dDRw9jyASC1ZXXZGbssehNKwya3QryO+VvLP6L
Y9yotXAxRlN2hH0x7o9TRbNAd1MzZtSA6DnWnNTO68n8NYwkn4TxprijNLxM
K38q+NDQUU7uGbS5vvFC7l8OsSf3x4tL3tEkoBdbag4ZFUPbc0nJ6vCioOat
JTsezBvrAXoaACxH6piJKjvWjPJkLp+rLuWUq/zSuuDljgDBSG8Br+5cBl8D
RH1od4L7ubKQC5lryOVCjtOkugGTtsEeqMZSpBDZ9EYSaLFmlfm/hT/VEtlU
3Jt1pBJXkUTxNkjhz6KDpIv2qYxrSvXcT5jkKDRROP+BZFtFl1KV+5UuBs1e
2HswQ22ELn0M7AAFxViqxodlrwSS36U/hwEBTPwMQUsBSbMdIyKAEuM98+WJ
ToGkQATBO3/u0DBxGfXhwzLgceOPnW1I+zgtHmVduZ5nlOhaY+tQg34oxyZ6
hVJB9N76iWECPgmZMYOLKshQ++2yTX6ekB8whxb4PXWYf9I0MA6hPDedu+ZT
JUjDBGSYnvb26thY3EQK6J11e+d6JvzXNmeBffPBda+1r0JQuFu3Wd3YE//y
tEDtf/rK0HlVBV9iwFezU90r4Kh+F46TTfsjV4YhE9X+upHWobybdJ9QoNJ8
v+4L+IWlHKimx0dIf9Eo6mTLldImEb5RMSsVZz/8M413BIivbwriuhgHid+F
45gwdHWtCIucOsLiS7qQyA8eGlADw+VEpR6JD8QMaUP5BVt+d33poN8U14L8
kIVchSvOCdMO9gsfLNqsFw2LvGX/lepVCve7EmX59Zyy7KTfechssGGWr2t4
t9EuP4HJTwamxRkdA9H1+DYSKLQyh4/g2wFWS3lJgXO6HZ2YnyasCGORnVXy
HGgz/3+z0HVMurY0ESuuDtcd7jfW3iKoAO13a50l0oq9mSO4BCIb1IFRb89F
GUXnbcUCoGqdFF2qR6cvbHUb2N/IOLxPXL9XNkM3olT/KxTW9nzfyRQ9d/Ph
cMhbuxoVTxAG8wRLk3xNRaIXHevClIkGM5W60dxmcaq5gRHk7krsvxm8VYWi
yGfd1NWg65RqcKvjFrumEuchfO0l5y9hwfgziPtMF8kDdQFm303Un28BTeU+
pCxwOL1JUs5e5OxHQQB8tkU8A3kxUuOjcOKz/KOvv8C/Wz6zqMe03GUa83p0
078EH6+xvaBIwJeBu6NywXPVmxqv00MVOwXmKT68jjvwIJ1x+suZrAOZHMHa
u1NmHX4ElvBx+TheaqXIEIf3wYokn+jYousIVUa4nUQwxbo+/l5CYrPsVwCU
QpzCILrDwyXL465ryX+0k49DyhG1lhhsA5IxKroQstZQ9BlCtbrdiOqwE4RD
f6u1ZhTw+sk+Ulrse5PW+hor5ED3rH8ckp3Lyyie3kC0jTfRPQGm8Pc44m5U
yyPxApJw/C4HjoOyCrjl3S6OqY5jc9+VVa/iIeWwXk+HaZhquhCmEmhZb90V
TAQBFxT6+i3r/22Kyy87/SWHCrO/gh8tzDh1yM6QghT1+BRtfLzU8Fj4Iya6
rE7aXRhGK0WyH6hvQiOZEEF9ROSeIMXSO+sI9qR8Ps06UFhrFnTw4OBl7/EY
31LJrbqUsuLUeW5FsqzLz6+NgvBnHj4K+2T1/1d7VRIvG/bkd6mfwmEHo7lD
i01lXcHbXt3fxd/AXJWKXtwDETLjbBv8uJmB7BBnhcJjsVhP6IpilPAPAosZ
cOMDAhxZ1Cha4CQB8ptox6/HPRRWlKsEsaDpPIINyeAw39TmQtlISwhjMK2g
59TOCiEua87akYysAMAyCF+knYd13QN7igW9whjzjDQZhwve33dshn4g7jMD
WRHGyX2U/MNwF7ACweMBk7ootfgxHLR2cWPHTQQTNqCH7m9cFW6QjzukQIOa
9QeNQa00DMf4Y/BPRQz405KXOIRw/HwZgUx9gu/4IBI1+B7dpX0SlnCmSrdl
pQbjKDOuXyQwnTz2JUVM5u3LJxP9OXN0CDlilYIwfIHgiIKS5/HTjK/KByE1
WYXe2KalH1KTe+gvemiTgU72W/ZvE3KEVKMIsapEaxXBqjHLuAABG1GDhr4D
MFvTvJbwV9XMJwGx0UOOJ2GbNtFQz4iOGANCekKUyoJ/sBvISa7+urys/8o+
WkzWGbbHU6XKHtHgYjskhv7RNaBtc/K7TZRutTYNOL3V42xempmGnmPD6teh
d7K0qqcLwPnQx4bTYs10A6URcrfkfSc6elnhGSvKR2YBpl1DOoSqCJOa02ut
gHsKW5D4PYI03HRStY6KW07+MMz8qXfdGaruXlGgRfu62+MU1wF6eXiFHmMg
2pd6Z0POOBTzzxDlOxanFAcudYT7SX+fpkoD7FkfCz11IuNkZ4Vw5Zh0UvRD
CapR0pDicfIdm09aD8U4Bq+o/APrL4CLkXalwg20KJLouhqItpz0AwoN6T7e
zTZBB4vzykfIbAoEcKFNW+0fNX0NajYIXxlLaom9y8n/BAD8UGcqsoZsfgcS
709blrOHVHmQithWk8jahgBPe/xLbnt4iUDy4gGYxmrA+nUP8NJLwYGZi9bO
YssvjuTcjlqOq1gwsCx+cblZwInJidhO/41vjBdZ4cBk+YLp2LqZW3KV5s/4
+77lVXYhxpwBh6Riik/HGCA8FXzeQFjL6LwAmmsfEI7QyZX18/nAb3R5FpiH
Qi4GURnw1en2Qr9e+DNSvQbP5n2UrMVGdlVrZhbPeqPj/Sshrn8TkSUfvW+d
sNcfWtdRIIf7mAdeE5MeuDE7rukZY/cQeKPrGExAeVjeen56mODfl8pmQRJV
sKhY3eLsSf6RHAVnItDVVMODVo75B2TrXk3iFhON6rjObR2EYU7Xibz9nhve
20+jnqlRGlYnvl1hZvjny/Qr/FGgSB/4rOUhWl9u0CdiFgaqX+t5xhd41ePA
eOHAN7OpBlKg1GItdjdldayA4wwA2ywvm6kjRovrv86blELbX4WCcVxR/DxC
wyJfqKI800qJNefvVkpzCEk7sQdeL8N+/2/X1sQjNrG1zbxD3yFsfeJ3QLBS
t4z/gVieTHZQY2cw/F5G46buQAtTAGWBfmQ6OKyP7lTTfoCyrbN9V6zpEgCg
1JEdiMONuIpB++MXQdBzUanl4Rm54FcFwqAVlrUBxFgMekRo6PfrYvBbAih+
oHfsJ8Ppx5s0GWrTYuAZWNpArhkEFN8YguhJXKMQ3s+7eyc0LfnPjsg4y0yu
mxzPCAnmELRhk/XNwJ4ShLDAmHWhOzH4EdGVmcVoBIvGsJEXHECq1vS0eSoH
TmbflMUI9hI5SKBXieWtyrwnIDekJ23hPmSR9Ana/3eO+h3qZXksddaBG1YV
PvSh/L56EXU++8Fzyn9lBgcuMddDA7xSPXm5kqAR29AfFHXXK/NeYXWDl8tw
z25vpht5Pd4TbRYkoX2jZvtIT1oLmYrccXJN7GleSzY0xJmF2GejwjHxk+fG
esURwiwM65gx7z/a8H3aucePTBfYvgvQIC5c5v2SQJv6dLapDbZfzyJf2fsA
ENkneokjufwla3wDaF+dOonSkpxXZXx96aMgIK5+KkPkhayONlWYR/7LONul
1x5nLMQAC5NlLS4W4jPKBfxe8pznwdpDm1O/iTytsXQbx04yoBwMhqhEOLZ2
oNrmhRgkEBkRjFsXFKjw+FBD82Tzq2lrYgvpf4cOdfKCEKR7T8kglgr8dM7F
sGrO+QIG9SjNXUvc+A/VsiPqykuw113jcZ65/wE5OFHUmR4wdrM0BYnvuDFO
QeYw+MkxK6i2iQF9wXzNy4VWTa9aOvL2ZwqvZyf48+3xkYATyZKyBfFDXkUd
h+4+XVEKGTObCP8q78IQMQRNc9LP1SSDRlDUwNXpA0wZ6qHVP+xqK10R776P
HvB5d6BWbSLXXfiU/FenI5KhoiKEHdKQFSToDOl3xpQp+KVIYvX5QYISmbuS
H1UTr7Mm1bKOkYJo8Urk/bFvJlPtmfCVU9KK6amEDR284qwsBNIUzDWNl2+/
se3h6m8ELluKYVp6qWc+ddazGTcd7BiXIXYUc60e6AVJYS78gtNBvSFrU8yG
GN4viLHMQuD/mj1KyioC0AKjWJFTiP3S2XUY6Rpb288CL4IqSzSnBzyNke3z
Rj0z00eRx1RjJghNBY3VkX2KBjp9QdBSCsk3MJ8JcZF/aETRuapneKYm4ykc
64dMhsKYyzHm6By0Pk47JUUBkd45IwUZbKF3HY5798A35XYI688KngNltP/k
b18eTb65h9mMdS78WbbS7c+l8PvLvv2V+QGeUcPULp2dTX37kx2d5ULF+tct
nHK/Gyvht1Y17Ia1ItkLD0DfghEYXsEQrt5g10vbURpfkJ44GLdDP247hkDp
n0tP6VUQ2K+YQJKuryNDzp8EGl4sUfDMfdeqHCTJOkaNlP5Bndo9bTNJNIOe
5P+eQkcw6c4qG18xGNT+GMsEssnGwApgE3ExvKMcKSTOYXAyUSWr9mT9eoV4
pzV6iE94OJVYn+ri+Iit1XXh6ME/TLxhmFpaAv5tAiIRjNPGOlsrvrtRWV9z
ZxSuZfiiB2vm1QD1qZJ3XzBWopcoxnPwyuC+BuDmCjXIKnv0uI4u159w56ku
nS8g1SH4f8De5lQKBk1LWG2fEJyRTWlXTtCsfz4nLmQgpHFd016RB1ZbjTxE
coeWI/9LD6f7KPYkrspDdkQ/WcdPb5SCr/5V07mFB+YjdG8Z8LaX5gFWVS9s
4nmYY8EdDSs29+R+Q/Z4NrIhh/W1qnsmunu22VIXQBcMvabe+vRqAx87h/2k
F1ZsHDnAUI9IohysH/Ra3iSp/W+qM0YbahEL5Dtsmj/viOs7gnXJrsXazfwU
NrrwLHocHpfM2AA0kteoZ9IZzmzoQ2rB38lO/+if4amrbNyu+aPczIem7h0G
2lRTV3Sq895NTPDZa4O/wsYnT08/hWKG6ArccWLs1akjPayYOAvXTh7LuaIE
3YMjhuSwDEWpFVgK/m73qp+A4XTkfkf2cZEbRhXJbLFjUVYGsJHg2PlOH2H5
TK7cp/i9404qRAvx7aK7P4fS4MD5nwmgSXVB+uCwTwkxcvpUv58OYddcWfCk
sjvCNAUtU4EeBdQBUKhic+n7036r06r+VCOQ4X06gmzNM1b/UsKFvoi+N+aU
ZJ86fZY9ma+GIqQAjwV4WctQc3vZKlebC+dgWyOZ9QfahL8DJTGlmZXnTE2e
xrBdELQAKiNwGQmeQ20jNrUjbzWmoDgBur7AyqjLECmCbV9K7VK5G0GRn9IX
m/mEuIwZi9FlK3+JMEHhpmWTCd95xm3JfoksjvcjngUT8toEwJ/Dhqc0Veny
A1kJpUpsHrRtZWYc8HtM5qsRvMXlp6xwn8SclJ8zCiWc5PiZ1ab9ESfzBymB
DbnljFSStI3Rlfx33V+VbR+Ig1d/o1SExXnKvue+lZxGDIMvEzKvUNdSPnO0
WQvt4FHj0rELe71x3dVEssJDTUc9IaMP+HLHe9pB1rZrr4PE0dKBxOnOyxYL
dlQcP+VT0KPjn9y2IfhxSRAk+z/FvSp9VekY93BEFmfhpk8Zdlcg3VEnxalE
fRb8Um6RiwIWsnIbzPSMEL1xf8rizwB7TgKa/ytWlncQzpLUXLN3EUIGdAHX
7ptsQ+7XGsNSj0dUsOzOyhkEJS2pflFWGY+qeX0Xi+S2KfmHB5fWQeRynMy1
AeYryW0Zph0qfPPd2NzjjTyCQmYScQlKM4wlw30+VfhCK1V+D2Dli6L9cwuU
Fy43EDC+Njlgk9RT3E36eghLBzkeAiUoh3bHzXzvXmWZuoDTUPLQ2EtZ3qwf
zlBWJ++4qaq+qmTRMBgrsQ0JF8Iy3cE4L4GL3O40DyCQMchAXKF12CfAk3bS
sx4n0myYPSgsLjwJ27InGWPQb/9/applXgJH8t0bKQGBSJdItXfVVODg8bBA
J70PNg6fBCJCr1jcuw+pSfJoUgKoKYcQyRO/2XyGh8umEAJ1WEJDYlha7cym
kRwJA1gK9AshGoYeODzTnW52daIcXzq2KnGrx5nH33beL5ikuBB26Ng3J77/
SEiNwh5SepJGrB065ELe0q76QVj/j+O/HEE4OUPC6iE/j9E8vi1yvt00LNTW
7xrRrQ5L0PWLo7u8ZlykbTgD7FSDD8oCQYOvf+IxBcLb4w/L8uR6pXPZWB42
kcWJZeaXItcHLvG8pzRERUhepgWtU++jdTydbz98oKLmS7sBCsoo4Br2usW1
66kS2PS+CgFQqI3SRyFwx8DD97cAatoz8BqeUCmd08uL54HVQTnQvF4h+sLo
bNONrtJ4/mcDZ57zFJdJKX1wXzrcf12ok0X1QwTpixhZvVEraCKnstgcnPZV
MQ8nvzusWlGOBIpccQE06Bkg60nIlXI0jNozAYHitI+EWjo7ayFIwfVoS8dI
Aa7A5n0lB9EeOZrSGOzFSBzbwLurvFDRZC6/o1HA+EVOEHKONepd5otikI1J
Su7SZFvzK7liVR/KX5G0+MxsU/M7HODQ4P4UWT2w1mqzTlazr9T5f4aMRrnh
raLIpCzsQYV7skcf5BOovcCybQG8pQSY38qyPoG00OyY1WLYbV2nQht4w0ft
9TRvWAf1y3IfFYQ5q2IFA0QITQ7htGD9cXJwCdO49z6owu4kXa/Hj44vMoMz
jWmCZYKNJGlmXMvvTgZ8k5ehhqKElvLo/NiDKCm02u5BY7yuDdfWBMg85hVi
Gd636AwfI1R/P4TMMykRNrzdMH8Qz3BD5bUjmzPm+og4XRsWC55Jy+rGZVBc
QPTJaXS/iuS9hw1ZNFZzZ/85VVt/H6rvKJpYPZ95AYA8Rxp5NLt8ptnIrC0Z
7rwNXcxU2gTa33BtCmoQPmmeCvlrgMEbWE33aKJOzGiCCxYxv24NnVXxLbaW
ci4Y2hek1QwBwZ2osoVrjgM/FJsz6z6+1cz5pRUoJ31VWwQq3il/zvMeQqEs
Pa8rC/7zcN5JJK9M12Wn7mR6q5+QhNY9onmfjeqhJp7R2+8xSgee770GiV5i
nhrJVsbicklGs2AUkUP4vYK8FdqM/4Xu1LmLpViT8bxldcqznmTSFNKPpW5h
OBIjm0B2oPU8BiK+j0hR7W0+ui6BWb3tV4vXl0dmi+P8Iiu/lQLAEBO/3LPo
WR6IkhzqPd09Nm1zce9y0faFYcXMueBd2C/OIcZYKkzoI4vCmD/91nO9TuY7
p9oFycBjkbhI48xJgWII7zmE9RCMzzJv1kQd+PmR3efbu+IsWXHZwVTxV6BF
Xvs7svWU69aNvKUpfx8ztMeSE5WroGNv2MNFb4XmZkD2EOEwr40b+/wKvazd
AzxoLLkRNgh4itITMFAGN3YsApy6nea3Olg+kTu3hKWnAyHSG88UfwcDsouq
jkoDaZPNMmnycEXIwr8fPRm0G7RaRxPMkksAh7peNt2ytnsFXX9w94QGZhki
0Xp2n1cbT2CwAPVZYJvO6ca9WhM/3HXRvOAJBDi7AEVarULPzQzRqVNDoRm6
8kZ9ckVI5axm8ZzmdpADboFtBieCJ0QjmZpgw/1whTSi+KNq2V2hFxttYkhP
D6cIkaNuXfZLRAk6B0n9PRcF0x8ocYLi54ovOFaQ0Z9Xh8JkCtuy7fMSHRtJ
r4QGGbQEhA+kVC90MgXp4l6o8lnJeJjWVmTDGO0h/xwgIYjsJ/Maj34gwqKh
Inolq9eYH4OgPTWSrYMLmeqqWBKdFlw/k6rYGkZN1/2Qq9xJAW65K46x4pHJ
+OUxYVtRCEzdX300oitVbJ0kASvzqDv5/9dcmsLu//lBJEw5jTt+YUEIzb8K
6kgcpUMyCI18FDLMvL/6nq1nkHLIElrPmQ1judc8deNsuxcfXwNtJMM8nAmf
+cYi5cqGbLeBmyJwrjg7K72HgsLi99oxqW2gBq0nK+x0tOInwTjohJvSpVKC
hBhaDLYn4qui2bEPKOThw2XTUIn72UyfPktPfMvMItyjrNFOOwznk1TqEvM5
ogUznAmBCwmeI0wC+iqMnfmR6daZ8Esy1ApKKreO9WSFarVrJkWS/HK7i7tM
rBSSBE7j4rfLWUAXHXQHuxSawtkq5OFyue+0RRyVp2voVq3wrTAKaaiS1hqY
M6UUf5I+PO6TULDLba+zIP/vD1xWyf0MBVvv4w9iqPNeOfWKJIjmWorAK5Eb
Nnu+s0dokbEURbCCYFk0F+3Jfb/3y0F170rANCmkSdxCYHd2JLo3+FeK0xXq
NiiBroVds5S7BVm6K5uJRRTM1IPlFau3Zx4wrnY2V7CSTYjCBaQKlkjsp9YL
GpHDhNAsjzHFSYqimLXGnLynXbMoAFT8rifziv8gy7bu1fo7+URdAZOLPoyt
DeJLD7jGOdtEXxZIqtSFH9flVAYI/vO09epn1Q9aVEujpm3OzNOq7K6o2UQ0
YavfWrbBwvRrPJKqgXEGbF+shYBHa0raT02ZJUYSUIq/wMqXKK+JzXWPLWlR
J2FHN26/K6lVLXGw4qdY7xT61e4Vjlx4KBOXTxmfYJOS8q/653WsVF+HA4EP
AX8UUDPAK9sx2f/NVcVBL/BjoUjqvruhKRqoIZ0zJkPKXlSRqBfGiqrmO9GQ
mz8j6iJgv3dqhHSW0cG2L1SmEksVxkWHGDPFEffgnzQBPuL5xYmFCOzBzIY8
m6J2AAxA92ru6K53Cxvh7snPpnKH3YEp8cDaqwttup4tpi7x6JDJNCoWGEt7
0gZSlXVqAP3RktEaFRj861n8a9SnRc77CxQOcG/fIoVFIwMf9Bj4ZFz+RkX/
tr3Zpyng85veDKXG/LzzxEwDL7acrlo+ehFa0XV+7VHi4JX78XmP8Sc8Kc2r
AyPgxTH4eicn9EICJWhdPrXm5wEZUvYxapuuf2Xy1qqnCJESAEGs0R/m5pi1
DVEPuVpsCaOyaA1kNzrs7qSv70opoC7tc0I30UCAyert7W8mEhPCU9ZP4EJb
o/fH8xKxUPTL8x8plkBuOOMf753daSIgQry4GQklYkoVR2LcL13vHapOEvCF
Xxl9d1yWE1bfFisNGECxuP39o96m6k00VEVh0Ygh6vD+qa+EOZM2VG0nXkuv
Htk5n6aZufl9/MUJi/WERENzyfFzKaIQRr7033AmnLBFn2WZmHS8F7vi6aTQ
yaO06sLHsBukbpgnkadjOdjfYBCWVqepHKmqCNW1/otakWkNaK1YQdosQtth
wBJRg4le3waUFdRRrrlBsAoRJaAvzc3oirL7lyN3CdzAYwbAjypbMvWVb+Dn
m9Z00TAqmuD10FzjMsM4Qjq4oOjD/oabUmIPI82yqMIT5JioDI7iCRkzujvs
y/GraG/dwTgD71cuNNNy5gMHMlXGVWesXwdZQz3Wn00gz7t4gRgklTH4IuJT
2x1/U9mMv9cMcD6Qhc4ycShYaR7v4A7QwJvr2kXnLAnOjym1y1XQ9kwJBxtV
38g9mOz8MiJ3pvaczQ2BPDibjHc40anvkame4xIwC84rGrI5T1HIlQ1+AOOo
iJPAe5s0Lgtu4yxf0E/7fDB5W16vEhItO1KV4Vjo/xCYKuE1hCi+jG78auKv
WtxOFGqlWkqvcgYgTI+PqfFk7PNj763jVzUF7PDHTWBEUB1exIor4PUyaI46
wUTg3HKr2PweaDvv/lxxvb0n15Rdh0vV883Q6VhO/FIPac6WWCBJ5r8nIagz
rELmx3BgCeIuFog7pMWJyLcdtEkSXWI87yAHynymatzzKY13H23a23OogcJ3
hKRQq/wf2hkZcgVlgdnqoK4/IU/mTJd7g+tuos1GnZ6ykrgBa2gJEdOMe5rT
gSKJn/2wHLM0U+6+s6IvjPGQsQHbwlTolAQXqP2v+RtUmPMQU50I6iRZ4H0a
0UuvyH9IhbDlDJ9RJ0xKQ4UFpabQnSBxj9tX6MMqJbtdWLflr8yTcKalUGkY
ISvtCP66+QSkC+Kbo7IRcaxA4QlEYpIhIBZ75GMjbRSBA5460zBZN933K+sm
OIgVEQ8BDZbKQehBR7Z6aCJ8ZtTM9Tjk2LOAnuWEclTN9MB42wYTCLGXm74o
iliNz32C9Nnt1jXQp8BctOCvVcG1/lrp8yNPpO//85kfO6qYyreit1FwJ3Bq
gT0FWN4UWzvkJcy68yqdbNtkCr79jeF9JvEoZyAx/DsFeuuQy0g+2d6IwjCK
Pdp4reaxMs15JqCuqtMctXeBe1Rw6AirX4mupBgjuDz7N/t+Z2Yz8q4OtC63
NsP4s1HGlrSCqWcY8t+FL9JKnyJHEvECk9q7Nqtn/btZMdk6RV3mQMCLLJ/E
244TzsjtTj3Hlj/zxeTHdfqMbCaMF0gjpwXJCsyw4x9tfI7VZhMw7VN8Qlmc
hxuoWB0OMk/Zy3PI23QApW1jHjuvDr7cYWRKUbbvL/sbNtqKYSYTZRnJ6hAy
VM9CBvSVBzsgcmAFyslAwCuYePhmxWNJumj+sQcKKZXriMmm0Pc1eK77D34e
7fG0BrvDy4Qc7RqFB2HwxINaCHp0tvJHdgqHmWr21JxNXxsO2EWYDFEXFHa+
GOr7MBOxRoyRgZSdDo/D3HTobmm5jmxGn/2CI3MPlH6oShmGmcUjjKjJ+GAQ
ruKn2uOukvpOJqZbZ1KFfiN3iGBsrZEUHBg2+wtw3v4v/s7nmMEzQl7dZ4HD
5M3x4ahVw4IIilxHOY57oLz3FvoTYe82EPGIqiXztdJv94yW18tEmIZZUOf/
jwfGuTBn6xDg+DtrFOpm2CyZ6zUoY9Gyxd1Sd3bfTj4fF8B0wdIXdXiNA09k
vmgWSd+G4NsxgwmQTQhDR+52+MiPehNJf2Ct9izkUJYH502YWYIqWO4vvo8P
4EIPU2jK9CFoA8tiEp4efxHJ52pBTn9UWg2byEUUiYpxpGAJ+SQ7+vQp6Gwi
MnFvJoNgKMv4BdjES/lQcLCOQam6GPXPu0585iYypRrfhqpQXkfa2wDIDi7s
EqZL5T4uQenm+Cdc35Z63b4UqujBbRrfZas5kWH+/voUFPyCcdYAnYk2dUwP
e2YRYsxVfnK69+UWU1ysS79jknoYGzWA33k/x6yviIb9HW+bhi2l2DujiWwH
RA10oA/xekeacbmehcYhncmBKdGTlZ22J0NWkxaXnlomyubG6uGiGcV7BVGp
ylP0FTtKJu2EDZilKO+bvUGLGZcOG6Bp66MtONq0X8JSW+OSZgBzYm18eUVq
EXKIHeETo28S9lqnHkkkisJUCY4UX7+0P2GDWx2TnfTjVMxZUKV9GkS8jzxQ
VjxVW24s2jrzahrud6yv6WwB0+RaYUZxkWLI/EVau2vDsQPoBq30RIJRm9B5
Sojvw2gvz2BOOXMyTpSxQaZYfIRNxpyn1HW6+64TcuZcfgqVUOkcAXAStYsm
WhyYM/YC0zWBsXtv9UHQMYpdZK4Xm7Etju2MaHZMpVvS444Qk2DCRlSwZIJl
3OYFpE4AeYdBEWjMA5EfBNn6uUuYoh0S4CgRSYVS10j+m64/1mLvLg2Rvagl
mJDi10OsixfKkpMN6QQZ3s2259g6c4KDWZvUFOqXFrzg8oJPpNO2xEMBoLDU
+6DFTydctQ+agLLRrkqeNq4hCDhZmYUKSIMmHRvDa78djAxYTnakKn51en5D
OGOLmDwXzuYX5krHm2SVnCB43ZwwTk40YZ2ZaKA+wz0VeG1YIEXvrOYsmKih
fLHpOvxMwIpBm7yUYo25o5n/1TW1ZxX3JEUXs9y6QD0ZOLfZMJwbFQVXs8MK
hONeUSFh5mbyCJeUC86SfAvwdMyYLvp3uvjofeFwz2EUA6z5moCSeoKWl6jy
vZkeFaedAtwjgMXdDaTkh1Skdv1eGrFyrrxvsKliY0SZMBVjaKoBjbZaXESD
2oiaErl/qAjEn1L2wgZNIoLrDheF1BjnggitpfzenJ9c32mCjeKZxgDLYg9k
2NKhR9YOCGIZ7V5DU7PzDB/NBhfPZPlkn/OqGluvmtpDQgzo2vH+HGVBZr0n
Ix5Atr4UWoXAreTFXhIaLM6OckjdCycvr+croip2RinlZWOSlYbdNBeGmF4Q
90M/x6DNfdMkvYr63WyJSGbb+wnScZxiPffwaSYRB1iTyYbWKcY0kf5Yz1eg
FG0QCeXGFIsUEtsyRnKJUhOBN+D/0UZfpVpRvEqHYGcRanDNKSX23yNQ337v
aoJnXAAeuBEduEc60FjStpxcfSgbAjfmS2cgJ+ulfwtwnDraPtFRaReUi6yd
M004Of7AZ6akw0hjWRUrdgiaASH7PIRO62lxy9XBPMvOcNHTlBPHgSciMI0K
xWVzIsYVEFTr9ThWYzLoSHC1cy7Z1drBODfBTioQwmqH+K93ADJ6KzJBe5lq
TBRs7s/6PwYrxlwugL2baWTbpCY6MOFXemsDsUfy44yjBg97cusMp4J5M76Z
PBUUAEjaf7MrIxKKY6WfM3j/TVOZXD4RbXAfuqDVgE2VfSw+ANJ5XvIMhMH6
fdFAg4jn9FRmhPvy+LMryO3TMg/vRoQnqG8HyDsvZruhYkR2ehgYTL8pU5Bp
v23HGGiBmiU9rpzGFqr8WoeKJlVT7+G+jRZOPrqXo8zPNKvsrZarg2zsWHxt
pgPJPmY1dN3Z0KxWtggTodqTVs/I4RPSb2IsqK/MmjMBwOHfmcmPvwU2fFK5
CEdkLPKgxMXG1oy51qmriAJ7iEOx0bWI1V12Ty4/QDu2SnQ13cuCXPGbB5ta
GbDS66pIwlPhNSTm/JzCbi/zmK5cPEoCwABgiFg2pGGz9R1DVCpp8PS+dhoE
R0bo3rVi4oilqsOeqMRjNxkOpGPrbWgeEGwnkO/YGuJJVEPTHA2yiLkiEBPv
rqWup74ysm2MnAQyvV4CEfrnHhvo5G/dxNmfmQXTdst5xKoknXY4svgmyEg+
dp5vi9B4Yn4nGwi6Z3rnh/bV4S1Ungz+LGR1hiAYBJR4Xc9pDqHSLEpGAMBF
aRo1dxU43q8pk3zCvoK8Vo9nEDFcTIFkpNlDBWxitN4IhPBHB1nf83TpfY/J
sJnPVQZPLO2lBaa1Ig7ABSfJAjJ6DiQ/4R/5h9b6+waroJob+Jp7vaHQKzxt
beiNShp7zzDR7HXhwvbWYojnalTS0L0QYKHTx15sbegB7cvb4NQ/C9HsDSkv
3jXqVhDtwft+pjIM++E9V3tLg9z1drUnHea2zV55SKLjJZ1BbSgcpElxUbkG
S9vPaifusLTTsj8+5jZPqRZtZQBKbh3FQbCvLbtRhqO6KL5KvFZRxfHoxncM
IFUX+ZPHQUum6SHfE2W+zGTD/tKLRDNTzjiLNI+ZRqRrL7Nhk8Vqu/AXA741
69nvR0YFVNeGgkalsMAkupmCIiaDeKw6+wZh1wnIjE3M99DG2UufjlhTrisX
2p5ByoxMCDxq4IZ640RO6oD0/Uu2Lrzg3dnYJREPIQ+vj5gMXLdSiFUXOO1W
f3YoALGvtTFnj/VjlxR6g3gsT1iNUKIXTvotQHxks6Bck0t888eSy5UtdKXU
hJi5dlwkT9Lp1SR7OETVG1v9hkhewV+C3qDfbOw7EBSag/ldSNObI2ITS11m
/OUlsRP11eVq95K3pbEgdoi9W+109C13etb6p0M6AKVQ4IJhC4VvH86Ted73
VfRXU8yxJKFZLLRCJrOqoa5qTeOaIVHHlYdX7PXA7E8p2+2i7CmWmeyLy3/i
cV70Wkx0PQfN90DN90aPimfgLc6P8gcqyFqqaId4MhJmxReNv4huCdHK9oYX
pDZqgL0GGTgjhcxE6vNnYSgwCoA94hrN/oh+r/8VAtjdiWSp/5gTMVo49zqZ
NXcNBxgYEANz8QqBGg16ov0IYJlfZVnn0U1gvA8n0Lk5/V3vkRs8rOo6Io09
mRL1lITkwyZP4ryE2fYrtmJcIpb/wGizZoStQNBNkZo/caQo9xPRj+IG1r9H
Dw36OFoSFzNf23rJkngR5OQj5NU5ko/4rZbWlHwdnh4/M+K0NeFznjIip2P3
Mvhyr6ZOcDt8WveeevoM1Z5CBcgOmX7WCMl7+u6eT0TCvPzqV9hSHJdQFVP1
vNPIW0/gXOvREUHqlzcuyXzYuyxkCsVQKWLO9EixcDbpeYffhe4fjMBF059X
bsNNTuSxhAAVa7aViTvMHCNeuR4PRi4GJHL9CcTcKZBq4tSDdnEXdjykZfXq
n7aMimh+spQTmJUq7KK8e0tIsZiZFiz178p9jRckWSihj2yS0JX10ltXdOlp
voCWoPKBzQfPfMse7bJLbjy1QSM/N2qzj65p4Vjl+Bg0ULBTqiAj/QHc5BbR
OG8T9VoyIsn5x4sZ0ax8pTCiR2M7UlF41ZMgbU3qhGs+4EjONTOgIFL7CIHd
wsPW6vBTPOtVoLvUqyU1SHPg+xpAZ2vgvSadeXektqAFpLF5TuYYP/+cRcni
+9ARdS+WBFfuyEDzF4+CQxo1U6ftYCbapj4sHZrpkpr8NaFrqkLt1bIjV9i/
7crG+d8E1XnsaTKwodQo3zjex0ZZA0lYPwh17bnFSJ4PJETKjlfFCwclkSE1
M4qe+c7kcCWjsNXgRr/ajR1kg1nQRuCjU73VnxQKjdNw5aGfZdFiMIdoTvYk
RciVj6azskHlweA4V/7odwk8LQ3uR5cnvdp+nop43srBI+FxKy7fsN319XbW
BMEhKS6aFfVctzC4lsG9bhCqiFv2fqanSpjNDTXyq7eYrFxINbQYJIbfQeUE
bQ9AJENEgWnV4G86FZfP8ralOCiwfOCwrhlLORyy1MTUSIR3xNWsvzakVhzc
jWJoQjOVxNNU0Qc+X7powqU1xf1CYXetwJBehD5IkBxtppdc2mXPSDVhECsV
sfco8tiUbeTorrCBu/FP5Eu62S6SCZNjpscokknEMFk+qWg1EVLl1xvtachD
i+g4YOjNXkszrhwwhEAruv+RUZByRC8lgfC5ZWVg0PAbhyqbr7mlKgZiwl7q
khnanAd+UxL+FhIFaaGTT5CejENNyTc+WmuJJ9H4qXdRwPwiiHOT94YjyTCA
QsQcc9YSttpCpUbOVJblI6honwbY0co4iervRZyvoBPAXwvMQbBoJoHk8CEA
c9lor9JNBOES6GwUhk3t9ZgLpiJ+9uF8JEbCRa+k005NbZVdyC7AIacEFtpj
jV0w2AHFVMVNoC13LUFOgQgiWVDDjPWrPple9hLGxoJEPUgdCwItYRW/FvZr
F4qkzJJR/Eoe8lYLJLJ13Dnq17v5RC93fzc/NN5X8LHEZdZlL7VNBIobe/ZA
B1IOVjJgbDH0mrE6kIOTvhyyz7ZdKL35qMnIGsCMyHGh0zZPowjzdEIrppLU
7ApgN7Zpd3t6qVJZ5vL1FMhMK1q/nlQL65HEdw3STwGj6DSyxShHR21mZbLv
vbPv2S//folFIN0SsegOx3pNe2Lgm9nwN73jrfHMO/CxIthZl7hYejQKOXka
T+9mOpPjIjcbjkUnhVba6bH0hf4XQ47Ufn2ngoRfS+BPN4BobEtB8Ef0kAbV
YUarCh80xjeShL3w/lmK99lbS2340jDXc5dQZHmUVRPYlkjCWHiZG6rTEKhf
6QJ2DADdkyRoGb50O20zwwLIfq47hrPCmOfMuRf6V9FWdFcNh0xquVJwUSoG
nVVuqTN/qucf3jWeyfSKNI+zx1TC27WtbXSe528sbRZEF3z+Be6vEFH3d5Sb
Z5lttblIyAeIGDDymXyShsP4/ZfeFQ3kGyNb2iLWoleu8KgAugolBRRZ/NLq
Nsz1BQaJBfTIcoAA7y0um6K6c/h3MUozpzV+LdXga3sg8Z8NSPqNROyYHU8a
TSxz4WqquMHmSQWSeYcxP9pCYcFxC3k+xkJP3XrxjMwf2qqtdXcnPKUIzila
4Ra6PX7bESn77ZlITWN5TghFcJQUFk4AaYk0ZhF+/UbMXGAU72uhNXdGWWdM
TUtWfEZTyaaBJb5rsOhu46p5I959DEJY17R1wtFL4iTTdXu3mHb2pXU6dfW9
OJczRROWKQPLz9V9a0yj62oCkdoAtqtCOW0t/1aiQpSp4n/qt74sD74oa6eP
rieY3we6NIxuRhNLxKB/8+eDYnynJQ92HKflEmk0imjC3QPKIPp9fBxL7VJ9
Ebn2JFfi3yA3nnFQwjTfzslgauJW1xBW84HA3QRTdHX148usGKzLvmsvzC7e
ANZ5+sybG8Ddiqd08faXAluOVSRSycm2D6Vmhg5AEfGf8/gWRi8DkBIjQYhY
52XyWTBgp8RoqqXU5+FmYc7JoRudLOWe5ung3h3F3yw0aIZ/Dmy0xLLPv0cM
bPrfZi/8J2wnu5DS7MbkXei8VApvsc9O5nIkMPFeJfis+55Yvlt5ZnRcb6S+
tTig7dKg3/edBVTTC9sRjotp327E2xpWyfuKyi8aZ6/0pfEhsXdAg17LOlBy
HItoCFbZwmdOO1CeKDZMSGdBRhX2v0LoPKvwY+5ZxqEYcMPsd/WhNNfFcTWe
pYYCqlCfj2Ndjx+201wYe/CAqOSSnDJOpw+VNtKHwY2W1eTWcwjN6ueYe0j9
bV5MjbY4wPiAv9QvjpjhtMqk5I5BW7Z/5oVXC0r7MSFgCLEWfeGaWI7AUxbC
HCvhmmPaYZjOmFZZYmzDvvoM2fvD5MQd6+UkxpwGEERBiRufidq45rQU8qkz
BThfC/oEOZIrqMPNCfWPCWosrnkufC8mTPaNG1xJr6AqsOb7FsjbkV/eju0u
pe9mTijlLaXt3pTVMBgK6LOXpX12nxtw8FGiFrbFu24+httoJDvudks6p/7/
g4CyWlry6Eh71a7MT2gtkCe5TZRYIO/Ba945lXQp2xWsxt7aKUmuybI7mxOK
L3ay+t7vDwb/e9hwdK0Kd0ZaisaEiv/u1y7cs4ZYu4eOMEGMj3/SO5DJQt+T
9LWgBrNEKI9C49I4GbmziQnAW2zbGN2ZTV8zZ8w7U7FAyltzgr5t0vBCoCcm
WwWVd9gyxgRsUr4ctFESkmJgJlfPjHmojTgNk739YPZjUE8GtS2l/23HTrn6
kKi4eSLbo1HylCabj/eodDQtqC4P7dwluBHsXqeMIX7UZ2L40sKIFxRP4xLl
lWNuNVe23ZtoszPiv83crH9U3+Nl3ka23l1U0HTybzgZInt5d6C+iKBhGe46
C0UE8hJPufqGHyka3Dkq00S7dBKCKKIl+1WTLwU1JSjaqMLlajx8/Hez2mxV
TBJ4TGBD6vhfFePzsaa8s3LiL+ROnCsF+rnoY7qH3sQdhAbI95qIldfotxhi
FUs1OHr8saPoO3OQMjKjZ1CpKOk6C+1E88IynYVeGxW7M/BAJoZveTCD7kam
W5hODpIb0pGqcORLnrhOqy7KMf9FSwpwpFNKZgDL20Hf7PrI16uXIMHXnCsh
97rPGU1vBh2OZZYGc8hHHhOESYji+dbOgBd0YawEWWQg2Ds5zKygFdOu3Xd2
jKbch/1f2tq4VS6yQ7QpGd5wx8ZRz+nYKKfuv26I7pSG36UHK9j+SL3OPLUf
aF7xELcNHv/KpRt2x6hrPJSZiwGuX09VkGMwLIQkT4VO8+4fho8zVBSOajT3
6qkW+wliNFYBT84KuebHAuZLR3xLlpKcX8PrwryYFO+g/NSxSp7B8/7bBW6V
r5bEeR8n2rKbHDzhgb0uT3DlFmgz8arFtNxFmaclySHyen8Il4w3z078tnlU
9SeBDfycdmjsXEKCw85qKigGixj5vV4avxFEe2QgG4iEnRk1EwnHJKwoqu5k
CAv3YHH3eh99jK/9fFz0gy86yaXejUG50Gy+hNYkpaX1J5zHuOlQPMnP5jpA
huDoBmOsE6IS45ba4w+eIH4HUnPRunVZSPmLt0mkVsqdLEd5SnyPmXVXIpz4
bYQqv+NacMXxfibnsXluw8gSW1oSmR7ybETW6RmKAkXVLFd569xuxBAYdCkm
kGQ5G8IOe3gUmeMmEJJZDPSSuavaIqfBeRSeORKh7z9I4MU74J88vxTbP2oQ
9eu+fCuGR2MzEUXF/+VhHR+WeA3Jpf5x5gGYLilHo2kjX1MEbybVpOOOCXeh
WOsvCrma++QcVRi+BgZdeQNhRWqE+WkzIqG2jCMcIryL2CbU6HFRl9AEzNHP
BPhl7qJslj9IXQWo5O7NqAywTplJhB5jl7XgjgD2qVmD1cv0TPlH5clhVsbZ
z/3dLxobAqFJ+VPJliEifMwl4TqhKr/tC+j13zTsVw+dsdgzYatZDiPa5tjo
VJuRiweiqRfuAzVUONLkYIRk0S6q2HdASW/4x6S73r40UXKhga9OPzk7FgCd
K9d1yev7fhLjpD5UljId99qTR1scy1ASw8V1TDBAbMWbNG4nhvJj6EChczf0
sN4fp+FKpra/tMVG2sdgxXt7I9w8PFCv5f/TWcvrBayWhILGoNgrpdbuVbTl
FQZt5syqJAh+pzWG31w8ISjaJIOmA3xELxigp5tHR8SaQYIJJTvWIGF5Cbem
XhIQdw2Qz+W9KkPXoZMPqMDOfT7vSne/u5hn9nJcbztqM929o7M70P80Ag7/
S8096bYMO5eV9X+OdIjzmHO9n1JuJb5iyAhw25otaYsItZ9pncjQmXrWtOkP
idlZyOCt0Vnwasbnv8WMZvnbU3rikC74+nErAUFEa756/sN7GoI/dnqMq85s
2AuYMDyO7GOTbbPS03hd+uCogna4hBhXXPHt0t2T+a+VUA21Q0/VzjUbg740
JuYxAxlB9wIEoptTfof0iDB56L+erq5AXQhoBesuRSfIM8cKH8ekHVUMMC+h
wL2vVlmD6nzUhXH0B975TapVm6e/SQR5wNRLQ8F0UF0QBdqqsB8NlfzP9lJI
PBvIAEq8g4wOIIhohpCnT1RvcPSXIWltoEbbHYeWQjIBiTb6QeG3z3kseKlb
gUVKksCpkaBlEftImnOMVfdcD/TVKcHYNDqIuG4zzP3MClMsMuOiQoaJyFOc
K7hcZGhG28YzEyhttuXw5a1aKZvtx/5tmwM6ctJbRMhbqQ+t0Jua+jrl5zpj
5yj6eOb4+8KWMDxu++S+ImoyISroPlVbDj5aQh91B/CS4Y2i9l1mJlUINbb4
6uEqZRFlrdURCTCmEGQjuKg0V9HSAdTSir5foOoy843KeCqRTf9kdR69NBr5
tDuGSPjoEjULxIYE2Ohe5FmPo+toUEaTKaYrvOeey+SDUmN78IGm8U8jp16u
5l4gmgbv/s/Ci0W5kMq/NyYpxdlBH0ybL2BqH5JgV7bsb/BZoyrg3gVfmMj3
ZdLzHcBGoTWdeQ7xY5hbM4OkWjegKyUEtyveSekBmVxQR3VnInlwTl3QTAxI
fhToRCgtXxI1vjdE0GNfVLd2S7KOZpdL4btwZnDrqU8ED/WUT2wnSRDOMkKj
q4mitJ+fqTlLlOAPczFoaC3FGBdbyAFsAgsUcUEKTWwAGUzqmV57ORZuzLfF
SUrLvWycQn59PX7rBQRV3nrATga5/3GYuGQsM4BEETT5MJH6W0gMBv1XK9hs
seRDkbwk0O+d6/VmgKD++qURu/1oMoE/gB4ODeRSXpcRFhfOlxSyJg5+Z2s+
zo/3M8ncGkNVFbuU+ndHbGvXqvZiYKkqZshvHTYw/prW3KR304meCFNDs3ac
yFZsGYff0WfDKivLmHGoZYcrutyjpyhDocl4J0PiY1ugfO73AVv0igMTGM6D
/oA2LNEdwOsE1Leebgwv2i4hA4gHnF59ARJOZRzVUi5HJnqhOXiknWca+2ti
cptG7g+p3bURVYt4IGe5kasvRLmn02j6uBSEzZYwrC1W40s9ztUPyGlabHUH
E62fUHqw9+UzXkzriTs3KFxBTJLORT3WqT/gGxOwWhWTL324wAdTdyPDyv9I
QSM5vaFzcSxg018Gbb3KWBZNjSAKqfohiopVxRRQOm9vH76rc2Qtsl1tlOZS
inTelRa/70FpvARqOMjbKUd4ntyCoRqX9YJTPW/Jhtbz2/5cxzBNX6i1H0k7
JxMJKyF9WFYX906gS34I0/GRiwWi7Emxg3JBc9JlDyCjVErrRug/eYWu7Mgq
qazCyHUQl59Z7kT6eFXCSqY/Mx1qmtzJvF9KznFV0yt+vuOR6Ngd1Pv/Hntj
yiJC0twvebDXFZye2Q6zHmE3LYUUnokpxhwvGiHteqd/1pDLl+VFseQQkNiz
50LefceQRcyWRqXmkMZPVnL13YXEejt8nm3qbt5sCjO3jcfbp+V+sQz4YbcQ
pY46gQMeFYQLYgqBdr9tEWZL4Bx+a4GweMF2R/CsPsBz0TzsH8B/m/4d1XF+
jPzYoqr1ZHEoG9ldSY++qyXGReDfnFpNoPAwKsLbfe5Z8b0shPN5VIzZAsee
Z1FfsAyT/WaU10vrwwygK3U2fwEcuzk1nR6ivj6nBVl+9pzii6A/tKS9+1R/
iZjY7MmgbN4/sc/osSQLBP2ThDgoiE5UHgIDcdUMjBGfA2rXR5aEpOSIm0/x
qG2aVxpEtA6BpGN3CHt0lCeW/oDUisDvI8CTo9PFuKc4uk88ngyDBP0rJrFu
vUf8SETEo8osbbzThWm72msc9RlydZrzAZRRqSnB9MivJO4Esq6rKniGVotV
j+jSBfIA1+iXjmY6wySrmj6jdOvUN1ggyFNz4WRU/Cuk10r9pU4KstDWnTm1
SdxB9mZa1TTpj8kUZhKsY5wbNFHXrmxq/aRQjScc0OIJtWXPlBMjyekCdEYE
kKaxih692IH9xNd17xF8uHpM3f1M9b1yYmuCLZkaB+shSqWShDRjs/ttOH98
/3x1bzoKfsndMn4HNGmEA26mwGqn/1MIrwFXN38Fy6PguizLUguftgd0HUPk
pc6bAc1i56ZCsXFq9PG+Lrutwyu7h10aHQKGmNawesCnk21AXEyaB9dQA2Cx
mLxfNFTRbHsa7EQWYf7EecwrSv5by9tWaLYYnVbUi5/KOuEToktN/FJLY2Bq
NH0eXw0ZfdHOPbiht+f3NjkXeP7Mgd2Qo1naKOSquGJ82M0KqUJK5hkVZ+zT
m9vjQcmJvgZi9bfiGp20ozCpE9T3fA4q/yMLE/vM0Zp/okTKtcHsrAh32mVc
IlDmG7BvN1vfHBQRUaXwpMm5ZcainZbz6eYc97motIZhau67yQL/T4wqIX05
9Rxv3xGm7OxRwoOhS10F+w0YornWfYQWHFxhNM0h3DQ05oEWFYYgcvTDve0v
MRWv5Ph9tY8uQt8gGSOQPWI7qrjRDQfoVTRaxlwCyf4t3G86wufXk+q/EDix
7060pa/Fug/xmnvoNq5y2/4pEa59hOIy/w1Zd4f3n0bTxyRet+I30lv7lej7
gT1WGIELVkpIGdgT5mrqiBBYf+AgltkyF/jVUPngjqjRMuBPC0Bn7I1or9sl
L5b+cKpcWtLlXr7Sb/S1lzaHm9DyWUoBTXsTX082HQcRx1MgG0SbhsB18kV3
L2wilFfI+iA6Z1c5Bh9KK9k+91pfsef1/5h4rktVvqpKqpIIm5K2hXovEthU
ZK0B6/ob9C5RtbLaNjj7dSfeuMJmIFVZv70jphW3gZ/BiYeupFnVvi6UVlap
QGPY1kHMKIMqlz5yBWOkLWcgRpWVhPLo75+75ossigYNE0qjq1ksLPi07meW
rNKxTim4JWlbUlXrVa3t8W9kFeMqNTKdjR3wiaOCa9e33Aj5QeF6OvovoPoR
NJNhzrsSoh/estYu2qjUyp1IHauZk8RsokKtHW8Z9J8xGnx9+SXBV5vZdyUV
oQBedUpt/Bw+52cGqGqe8YXrdqs2TE9KfXcYmXQirsXseH9RySEYodU9eD9T
RumzeW4irBRUPkCaVgSEYnkR7o/ac6R/d2NQg1kUqnrA4Ngnf9R+tNqZ4k4Q
+u8RZMOA5vzJWCdwWWjzz+W2fVAmCSIUvWnnozvxh6deH4DAbRyP4HWMmuzE
fyTlyg3p1+075GAtP7wN9WwtB2tjkljmKfTHrkPiAr51uQTvBV5ytRkc0tyw
WLcRC4BymfZLVC8S/fHSka7k+pSUx/xbxhMvajRUiZfQ9RzaX5FWgnEgYped
bSSnUfqHHQNqfkJWGh4lHrZ6mMiIndWwbXfroCY4XSg1opaIX+K1PMcsVtZi
F1cHd8+O5gJk7lv6JTlVjXy+mdjk8Wlg4SQQDzvUsQrTirQO0fjEjODagCNL
uC6ObCTT4xePpSEd04MiaMBjpdSOks9zPzRuz1UzfxVr4hfcMD/WB8WW5PPz
ZvB+pQOoFazef7DFkK9Qt+viTDxiRSb2ZoL4hAENn9OZmr4zhNk/AY7zj3x6
+qtBdhj4eaZUdNpmyPO8BPA22OJrkbCsErb9vI4MLdis+YTFa6LsSLUVOM3M
jDlgPQ1/fBEvYB9go4NcX0xCtfgIDl3fdNn4sTuQU7+1sXLNz9PPA0KyboYN
Y7YLO+XBBjpGoUdavw6Tf/mNNPKBO9NsVTiOUjNoawmMvkER62ApI7OwD+Po
86/VtzHmIuIUyZzK0PtY7U7Q9PL0Vu+or4Yvw46VskfLKthLjF73I9pz+JQb
IeEBEzjp3y9QQfYk+U0epiOIo3cVT+dRpBf4XnpzyzFumXkhg19XLKAFHoH7
ey3q7K8XTV57KBydPlCOaWihZqujO3jC7RiZaxmRaT92LNbOLc7x7+W56T+E
cM5zrRAp1sMglWKSTDDa70xSUI3Nhcmr+3/y7Y4yxdS7z0uHuH7JKkdwvzac
thWczLq3jYsPja7dNA6SYcdSn3IHx2Uwq/ZZLwTWO1oczrHRjiRnzj5cVUAj
zQtTJN9WmnyYct/+/ZP7N7OS77BIep7HhNvrJXrbbNIdMxkbftVuG9hwPGN6
17pr+P+zPfEv4c8lPcIvvcZc8G3d6PB5j++y3QWIQ99NOT7f+IZVOdzkONje
q90t6AsxPSehQuvYJJXCmiWlofMv1gn2+ot8APFsm5k1zCaggCC+xuJtM0ye
hSk/srWtiIMpFzWpnty98mu+yhAEJt4nK4ye5vbPp71P0LvNeinzOToTmRll
KQflgS7RAjvKLdA8pECFoMKk3HHpmnEY+VcBTbYzIGMWfvbEuE6phzaH0QW+
pM1MZZQBD4Vv/YRM6f9R+GP6soSN7oA2PAV6I0l7uP42PGE/0qI71981N9nT
jDOj0RT3f+ZDUZGSBTM8BCEzDUqleNNHS16gd5QBudscWPrq6KnZfIKN0BmQ
j22KsOop60tcwJ/wrWSmWmZEPhzcBiAQMdFs/+/EpuQ5D1J44ZqvdCtwbfGp
r4830a5CSR6bQD1g18XXQQsZ1ECkP40REUYijXBOHH1knTJnfyg92RX2Y3Ov
o2MaKc8rWMGQOrC/34PWyN35YTu0re5D5N8CkvogetBCwQPjUuMDtXNlqDgT
H5PTj/9Uxo+URikMVlgcXMJzw+hHONFNA8/vZQkBQ5rcF5q7GnIfIQS5v84S
fRBlVdq5kvO3zoACFghIYUdA3c5S+iW+qzUSTabC2H21ze4gwo739Trz1V0i
zDSvnFvhri2naDvHEXGIEjZtHRKDLB+oD4gucXpBRphJeRHpmqjvUTKcbSx7
+k4kyqTkpchQP8gwvXWq4kU3gpGhrJWjDEoU0pmwOxPicEF+z9ZXVlF2leED
kGZzTwwPft6KId5WQzDUu6BB18TeIB2P8qISR3oWTzey4VN9KoIgZtJ7yvuf
+QzTQ4veqTDD0C2jJSEGop720lQu6CJ1K8nmty5HAbaPQFL/wDUmbgHMjbZ4
hI3Y0D5Y/mez74sSxhW88nor83YFssRf594tV6iB5G0OeYjDuZl0AgOfNRuA
Wc6tKm+W0cNnXdu2BrSwHqESYBauLEmzvuWqnoNDZLQeprWfBIXNJEuufC+6
YLyVBZybfVzIMh1GNLgTwGtreSoZ3HSvC+XksnxuIyYFOMnMKhk5iu2nCMvT
vKNtuHbygYz9sR5VABnqCiqgbkTkA3qAKsnz3U6YpSJXREXjisUxM6fMxFAW
D/0yhjWD98/KERvPVm7j7dlmq4pPSr5f9DV6iSB4UPTjw9AefUm3qcetLrMB
B6ZsvkVTXIcsa/E8SoMfnPhRCHL7pR/fH2ha1BL+sUGrKimey8MC1P5QYqhY
dWuy4J45bpx837BBly9fI0FYphurpAes+48jbvLoGH/Xgp6RLwwL9XSwSu4O
UqGOsY1fC3r5MSK2+THOkDP7cbqgY3huj0hYtbHrReRQoootubK0pRREUeNw
YBotg/kUjWfOnN+0WxkzOXE7smR4jTbICcNCB/lotdX0M5rPkmHza5bTUVY1
M8rScMTTN6u06/XPEDpG6HFD10DalTCZNnp30UZjxsvlFpz9BpBhRox+jLuO
UIR4xv1/vmTZR4a/fVgkWZ5fsy5t5YUf/WGyRPicE1xuRRn42+ovaRWqj8IW
lCWX0xjzJPL3hsMRmb+DCSFjv/e1MzJ1J7X6zQSp5RR5JV3pAd5azUtW5u5F
42uwAK7A8N+WJzvFdNpJiu9O3zBkwBWz5qepQej31Z57dXOUOoPYlkkK7Us4
SvJxLOJnTs0ZPaFJNKrz2UUgfgXGouxMmbbZbDJBZkXBKj4VEndyevr1VUE9
+tfuHMGod8o/5TFVmirDNEon1w/dSs8hphY8aeU+xPPGoWq6FZyKhv4N9/xF
/+poTvCduc3RFAGHg4iSHeuCAPLnFbNb2Yq7oqn0qzPvPrcWDkXLhYPVTOvf
GVPQNqNLEoWFRJJcJxceHDvX3MeghNTLkcBvFOlZ6ExpNOI8tZJGfZ++VDC1
mxmzHPpJKYGyVDtXIMtQQ9IPxcrpgCygso12rQTI2EUvr7IJWw39e0u487c1
yt4w+tRJ68bXEBtGx0MlH+NbuacujeSojYIUdvBZGf5QZMyLiitwxARh90E/
V/3g789EdL2UU6wEPpsRnKO85tM6c85QJ9KH7DlfOf/71aVoOAoTjoSro86T
XhgR6+KdGeNFxKnX1RV6PgJjv34mHJEsWLsd1ozwfrcGyejf7XbdbJECRYV3
mHyXYPbS/Yu4Dc+JzY8u0dGxxzlBp9Vxb2fofpVR98CFPMhr4wqzeIu21hkO
SVZp9iRt3q/u+Nt3PEDzS0H2Gva/VYb5ko6CfFNhfiWJC/iI/cmLLeMDsfaI
WM60N2QUeyRWdWwcipEI8D69ksW/bA2YJQZbJ4r6ww5FDrW5nRVJS5KzK9bD
z7FFyaMdipi4AD09EQbKN6KLtTJCA7mvXEmbg6qBODkj2MnS2F0i3Pus9/ao
KttWyqYqVmZreAXhGuLm36crMCtjRIxCt0Dn+PbyE4x29Lrzm0zV8dNzj/RN
aOgdgj7K0zlaePxTkgYE4/IKxydTI5Sqzf9yfPnakWZvpmeGnbyby/tbnff4
ixnif7MyujUrnq9sQ4n1EJLFpD4II5yPn0Pg2RnxjpceNtgTFMiq+93GYHDt
MmQlmOWGvxi4msEzuAFC4SYqgbchqajdKenpkcS0PROLy7fIzsm+hZ8s4eQt
KTsP8UQ5Qfl9/zUbSzF77K+6Odf1/14SEBo6gnmuaI0Z4xVcGbsKu17UbiOa
tuzJ4cZLAUnAHI50geSjnOJvSqO25mpYfz5h5f/s5+bdpaI99VRenzz40vkj
XKThba+GscGX+BFQQxAdBsvf0XXa4AKl1CHVfBfneliTdX2i6cQa3Rdzo+hf
pPYp9H4ixfpO7mGYXaJH1+tYgJbgvxNvSZBOzn501IzMlyuRJ/ApUFMzjBRZ
L6Lbca5vbf5BunT53UtWL966r7cQp8QXaImgivrqBHvYy0Q2ycG1re92xVvg
jkNNTPGIbFt+4cGK2JlEiNuqdv0KsRTzfRNnSLsKrMdBwC75OMn60A9vbUMQ
UqFQbSUcIuWDbkiOsE1PZMPD4ORjiZ7r+QIe41x1BOOZ7ZIbrt6U5ZpwZDzk
WtR/YmyEVOsbsewtYHtq5aPz092mI9p9KEtxfrZeva25ha4qqRRFhjKbLbpQ
S1lWv/WYhBP8WzzxTl2xh9nuRhMaRAWn1Q0WmZOQtTs6LQN3/htdWpM5J3kK
rxCcGTmVXW9T7myiW/2NSKBbHdlatgPrm436PTSWMezs55WOKG7e5jn4mOUe
3j4K0FcCP7IoWEcJhKGMz98T8n2UMWl/+CkNjjOOtldx1C8rGGoir/23op4V
8a/A3+w0Ds3KRdFm/7CnDGIN0ixosfSmPTu2xIyYXm3h7IZeIRjV2vw6BxwZ
wofLZj4zDnunYFKrKHfc92MVPzpamkRDhbdA4Vy0NuGD8WrpUt8s6K/igHi5
5RJibS7WDCFXFZ2HNt6md79MaDo8VpqJIeO3/rQc4h7A1sumLxWOY8YzzOqx
13nj5S++c6TRkPqTmofGfzB0Y3U62PQI0kMOh3S3eHpBvg58a+YuAygPT3I9
bapWAKz80jSE6f8AHPnR2+uM7Epz0neflJrHwJhVWy79QwlvzppDrQ8hTlBK
K7n4xl+VL8jh/6F8kozkeiTJpTLzfAYIP+QzFMOLfM0QZag4OpqIzTbX+WfN
kAynwm9RbrN8yowyse/C8czSjd7jAATtAs6dOTUGRF7enGuMnKYHwJXGpBG0
zms/Sbg/noj8tqH9CDioeWVr2b0FuETsKMQgPma2khVAbnjygmpHlsckgoOW
gm7DyOaAiozhE6vOT80BHRpRgqUgBR45uv+y5cWSLF6FSRudJc8tdbOB3Obt
S2Y1+IdAmm9P7flHnK/mZRGSeN1ieTqp29qTzgJjyn7tekuNCJupunsWp3j1
5fl+zAgpkW8rNdz0v/e5/xXWezbpn01jqKlWC2gxGHxUceDnf+sFjna4GHI7
njmRqqrFAhG9UF67j96XyP7mvL5m0uKMDskXShQ6fbTuOKhLivQ2OD4EQ7fx
S+jRD7M4Rc2GnV5ldJOJFlx4dEtBEZtCC4tT1gU67Hbp2B74zl+CfbX2O5zM
TStMdNPARPbNygvaeUz73LO4C1min66e9sI6t16jxYF/z6V1RN9WC/qrMa4n
6GNj1sIMz3lQ6fKOpHzZmEQltnWrPimfha9LYoSICbV1IbqTHiPeOJZGLP6T
lSMRY0AwbyCFuAa6fuxolUXGQUhGQ1cURAPjHo/c8lQWnMxzm/SBCOJS52ZK
qNHXspLfeC2OW/XhO1mgsueHkailtn1L506+7zyJ8vFIZYxfM8xei78yk/o9
cL/mQ/QBorSk3pdopswnSwW9QkDH9juK00i7+u/dAJY1slHkDcUo3ODQfdfe
ok5UO6U0O0kovME8hH12X4D0n9cdQuLDZvKq3xLEe98FqGD0DumdfWZNutl9
1t5B1+Ty68Pn7kfTrko95QUPOJEkwEvllS+f9Te+7lPY47FnPLzS+gj43dVt
k76B+w9kJGucMffhNT5fwvd9wIazcjC00VGfQUK9C3Z8fD1KrumpHefCSRXM
lK/j0/2EkVsxkReWVE3P1MpYptD8F1wGYj9FX0TbYBBio+rBZZLhRR8wyHR8
vND5TSUKMvw2HaQfEt4K5RPfO0KjuZpw2aU1u/dVsNLYkVgFCuCGZArynZ7y
evOk52qJGzUZ4DdSml4Gf2b8CXNZf1FVjMgc8Ee/jbu0sRCuGOs2EDnrZJAL
nbl/EZllncIPIqKVkw03eEruZzhiul+EUlAZ5muCcRSPBntLIlkHFg1brle2
KQRmo4R/hupYq3JRebAheYPh3tqZkiLEUs5qQb1otutFVjTA3H+THE8UNuTG
BnL9ujITX/BA+3mQdc4CxLnN47IUu/PeRehjjFe5UkOLROZ254N10CD0y7Bn
KxNtYR+iwrCWprM8pNd/UjMSaRMNnE5BqsJY56Bd+eHOlVOF8wTfSHBarRvf
HLomjeVGjoWWw3l0WAzFj87jU1V28e2KHmUZ17KrA05LGOweko4IK1ETTnEs
E1PhFkSHiS73+nWT66Q5lGDtMhowo9hD19823INA3L1rUuvSEoWWlwXU91md
oAEIyku0s2sL187O0WLudCkBE3JgHs/yO1MOZ49oLi6fcF3JnYZUVJJ9Bkb2
IoqFtk6BO3tUUps6nR5LqFFxZraRb5HiAhzypk3PSipy8q1NDtMKQw2Vgdre
TcRsKh92f7ue8go7UG9mPAdJbDwtkPvVsAFFTbnlhfOV5XjxpSgbez4uDNMj
PympoqpB+AUzhVB85yQHJGz+eVL1ZbZX4a6yMskeHk3zN8VWBADmJW0tY5Zx
b0gg6X89wgDT68dit+KxELo4P3G+3+SD2p2vuJ7/gE0sgY65vmPajW9y7nsi
oO9X4gOq9xNHL9ifRJ74yfiIB8bB44x/Ymi0mdJ4gD9iOe4SVryKSzg1fcGH
qVqlvQmZ+fMWmwwr5SXCy3cqGeAq+yD+F8uzbdUj4xkcvRGxkGavnLZj+5vE
vpnVN2xlsO9qdz4tlJ8J+BDVcGIcCbT0F16Pmrzupz5LA8QOiryvZxB8s7ZT
b4DFgPpI71V29GWXN0Owic164ymRk6UghiJ1QpwENVX0anI2qq7GD6HDw462
ExCGMycIEqKSVvYFv9BrZKJ6M4YMfxtrnn09kPesW21g5Ny6MYdkKvJff3hm
iID2VIvV/hYM9szCuNUP7K3gS3PsQU+Dl7BZF7xACosrCC9qjDcd2IXCWzj9
JgHRsbVNs5Cee7M+cP8QG+Xco2JA82N+hvILV54gSTpN1IHVkt0E31Yd+wCQ
BvtkjYUzVd8/62wTwP7ZSfaHiXTr50fMB8hjvXF93HdN+6BnhurAFjgoUfla
2w8AOAZMbSrPjeWHgmnQS2eDou41OZNLcRLVQSO87EYVz/Z/ex1z25kM5tNh
PhyC10VBxXK8Ht9NnT8LhoRJexKeDGx6HvWdov0dgMXJf4rPqolp8qrNtkyh
zotELjOan2J5r0/9IyMeFYfnS1U3XyGOu3WoHlG9SExR9sXmxpBbLw9c5Bhq
9NOV7hKVsgnfYvjN8MgJz7eM0Sw0R8kK9YqZdaYEX8z01Hnnz4WOyC3vJZwA
pWt76kenduP9aJrg0QUC2ytoJC1ANXj8LFIJoQDYYYhPPymf3jI/NF/cLtY8
uwB4+/m/DNKPkzYISC0+i9DmEvpe0IOMGM3XJjt7PT1JkkjN8Fgf2CePM5iB
a2Axn2Ohtuf0Vn2t5KzoHhSJsrVeZP3A+UUKp+MCXieu473NVbbsUfEwhTsV
jzAFgbjLD5zwkIyu/1NooN6XqwsJCpoAq3jSV1ZTMWVX4FAsoomM+9NL3wo8
tlMRBDQuteT0E2OlFxcQcUcEw+aQpxj6B3RjzjytfrFQkBX5jMWhg3LpCTyR
cEOWRDoOJ3Fnwm5Ho6ru2Zx97RdW1lrurdwi42MONU2Aemdy6fog3N0EA8Kd
utzUSRsOfS+kQgJj728w90S9yfupQa4gnxj6LOz9lL8V4mHgiY8KqNpblIhk
UlRmFm1xiXzTHtlkcGHnHaIz2czpNXx4awSUZ9XeSxRBvXiFjWastb39LiM5
brOmcqaW4CvrfpEHWYX8LO7d070DiZH4emMVwgKpP2nrr4eRC6bv6jCcXheB
Jf7vl0WNUQUd1Gw/d1GQdBnK7olcouO1Jd89DvuHUs1doxWB5lUMvqth1fcD
Oy0HbJz3lHFlIr2y+kYuuoLVbsHXK2Y62bY4/ZULLe6w62bpObDJMdBhltj9
iI+G1ASfIrGSQahclZcuDZ01WHcSwSD577mtQiRkMryXhD8LyNx0dzvqF5Ws
JhMN+vjtLQugfxvKcMGsL+hHeiI3mTAOfMj1YPSgb2cfR+Op/YCilie8p6jX
Hymrq8tkOEl5VO1oFeRJ0g/a85oMwcn++e15iaYBndvTiXayn7kHG98QC1+u
A1ql8DXZKXbCDvewcDDd3VqX7Fe8M44zuCym/RuqsBIeQ4eA3FPr1awbDJ6g
K+BIc7UwLx0POodGPwT0N9MO5ER38ufjOfamFTS5iVVoeIcyBbWR0gl7/Yi9
w6tM8Au6IcI9AdVyQQxDNrRwQ1gbe05k/PRtOConh7vmBFYeGi95vkBYTqjV
7fRYMInivtesEXTfbMUEL57JBYinL1xRmNWu/9JNjlwyysiuXh6en63qmMpg
TVFWEP4Qyx4IywlxAO+Glmr/MueS9qFfGyK5dIOKXI0ZLGYVbOrd852sizCQ
dcWRxESR7A9Ba4/+tmWpYcX78+3aeSPQrT+cMRS2z2+vmJUF8UHSQqDUXyrJ
yQ5tF0HRc2i0rAdRGx1FCuFbebdQLlCml+kqFynX0sr79AjSVgNe7cLwQZ+h
C7QsvNgFDmag3RXkRhGbnCVccQTa5EaLcL8cJ+h+8GJ+rYGC5V3ZKjfGRijV
+3K76QQPUpFU68Wrs2Ypr60pY2EwPCMC7i71xPr8RzbR5OMD8zb7RgEXMkGz
TIxWaEBRFxpD1DkKSR1N6n3CnuOWVa56mb/bsRjKelGoh4oAG/jU5HRDia00
ObkVIcNCWQwSUSzjoevAQzSEOl3WCcAlrBCnfDoxg5HY4twORL9zOXZs3W1n
XfYz9rBe7sdr5tJdx8wN9qLS7m/PlVcE82y8ju6JFalMW5JA0g56WgdXt02u
onTyHKCkAWyA3AM28Zmv1XfCkViTYy8a2ZM64QUb3P7p5giGVaPEzd/wv6a8
76rdiDDoPPcP6o2v2L3Rt4xXlPwkKemMb+LbKBafVLS9mqeS7r4eRg/sKL2w
zw96hoiTtKya0KPb6LGYJfDqbDrjgOPcR3fC/FH4S3zSZ0QmMzeQcfYm2r4w
EfdtOdEzgU20XTYxK42E7lsHALlw7VTGgdoO3280BSKvI/tGws7hQ9P3khEH
wRw0TFxiSIb1Ntf9wX680YKHpe27xrIuRopy+53uoC4Sf1JJ4r4ACJA/XPcf
e9dRcKJxBOl1f38Ob6ku4eaAuX3gnWl+qZl2jYJ8PAmARyIzTIgtaagm9M0Z
paNAkIJW29zr0YCFnaIB5c09ulwrbmHSUxr5o/GDJReG3170oMa1RGhUApAh
vTpQdWfDg/sJph/DBZPItOuxZ/CsKQZoEK++EgQbgTIygMLauaD2TiiAD8oG
6kd6a/4r6AR0dWA/xuMMLcAN6EKX5H9hsvLMDcJLCRb2wqjIgF6p618CgYE0
z0vsMvvLV61J/AlAf9FggE7yAqt3/X8Dp/UnN60n1qJLMIij145C7qoguTz6
0SaDrnsZoLCFp6VU8Fp7alOyEziVBcr9DviTergMY3uHpkU3vVqXWTtfnrE0
yyIgGtYVVB/NFsKwkNEAcFk+tAelJ6KBFSsisU+8t4myd+beF03nyYlpAm5l
qrypqxRm395cB8/uoqcUUU3lgrlYXS2SMVPQ14cLY6O31+PjymbK+/OLlsc9
CdVQvHiLWMCUdSc+TJEBq8DhNugeOxUKKhCEh9H2S1fGvQgwMLy/F/d4xQfr
IAXtEZfUL2RqrvISMSfRcUMkAh/ian5ilL8ObrRRePxItshEUh2MWSzHgnOB
CpZrivIV/lirzh6OHNVUuyinEDmMwQDBTh1v/iZeODkmZZqdmKyiRmpg1UOS
B1Jv5u5BG/Z0HIimVDQNFE6/a8tDadfkRDUXn16SX8hVEy4YsgWEXTsw+Zjz
jYCsldbFo2J8JIoj1ggKCm1L3d2TXaT4i07gA2qmozxPia10MqkC0ZwZiabT
rCMj/g1H8RbDeX9s0Esg2MxLlkAH3wF7H+JeL18mCGRV+g+ANoHMpGmP2a0u
njB3xTSHyFlZFGqeTo0nKdLcW8BdMO9+kSVVk+IimVrfnLjE9S/CXa597G2p
REo0WrqlJAFVQitnCm85t+OjYue0mWfng7S9aXXB7DNyXXiMUesUzH3eaOXP
4lRNCGCLfwI5wZFyLKWlPOf8NRlpDk8uAEVEABmIt1OjRUmz5ffKL/IvXoJO
jjigaapBoGtsVYUnEaWflpba059MWqb/D+M4LjxY/+NrMoHASvfELR1sK4Ma
yA69zPYTqMXcI4PLmngJhChNzZO/U51vB50ImU/l/t7LPxJzoHnsVXs6zAxx
DP3n9uUs65NgTbRqNu4+VY0jIFolqqeXANdbXAh3uMm0bNOxk3BeUKZxWLvL
fN1ITks5nUNGbz62kQF4PDD04hBlhSfZiK2RfrxWBn+vIw0NaowpOhXb8B0O
lD6DrPXc+D/e1F1A5dFpUqzWx/fkpGTtAl/tAAgKrrukf8xatJZI8ySBilMT
MYiXpsyYnfr7mBGPUgILXCVZ5nSvgdsJti6yp4sEOiWV+7w/kaxScd/vTgrm
NDpEQcCnc0+td2qsj444O5GbJJWtehEHtx/wbV6BBVk/Ch34kdrPGiAbpKyp
QHZQnnnRB29WtEBITjQDjHYjClXkwZBsreC2F2CQ3vZBW3HFcP+BRt8hQIYb
vqwin+xtVTVSpRH5cDIxbEHSehRs36cGbThTi7Uy/Irb1JZLYbmOKqev8+Y0
R4HRDt/IORVnO/l77FLu3skuk8DkraTMpRFZgWGEtyWKa1RYDiRnSRdTqXUi
Y20cBRjTx40hdNLQJkdvKWGlsLLE9LaFHxSJY8Kl5CbZzKL4oKXL1k7RFXOC
WvFK0J4Rnr8RkfdHUyx1Q2oOs35qhzhPd+R0epK474FTnIyajlwZT7pRuNta
PchfmkFcEzvB8kwfQI12YOC1FmFwxTPrzIAR/DJSOU4n2qOOTK+CZS/CfnsM
11paESotZa9+HVoF6kLIKh3kNiBYCkCJqbz698JJwQlgBwLbNhXvqSsg8WEb
EallFZoQDD3tqJd/1Itf/9UA0fFTYeEI+wbW+jvKt0EkxmoruJsVMRbX4eI3
RX/QV3AcUkPV7BkkxX0RksXRD2gQd5ExOSfLy2x4Me39Emepz0697lqigO98
9aXwr56IM1QDWbWODBQjzAZ9nE767bBO7siQKGbwwOzJnylI9iJaLcMoigEp
OlX1wRipf+35bDtxsOWGxicLh25NxJgY6iiQXOZm0ktHF5EmADpqFZLfLXGI
ijF7ZIOAt1awye0O3ScOvh4ItJn/uGqJUjC1uojrHocNHv+R0mIOI2qT07ye
c2+Q/ykLkIGUu7fSxBB9tp3TFi9myMQKC0+An8ANdRM6yYrbaPFxqPNxV0RG
vvm3zY9HYLHoifM2PhCNjmQRB0BO/n4Oc7JJrGsvE/56Q95hvFbkbZDuSVNe
a+OoRhhDedwa1jBHUUBA9uvv2+b/XSbOlpHI/YXOaFROYUnBBzDKs+hIUK0n
zHJV8prgIhZkGk3GMK1REvFr8xdijjuoTWd2e9Q7OA7U0DSGbbAJdVaHcl8l
bsEGG1IgBDq/EvUOcVpZcs+jOm+sL8hMC2o4fYGrPkDc0o9klQCAz+2UYCkn
5NWQqdVK+hKg/i0tImjNQ8jIgwtH7LzAkauTML2XHeYGorAQU8naV0dva8oo
0ptbT/N2xq/52eJL56cRT8ib2ahRJy0MjkvmE72MOwO+dor12PNMrY/vwJ3B
V6aimoswIftLU7u7P4elewghlBSazvsWpc1Jq8OgCFqytD0EwMtBfvJEkSQp
+yIic4wPpZ6+SjgvJNwLX3rUlI5jiRTfhN8++L+6qH07qBb9mQayHwdMlOnS
wgfwiKKO74TqXpS+M1tGNDO6THfwGaiFsxvtt+KZZkUSd2m55QG571At4m1v
+RfyuzNMSfdQQFSiqb71vaUvWlD/zGL6G6thzF5x5rHklCPRuDDfZpiDS/k/
IznheKNdxJvQlJmQmTHoL5BvwXH1/pel0Jn6OEyJU8V2Ymes4FhF8YnyARgw
nLgVvloBl0IeFT7X0ZDgvuU58ORcRJALU7eGBDa0SJ+IOJqf+USx0ekTBY6+
J2vnxVr/pjOARKIqVqjIv4HMH78f9KnQsHmreOXIn6kD9uZsflwbQyoqVGlF
d31er4Hojv2IRW+Ycz3Ywsi0rtJ618ioLfSL58LdvRj/hzi5mQKwGSryQDYb
N+mBzQtcUSy+vdJnK9xORbKveE5W60Xbd3NlFm6kkyu1b4A8+WYaLrTLu86a
BdkHZF7AogHgSv2A478udbIuCPxD3ZgtbD3KrKm0b+byQHv2MVlrdooCQNLf
NWIJh2I8U2hf68bWdUSa7ole4caWFAm98ihOEAoOxk9NyohguJPz8kWWmCDY
ix7qIzIShyfL9Cz6SRxtMbYorRR58hoSs6H9cyyNKe8GJ/HI7+/6rhWLLtcV
axguQxesJx9XsEk8gNCzspIJtVzOvG0CW/VNFjaHDwxJqBNfO531w06kQ254
ItQsdgI5t6PshpCb5BrH9qreo5jBXVf4fogJ/GHVb6mjHLDjfpTwzhJ1AcjQ
uW7Kg8qMt5CvpkkHgEfOFEx/hwE0/+hkCBL5pKM1dxcvwf9YFXqPoDqGMVrS
csT79MOjH1XWSpxuGirYAruKSdFiRUXp33jHF+h9yKjm8wDfXo/R6Fr7f56o
LoC8CfsMgJTZHzhKQaQvDBGrCE8eOcZ+TvERGnWE5VZv525v6Ni//iK4zUSk
pDIekvhfPK8W13utUbLkbNz++SAPvi5oMF/I+4YI+bXRnG6YsX7wXqW2XoLI
vPfxsiMOHoXc377vCi2gm6LeF6COa5gmCrBENzClqFWhnpdj0uDiJJnSIKSa
ejnfvcJ7BWz7doY330IIwuWlKLLX9bgQj1ifuj+ijiUIo12RkoLjyH9eRjoy
zVdTK1yWufXnctpbqfDKisbk3hNMoHy6IO1QEJf1oLYT34gvpV/y9LiWe4fG
bn+cgBlZftd4D0GVaivQ9PrO2grnTGHNxQXAukEWNwbkTSYFZ40fwn0jM7We
K6gySlDpMskmZkN3BIKE9vnbi1PYfKjMteIoIcyqqR/ZHkZHD7jlvnnocGD/
bSa40riEXQbUdsHjn8RFI5wy9oAPxlLCAFvOUaPswCoWSPyIFMZG8LwTo6ln
zW3c6jMrjqiAOcrkBzJ2vcZ9vIdRpObFNJO+vTiUnCbibadQda9DYrJXioB9
why1w9iKV7sOIoHPWUtzAoxeioXMHFYrVxvG3UKu/iL5Rd29iWiwluA5GQVG
ujDvLBqFDcpowQwav4VZ2aQnFzwZyqGsRjJIBwjifMGX6NDSevZtVUU6+GER
zMe3Lx9GwsIVQOQZnLjZQRI/5HijxJ0Jr5BIBOrGxOc/uy5+IaXR6OWqsxdB
+zgu6QM/laQdg+126FljkL9Tv1lyf7PjuSCqQzw4siphvWAQCEKJcBjPhcKr
NlCinX0MGvbhRCiqG9pWjZbwzlRIHLC/BiEAj1tF/r55Z1y4pTq1CNpge9BR
RV5cns1Wa8QA/Op0YHIEFI+Qp5nOsQVM5K1eDfF167Zyic4kk26fsCJTux8n
704qEp6Tf3rCatZUpaXmx0dwu/uzj8SxKV0ZArT7wJXOAB/5AWipw2ZduQOj
++FLIiBJ/7zZNFv+KLcy+ZExRt9Lpk2suG8My5ilyb3H/xvyQRiIw2LlWPyK
qik3xR2P8BRVDgP0XV11uIjphY4F2M4YWkwtseLVJkvIEWMXqmHqDjtnGISU
lRQm1fLYvs7gu8cgLtt7kFjGaHoI+oihRRBesO51gcns04raYMAsPQ6jM/kl
iwKCSwWZNuNwVh1e09pV2+fXv5mqZSVSuRPpgcJ9oFVRhKfqlct/I8FTG9HV
e5ZoRJG2gth+Q+6dcjXV1yo0vGF8wrrU3a9PzLlMsCbcVlyNZryZEbVTTL0R
1pJF8I54vsqsayp9LdU3MNr3TOkXIGBxaunc7A2IrgbbOtD78EOogY7lj31M
NNQNMlhMK0cYMIlQc2LMSYGjbfZrHoUZ8VtgkHf6TeHbP4SpN9J27dX3PGoi
a+k8K+HPQiYv77wnU5KCv+jzoEfEVy2ElTW2CbAlwF0FjvFsYnUYhV+44sJE
OSSJrY0pF2M5GiwPhKsG8vXPKOSSiafSYs3FhbS+c3XrfAp+wkD96D70e7JK
1X9Z74bCblkzbJINjveoGRQGwNwut12S4Up6UrN3DQIxn8MdxB4qY7tYde4c
MTsV3jBB/s9dNTgjMFeFb9yE5g9ucZlO90JB/SbgNEmWGjFE3aI/pcIGE3Gk
PvjJho1rBluqBox4RbBc+SVlGUsk4Us2mBxdW4LFpkf5TheUFUoO55374ODO
WDaed8uM6H0lYX3TWxf1DJElS1J9AhRxauKvgRfGWcMBpA0zp98w8234+vwG
askW7w+kD+shwz44Xg09eskRM+NgrnSnPJRAG3PBx0r6XWiPFpkTxaIABpud
iOO8Oxd+gCXYpToRqkB9c3CHgaFVKLfqnyhc+8+2EqbzVOtIDLSoDYV/NbFN
0cwTZQRbCpyNavrb2b/npuWxWejNPIyt54eEcExE4mWRBSEEd0bR5DaJc9X1
w5OEWw8yxlxSaaEZb76/S42itk3Q6/CWUxJO7x6mY6TAA3iPae/LAsf/cRPh
+ftTkm4vEQm1RVDyFF/QEvifLFZ1a8IJASys2T6gmDr70VSIwbGAigEakwdS
Ts988qol+UYbCcvNPfIJ3cGwYKP2FH2sYovq5/e5K4qeYilZbjAIEZu7NZuB
YW7e6V2uJQOWr19B5SO4IplAKqRnGMx9hGvuKHnblPLKnO9WPRXWDf5xmlc1
Z3Xy/TgMDnkMi+PuL2QerLs88EKRzLqVLOdirluOXKPKOZjqZ4mX54e+/U/c
eYvUwiNoQO9Cxi4etNzJCC5njhj+1tARYMv6eK5XKtcrVZEBXvCBEWqCrsDa
jqlD/NREY2BmfGipbbYBKP36r0ZwOrfMP9XWPDgyxp72O97fQW/OBur8/xzp
tMGz3ziunZfD+AujL1VgbaDfsp3OlOduBdX//rB7+BAxIkUPZJ2p++hlKJvQ
k2euSQFlqnnmGRNrEknZdJ/fld83yo8f7UdyKRE4h+1DnCM+ufK5NYJiD5j2
rgvViTVa7oqh1EbP0jN4wf0ThlObZUCi89822UVWfjugLeG0CWmGWanUJl9M
jSbcmK6HA6hXO6RFFwcIsKIcJuRcb2fpSLZYaINkkOmBxdd4CScgM4kr/jBF
TQStkzuv3egTFzHrFsWrsDUlIVXz2OlndxRrk+DRS5glyZIQ+nG181NhHHLa
8MqszYXxmOzlPrXRnLwXMhvVNayhIMxpG9ml9S7uq4n98jQGtiwKMp8Fczra
KNeYSob1iX+An0z5JUQEeTWe2yYdhLS2XCh0jqt6ynW/WzWzSEbMesA7RwnN
Mlx4V9sgpn6qQfc3CdIEYmbdj4PRZH7EDIVu87461ohzctIRWP6tf933JIYX
raQENXTW1WVIEEZyTxHv211po8VbKZh6LxTRLs8g1Hw492YabwMwyuuwzv2s
z8cstMby17msaWcfrOakyOi0uUinG1gQJiXKg/z10ZY1YXVhBtAWeAErF2I/
l3UFGU+C3aGxXTWWlv5ID2Rd9WZnVvbvcRsQQG4w5yLhltZhvvhj4G5Cfs8g
souhfZGPsfPeEZcUmgTMIGzE+JV+u+w6q2KJfs0ghe4T10B83ahTv/m4ZbAw
CKdCT1HYQ4wUhg+C8FwnTKkkRnrkrXbsiq1yQlAx7GJUPbbpqsr21jyC/+aX
c6VU4iIlHguA1vGYXPozGYYFatCj01pZbuGxBgbAZoFOrBXFiuk7vC7wAMMy
9bA96hj+qWJGAHW6zhhFT2XCVZLbzOG2Ho+9Ke/u9DvT/87XabhV1w18odVU
90mssPUc6fPXpKXmajAG7kY0Xg8oT7VT56IZTe9lxcL8aLO9FEK3qPLmJlLC
5xlgplU3Hf4gjgYINwFsqxztXVUBoMY6N6/COxqqzKB1v4UxhTu2Lw6kwR/A
e62Q10NtwMln8qMK1lT1lA8drX26YIStdhB2PnnA4OgF46BC9A3EsmcOURVH
oW4xWCEMSOSSzFthNgi6R99KElGafTRdwhpDgvyshF7KED9tAz6ndmT835Ni
fsqmKfNtiudnccuXdXNhA+FTjjfWT5wnvhBuCCcmlPjfzpYux1nnyquxS5yc
3g2aN0v6vKp74hiP2jZwZ6lrebOwKP5CALpiGMKMh9KSEKHV8+1pekSSqLpc
EHKhTOsVMOtPZapxxwHHC4GlmPPXaxEdpzTh1hVOgGjeNq1XkQvY+3+z1XEQ
5uSsPvWbACt+USLHY7MEkR6RZuCD5sEGJzVn0osu2Ea4t5QKR4/Ij+wF/LC1
YlK5iYvV2TEmIp1At2ZbaBghlK8mK2ODCcTpg927rSYXjZYmZT4nbctEPqoX
IXaaESPhgOFwHeZto8aQT0PpvGhjWIHre5Mv7CG91udROi+XrThDxhfDdrz7
dAtxLJ/RWbi0pKllEZa/v+dWiBOFfYm5CHl+QV0m2kqx8gzjxJWMVt3Az3OR
zcWYqgVFTkcVDyE6qvm6SM5TuAzboRlY5r4O7MQo/2Le2YPPwEFCf9BatzHf
Obcd67BjMpiWZNwH3wRdaNs8HjMO5wuONw517Up5Oc282rp/QbS8n4Z6/TtR
j8ZGiDtYephV5iQeZPA0+fypul2a/b6jJ/kvuAXerRF/+01pHaQzS2TCX/Ap
y3sBSQLgtyI/1voH7b1/Rz/Tzj8fIlzGM/NV8v5RfZySg7fLVCX8WXIm4vfo
G3MDpmTNxMhI2BfDkaJhSgbkZEeIbW8Wz7Fobl+je0wiXwqPCtMr98TYyyvK
+6njrIPu2upyxVJso6CnC/sQdR2oI3Kld8FGsuj4RujfSyBBc/PgYcEs7Tux
KgeI6rhKCFDBbPQfK13pw2Mdv31iTVMalR0k0Fv2BUCP1BR8ntc9XtGv4fTv
PKOggOymrKRAVrFzCWgmU5zPY1gXlH77SQwnzMrZsjqZW6CrduvIEPjS5EML
fpuYC1Ntpx56nwpTi3qqLw3AW5r1rdjbpIFZZ1qrGuMHXB6zLBGqHTRAd5fC
o++QFIEK90mQMLl7aDpZQ1r0aU/w5Xcc4IxZLC0bGwa+MPmezzZlkFaL7XEp
u9eHGf4Spsbuwf6tJk3uyz42gnodac+H5IPMdEhiCAZ53d/GXrNy7un5nn/C
Jx7975764RIUAlNhmWDm3XKRQGyXHJxEPMY0HnVzmw5bl89JkvhgZjnUym83
gys4c9rm2bv9le6w9/slzoSaARRY9eFXOeC1Ht8B9h4mmw20ldAbjbja7lGY
jGtnsbdd2v9O/cFGPYUeBe+uIZ2mxWVY6AfGxSigIbTpAOYGPPRFBqD1qdE0
qCIZlTb39OEDWEHmRwnYWcki7x76dz8GQHizPZidvc/cLpLVvmtAPTd9btI6
lJZQTpQSYicnWXCMyqg58r6TwToAZRDrMzL9Dr31DY4c6ANZC8RGKpyxZRyf
22r9UrKJoQYEg6DDDjWXLOArBrPx6aFUqnLCdv/1xdWem9RzfflQDAiEZ0jQ
EHyLQ2nL7lTHmTCzG2PRw2rE4zOYmlcMSbNkpbjSYOVjSF0oYgiawCE4dk0/
cK6O7gKQkVXyGgXS90zBLX1r9q5fVAR+GXQpuMf6PAid8gOqVjV3HHFwK1jN
cTVLReJBsk4r3Lu1Fgxq7vil++Qs1pxhz2WLl4VYw4jkK215+5bG0SFciWuE
g4Sac+ixr9Y0azORdz7NoW67JIC3UEr/LHXhPwO4sOpnVjo4F9109OVFkNCs
ElwqNr+5u/JxaUomcRr6i0+29DusthVSSoKu674YSE7cLVCH1xfesfSQgA34
kVETiav2bLnJOIo7K7DRJ4G1OV+7knsJdH/0cnkQZG2GhhZPKf0XUtHyY/0B
fPLrAmlQvc841OnG2fhIq3hpWBwnvpkpI3+gNyld5CZ0l7sVLynFKknzjgP7
lLe+sPNhn/KGAduTljYFI3a9ymx3CFczsAOQd9ZT18CD9S1xbbk997JKFolG
caYZDazRLqV07Ul6EQuRaPdGJzr0mZwSL1ltXLsn8eDY7YU/3Ur4p1EHnI05
CvNVC3s19mti/2RNy5S22JvSa1/nfKkjfy/SVIq6T0k3ESibm4K6oYKagYn5
/cBgO/rLDP9BexvSbCgFf+ETWXlyN4gRYvN5f8u8vld8wEhJ6o/bes84MNKs
+07G9Z5ZIFAQuhGFqK73BdoRCb2qaoWvJ1Jk8gui5/dD9m+1lARur1/CwvV3
aESdrC4OPSPpI1CjakDqMPRcsA8nJty34qo+szoMlHQ6iBuePzSIqfio2naU
2jnTjaKhkOvuJI0OekbJ1W4bFHeVu3lZycc6sTsZJRgZk/ojuodQGqXXzfL5
7IvSVcZk6+SQmW+96tQBiQ1evwJl78aRO6iF18W7Nyan7bGnusymSK9cas3w
k5hbfKBCkxUrZZDv1YrN6vEIAeeERDGIK/hsX2fF4TwQRyqqkjoPfW1gfULp
rmPANe4Tu3L3OS0oFYX4cjat0nYNfCAXNXFjwkLQfC/9hI3OyYkUEHUeMYX2
w9Wogt0kAp56+6NtFiY9F/WqBsprRB35R4byh+urHKbnSQ3wHgjrckZrTw6h
GSTyHpJb1ETiJZ8immkCkBPfoMdBZHQ7w0yZslrrazqwKkfRgKDOVP0Qbrm8
UVtk0DEz6P1zqSZ1ukiwUnp+Q0ZG7fSRDYidRZ8BwMYLPcVso1O2Z8+z1sEd
zSO8zc2eSwZ4rVvREyJhLQ2EgPxO5tLvnnvOwxR7+9gB8kkLE5He11T2GMAP
rSCsEpLFfdBEeHo2KZlN5s+0ZopDWbV8XuvuCqPodZ2bNHYqrfuKgc/ttjms
tbpNpxWONiHzHi6TcfriqzI3frowY0Miu68Sky+b+fBGzi7n47IU8Rw9O3BK
5EBKjZK3+SLA5D1iT+ZPok0SV+xt5nL7noFo0JK6w3sPZCckZodQkG0fnVPo
u1WxrDb7WDjmjA9fvyFAC5azBmCULpwx4+jimw+NRUwYxBz43BvlvQEYxCUi
u6fZFnq7MAddYUAL5IqtpavdVqDb1xzUVi32pL2bdYaQpORZcMVMfPMCrsr9
DT1DtF4/oVcvN3UTjrmKJIUZ01lf9CnOWuh7fl6Ru6p5LhNt7c38dZziI7dW
8egmRD0rblQsON5MnG3ppLTcPoT4WIjH3PxN0V6/mL8Gwni3ioM49sUCUSg0
ltIYHWcQZqXItQ6gTex1DIrz2ezhhVh0ocHm6rYOtfwPWRzHQJAfiYkDQ/Mu
vIDtRI/ktyOz6tslWV9Y0DPQSnDTelv3PKUDQJ5Tms3hPwblaYAHWAAJX+uy
dZ4XxtOisOsaULii95hZ+IxRtEOt150Z68EdDMGnA0uUeA0GkJyG7NEuJ1QT
T4ZCgM5RMR9TnU2Rw8vmP2EEPFt4lfy+p/4d2tsfwu6dL5K5rY/piypxlsGo
ImpoxOAXAH6icYsMndv/itiqVgdHJemLsFf2OlL0F/xz87rksh5nHwDug4/T
J0JUDLWd4RZobIMDFaTxmAnF3hz7C4Gc13HNTp7eaA4eYKSruQRmiVwTWc++
c7B99mBfyId2LyJSpCH+nug0ap0qKAcTFDe3I+1NfzuENA4vV5WDmfcRLLZD
fQafw7eyrxark2M89H99lkwyEncSRVeaGfDEqha3UOGV1Z4FyOsD+KvzYXX9
1O3xOuALKK0Q7us4I93BrE/C5c7Zpi6+eMJXHlXBvFr3IlrVuNnsFQ54ZUnb
qehs1qdCqEQICQCPFrbS2PA6Y5Z2pJFUGvPPvRVIa3lYdpvYk3SfWWKat92v
FeX0twvzxPVEHeIZ60PeckAGbYZhnysDnBssVW45bqOBvnyv3qIoc9p6dSzW
AsptBw0VsFb1l1wqkngjalno/WSkizaXkoLNhFyeFnG85wSuzkZ9im1+6gAh
NYu1nLy1pgtliyjZee1U/AtD87qNK3oH5fj9JqL1uzpFYVwxjqP7Gsogf1WS
+7cQ6xWIhdECSyZus7LwHphG8kVwgZlW6fygIjjCk3QOoT9yA4wO/pIuWtdA
YI23/WSoEPmjShwyL6EqdduN7MnXEYuaiQARhIRN46CHSA6z1Go2TpziLxa5
oQj/nAqWWFc367gd5gGbipDioBdtBU99QxnZCNyEggSyjOS795H64gO+AC4d
M3+If+jPiKPxeH5FX2pJRA1ip9TXpkq5AAZUfm8oUPiWMJGrG9jADFUXACds
f3wGUCPj2GtEDe8YKr62o31LndZjgRUx7EoSVu9AA8VlN2QSyjTMRdO6SFRb
RqJOIu8ZJCeXHKLIOb5YCYIGASz3doLTxvC+o0kFTr0U8O1MJC0nj+RpYlJh
9/2+R8VMXnRiiUPzbMc1vX+evug1edSoHXrq6VkFV/n86QflTyDwv2Qj71Rd
oNspRnOdkwRyL/J6FTmAhppze7G+VSIN6Sz2HGmTO0csnHAKYFLHauBYgS0P
7ZPy4SLvmvKyM+eA0JI9jckYPC2POdtifF8lCgsSUn0RuuK1vd+pYjkkGAW+
ENC7U0vniMXIjJEVDrnSeUJx2PyKkMGoyTPVFB0ckpOE5Ki/i9UtrUwe8xfz
MHb/cLJc3ViVf9QjHpi9YvFvUuBgIrkcvEZoShhJrvKwa8ScWFaXZVZeJ65Z
dIqwvSPJWPfFcRPq+wToEWrKVmH3WkcDBkwIc073VMyjhZMiEyeaZvblNyDR
JQGco0smgTgDw/5h/TZhpoiP4oiOS9zWuR2MZ7peN7jsg80Iao8+b9i55MCi
NdRqBqHY35WecJtTlnhlM/K65e4rgmQ/WMstzTr/jt0srUHI4v0oXbr3kzNx
HokWav4WCOC8jRBCuxrvTw1sOg3ncDoQMbWpicZqHqFUkESi1KmXCE4Gj67+
pDMrCjm5jsjkIf7n7YTP4+7pRfZpW+skpH7QiNLpH91xfHYLtwO2zxpdItwI
PKOO7EedprxICFpoMh8IBHcFvtdEXCDjVzKbsJi2aSQDUYFhWtllw+fO1lFU
kNynBMcAfx3gXtUOTC2vSbrfaHPBgBUAyF084gl33Hvt4sBnbIoLEm9Qzz/8
rsD7qHbF9oBA0Tlri+i6o/LWybqajVIEgPXO0UfrcUKXT2P3UpvTkhnbIVHY
fuPu84Sd9CluSV/yIQd+oyD/JYPoWpWMI0DFETPThfuF+ktzhnjOMdqvOZRd
4LhTRg5iKpn5hUytsWO4djOCxkq+J5HF6NbHSg1bPGSj590GcB5X08YHMT3t
aWHcXxhvDWvzc14juKJ4/NJlyV/+uJMeYLw3LcE3MmBTD7dTk5NfQQJRvRB4
ppWRrPJNNwyPsstn3c5kAaziQEYVOPcq0PYuCZN/WKIlZlBnl0bVTyUp+GHN
YYkI7YZBmtzX8R0hrOWclvv9uC4AEKnbZvWGMXHzBtx9Rz1anRKroT3ZjfFS
Ow9k2hOM16HGnrdli4zJqpBLiemLcpUM5hDXN3ilk58FGOWFQvMlKKYuMknk
BtoYfGr7vyIFSS7lI3nrMrQ9D9OUocOqoT2vzYr3Upow/VUT0UiOyeUwfnDi
Uq/0O5GlM/rc5MLHyCbJzgQNp8kCV1L2RhDho/0W5TfcwjPMGgDsltdBzHHo
GTXAAFt0tvVTEP6gC7bWXllbTNM5rvVIPtyL6j/rn3qMjDTWVhf3tzqvDc8q
nVt3/71rQWAP+Pm3jzG+zfuAzu+iETEzz1ieEVXJ2sVl+54YGS8mNKHqe8Ga
kKwsP7lRRCH/NIFH/Mcotw94d90eN+u7FI122wMmJHvNw+9GvmnF2vU4i8Td
IymI59WdfutnT07lXPY1HCd8NeVYu6mLdJFgkfmPZBUbMgZfRAGhqZSG0ugB
WjTbZAcvW/lkSDg+QY++jR8Iw3cscGfSxSujKCftWilVUYNW3I3d8LH5Tfi/
sDPTW8fEjYyafnNPHJrZNab0Hgl101PXxkeSdSr6u7Hfj8yudpc8QdJD+vUW
XurGXlVmNmHQstd8kw3iCaZJS+rotUystfyCwXWQAKqtbwkzXzDwYX6V6adg
VcJ4Ir1KiO6rxbnPrv4vGtuc1eGSSZ2jzM/9sObEGYg82XobDhNYVVHRsFJV
xNiSmeIFr5kuRhTqxvV+I52I2e3D12MXb90sqWicwmQNEn7D5h79UJgJjfwS
t9rb/mhDF7h2hjqgmoZ8KU7eUfDGgNj+rmNc9d4qLw2dOQ/xXNzhrH+wXWJe
IbtOLsrip33bcQ/4MgXAIpogQilhWh8RkWnB91Jp1y/JswDFq90yJtIEiQbJ
bVNXoJwEMGjJeATTUeM6UBOYM64+7cv2XoW9YTSSmIKstlYmk9NRSUmOvGmi
EOpu6PcPvCp3lfBXkj6Nezjm2xl5JKEOdTCYXOkoXtsdimb+xiZ/+K7Og2Ld
vbCn0G6UOj8fQYaYnB/XSF9+82GL5mxEI6kO3WZbBBRnQ9v4aG6Jb3mlWAMK
j46BxqW8G8Do75iDGgL44Td3yof0bThTYgI5kL83t1LpEMaq82hAyFcLJHAL
HoYsnvIqO89vbTOiTmjXjVJ/W7WUw9PzfheKmoKqAlC8d2e6OJ+YH1ZX4wCU
Z89BEDMqUpByyEU1jcFEpoHR9PvPO+KmEXU9uAixGc95ohJ1la77DVddonCQ
RZdiwwbWsR5c2CHEiNlucCD2enxbyb2dMi/MHd2QKfGmZclHJ+CrxE4XF8CF
kLgH/lTJOFXhhgyjrgZh0kYiPWuLj7rZLEQEsf76ozbCIUQSAyJrrICHxZlm
zyK8IjHg76qTVtPixOhVR5YjNORbrbOErXdSSPnW+03NXlhcuNcvF+FiUW20
2B00kowEpyyr1ynix4k9qzgY+YL4WCk139TTDMZfdUnjA4Txmaby7qO2Gb/r
E9gRpWAMR4ZvlxSAK9k8CP7vRZmZqnloTZlYCTUHTVTk5RZqNsMPeX88E1+c
GReVpreYQQBSV8ssEJHwNQADLDp2d2CDyjibW45b3TjArBYVEmVcHD9Plo8v
DN5ZagsQp52fT1mBJD3++uLhKBWWHEAq9Onr25OBhsUPp33wYivlZeIZjoyS
Sr6D75y042YuyKKQk+z/8thbylfsjV4jAZtUK5VCPl0HyIVMGKrqJsnGeg90
qmwyb3dMLeED2RDF7MTeCxqTVrsWUu9/WM/MAtwXECLgU6e6GOmXNpuZlfL4
3dMZ4OFqW1FLLh8lFCMc3kEOy96ZrdlB+G3XfTiV+hupiHFiClnwttz1+88u
9fW4IGSgSsjMGcdUcsvO12KfcvV6aWXX3585ooGKDP5TFzlPWhCwTzwDoIzM
gEaTHRs9o7iyF8PHWbzH4YqohF7U6MWzNIO6Ash+hUMxEEF5QcqM92GRSmXl
9yEqENnaYuODgh8FfBzcle4iFGU48kiBSeO+vMnxvvFHr2kWy/UQvftB3t9Y
dk3LQ4oID0/fJsm9m5Ff+aroEbaBybWfMIWOVh7fLr3i12yyDZylzERIhuSL
H6uRyEhw+Z7Q5Zmb32MX6LAoMIXpBp8Veusjavd0368bTnU87Oezb+Afmohp
bXgUfZ7sz+wpR6CWw+iHVsUy4SWgS8/xH/CpYfMZXQf58+H/Y+qJlWG+Bid+
wISjzCGhiZmiPRUGigIulen7XOKoEANh1iWOaLX35sI4LGFGeTJF/G5ki3y+
Ww2cNLCXHNRiKVB4QUqdfPTd3hNbJyncCwMySG3Lymwo0KpbQyU9KCQWUkar
8sHpj75dZLtl5np6lYymMiNic1T1eVTYuQWkP84Jn0APSV6OWrRGKN454LCj
yfhRvyVmtOBVu8/sujmOCU4nbUzGJ9CKC5PP7I3GVpqVcBMhD/RWprfdLVeg
kIEPh1O6FPBoEJp1yaKCBY/E2+aPuGKxAlOuU/d9VyUBIopNP1oGuie7AMIu
NFv2yTR9p8fmamb0wXxJmE+lHVXIzb8XwyEdkipIokedQQDCl00jH7UKFtHM
Vtl7J9DIx5SdCwa9Crqof8eQszKWUq1s/h8ZJIEldCyizYXTCSgsiN47yNID
2d8/QgiVI7hbDbO2K5dXel1TrDzqBJ443DKYximGyi7uxqYl6irqBqants2z
HKBgmk6PuMrQtj9U985HqNB1Yqyql/QTh6FofsPXZOkliw4/De7SarxtgEC0
YaMuJ7MLux3tyQoQ0gcMjusIFkKlBr8w3b6NMg1PjfFItxzGiEDaLpAnqiWT
DtFtLkxEYawMq02ypGbeP0PiaDn3RZU775IEXubGu750tCuJxn9We1Sg5H0j
TOyoYi2aZ+TZnENWRS78LEy5U83dplqNo6WUqu8/dccY7CEDqKCxrAQWouLY
XI+R4TxXRw2SvxoLO+W8VUsebhsHSssBN8yjm++bE+P9QZxB/AHZJVvcIZ1m
XqIq31TQLfvjIRmYq0bJq/H1hNo7845Kx5q7bOi0pAh4jraB5lMOOr2SYqzp
NDokreoP6InJjf36376ngCZ+t7bqdyVV6REezhFZDwt/ADrzA7g0kTO7NscN
JANFVU01UvaBRSOpVoIIe0GYn5cwOwp589iA1ThXe6DxbyMDS7lN0EZ6i4nd
Yi9hDmsqlDUh2VkJE/JJ+jll1qNWgsVqByvfTa8b73bOqyWgmhfPN6euVxhr
t090imVOmu2W2WMQPDB5srRnB3gsfvc9UgnHKcTiog+D2rVz4orgWn91/VNc
hn9CJ7WD2w5G8FtQci9jW4vk6dGxCfOgcntpJZLpadPPjjw+dEWsX1Oti/gG
toqT/++dA1sWW+ItXFmd6fBZah8LN+hfNnS4o8UPTBcBhGHgwAioyAfDa8Ru
RZItFyLUBldLQnGtoJzNJBCl5bcKU45GIMrQGs9/0XvRuSqfMboRZ7iZB498
ln7w7FLmOAWnMWGUnfCNNYkBmAO/VF5jQa9A84aExvua7y4fVDz6tlXUxzcz
LQFRUC6YZRLlnIDU2gb8QCuVpI3kqfehZPwtERA10QeA8bT39pWIZ9GQ2aV/
WWfTk65VLzbAGq8WK0CBZPKKgy9vYjAGMtfnu2dvTRDzPFc9ksZcApU91aXX
uJmwsxbaVFf/T45wPXJ96k4zFuMOc9wQs6cboypAyWuqGbczXQzVfZaXP8PC
g48ouoz608CEaLYXwvv6ysAt5DO2Cu/4yZF/vxvioo6/uLnX7/Kt8CsXImjB
MyI0mXvK4sk2TX6zlXTDfxjeUeJjk7ypGuiXTLWKeGdl1BKR9z73XO9WNXvu
ntQc7JF12WHsCM1Ka+5XTO7FP1Na396Rj27B7TKoTt4ch5/640KmCCrM7Zkz
2vtc5fWyExELVM91ctNkIvnOfRQ+y8bY7qIb9JjE64UkoG0rbrB+AliBiJZ5
NumvhCSWRIWk7zvR+4n3FH02HFiROgvp5UhqsALUh6e4gabu3lPwjMiFnoPo
PogE5WqQ4QKCRo+hutJ4R3wQ7Ov0am8FHIK6BR/eUDcQDYosm9kMfPRtNh+g
9MK36MDLGrlGo60ORV39QzwBysEqpMEoR8ZxX8X2PdTYmMvGxWx6Je/hQqp+
u+DKucFPO+tDrQPXkeSi29ZT9KuiXe+qR7bf/sb53kqaxeeUUgI4zD5zxrpq
10dgXWp574+cLLPyRaTYAELNYvnUFuLX6tTqNPLWm2xK225tsrcl7iAmhksb
qizh6swcl/c1ZU8UczR0zUF2i0ltxQZrA9vHLGjDyshGTNHdn67EAC7KPZD2
cEmkT6EVfBxOqSYR+YE1ud/JJONzXdB/7GAy72P8MWv5m0+3wkpkHJw0/EBS
29aapTiGRxfUjrjhcbMcutk2g1DJ8y24/vvHDxmBniZ54jzXPwiGS1rZuP4X
B6KcJxR9ZtEPQZnpfT9uXpowA8qkWyBFnSERhM9YzoyIychpAL9j5j2hJ7CP
t+T4ssBoY3b0bHC6nLt0dYQ+uaMNcyFPFL4pnr3+jCKyixveZX+J5aPstBSk
Rm3ke6SkZ34deNHYLHRdRs6kaSL8FTyJ5bPZ7cO24dNtSZXvHod7xoIZBX/U
opQ9EN4sxycGe5N6Kzyr0Hd+Nt1zZFsoTupXR5f17MaU5J1O3KZoYE1K2VeA
eRH4OvcW9LAH/hR13ADeG4ro4DiJ2gfoz5t1zKEbzyFsesM+dhezemWwlvyG
utmg7+AUX6yIpIo/jqA/ZTYAIElJupRi3XqOjVnSn1lKVbeJ19wUCW9I/f6s
p0lRsgnXij+9I8uacIDOo6lW1iugGTJw3tzytIhRSE0ppLhtff+UOCgCTg0O
4+d8QCpMGra4qijR5OxLqsKjFAPcwre0DRe72PLqhPuG32heaayDzDit4ccA
1FMBJvbWvHna2pUd4cks3svTpxrsAdQ1rBr+NYfMpfuNZFK1MkBRnECB0IKA
nROMrxICwJykDt+cu7iy2tYNO0hjYFM+P6QRNASzUV5tkujFehT+VsjrEfm0
p0hFZxwnXzTYXVM127qPVhTGsMqIAn7l6jqatUSC7j83a99nV57hBCWp1hAX
LOjwsUgigmxcyA6jVi8QD6yWrNH8MAFmNB7/O1F2UUHehEERxNkT/bt8RB7D
TvA4hbKxCnAso5D7ElF42WbbvDHWNP3Hlrke57fSjNfKO6A5AiL1Fqwp8OdT
rkD+/Ad6Y0F6QzcxOXCxR27uDSKDfxLBmxZZ18x+JrAAaIMpeVBnyeyRTmnM
XZQn8dfgyCCxEZybo2Ndootgfc/g2ydLqo7K81tpijRq/ALQDceidD8e9NU5
KFnIn+rO1ygFM1/sNVUaXsED48H/FEidFmlD6ojotV8cTHfRu3j/rrTJB4Ma
zmIanllKj4wnob9L2/tHd7DdiAefqGRY/QpmhRT8DXvoi9CPSMk8QCLN99E8
TuJUbIww3l2IvLW6F+XY6fL4N41YUEK7epfnaaTt26qktxgVZnXVETKz/yxH
mydTj+rtP2FrmngvZvA8yjE=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q5YMHLNx9V5HU4zxD8Z583suv8A8S7RMtPiz2Ty1SSLRkzFdthnwvWKzPhVkdqnJop8MfiLtFAOQt/hGixYIMvNg1Ob8xdrXx0Kfjr3RelvC9A5SkwnQUdB4aV1/sm35CEpYCXeyt9OloLbiL68r47vg5ZaKL/SKsE2kvdDUYJQLz5jy94MM11VDqukCofKS3J/E1XvFBrBpYZj3EbYmggvroEBSfTH/r1VrqebApOqWyI9runz1MWMcygGgRvStoNmOXVFZ+cTYx+5ECJbU24KUWL8nwHphMnvfjmN8kxdGJ5hMlHtKHj/o2BCIPWV/b1jOfNmkEp4LZEY7O8hLWYY4fTPG3pHPbZ+dHUM+ynbmIIvPe5m1l1QbE1fKnIVMIGUAFSwJXn2GRAIHWUq14rlEoDt1Na/NIR7Bi1HsiTAd2KIhm0LRGDfxrW2D3u1xLXICJ7u1EIzkxoprtUvvTfRiQjRYEJvaE4QvrF7/MNB3Q3S+LEqXjIo61FS1z7kJIXHHTMZ8L6+wrhIF5qdXtCODoKol4S65NnTVyBWDn264UW1YV16QAY5QJQE0+IPlXVwD8PG9+MvG0xeV03U4cydGfWvEb3jc4cw8WKR/FpLgtmiq/oYjaHrS9hlGvlnW3S6hwhoMcK2ODbNY9cqwZK7F8qx+talXCeJOvTDEzBFe/lJ1HhHgxn3zfNRLuPivmoMFeTCgkV4V0llI+LMeHUkKiCBWp2jIhvLC/8SaE7pgpSfEIayzHBoH6hOp2TwskiaBW+AoW5D0sCPUKzAiePK"
`endif