//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
wqo2XIM6YLLBlQSEVebWphUBxIztJ1wK2ZDex3wCuGbnzsoPl5UJZHFgrFOt
lfkjqJn4utGf104CnJx668JpGHhM7wA6wLiqjrlIxdCQoB1wZWOHn23o+EXl
UP0tDSfcPtwJErIL6IQezc+NN1TDb5HK0AOOQAHuS6K0GxKGyV9Zad40g3Aw
LUgeUn+hjTqVs2l1Kjs4LPgjCBXpcEfXhuVgo/KbdaGuWIb5Hr00BZIbl63Z
IuOFRgAvm3uSYZd6podtoZYkYT3OZgyoLIwkGANk4AHZY5oWZQu/t5IKdXLg
gebWFHxzH6U8nlQud+7xkb+GNQA3fbwzO1fICPsuJg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b/icV2ujnrhJK6usK0EVpci14ixeWxoYIJMLrz13t+Nt1sHtOhfCplDZCQfe
dF2kjxO087PtiuCMtYWZic0HpMOEZ9/2gCWmIRXY1OmkJo2DPSpqYKrt3+9p
JNlOkenOlbQyVOvUnxFQBXCB5ZRUGH9uSXw0LmtIFEMqA6ftcNJlZ7KWZ4Fz
pOaTAxibE4fyBIn9HeQGaUWj7mm9DeTic9yFWDkfjOhHNTBEEfAPY/n+L8eX
Fo094BUEm9VTX0pbRQPBtuQGpB3MwvolRaAcfWCHVQZa71DW56QOw3I/nxUP
OBpmyzdttP/BDtr3aO529negRUexyiJNc72UDZg4qA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TdWCWelVO2BLEyNIpdQw+ZAEcKdpz2a2rXHytpm76cuPLCRDusOo00MnfZDE
FUIzpMSgdP0pAa19kLW0skE7yK1DkSWC9cs+1fvzVnSOK2z7MHEeEGTJM8qf
zLm7yMFusR4U2BPOqTX/BYzRcNvWmrjCrnv6vl3KZ9miZ6EjluYAPLSCbG0M
UuvX5yYQp7vgA39vPTyPcQQWCnFaAze2bNoKRaxFIBid3vMf0xQaigUacybm
fms4eK/yX7R++QtEKVZazulkHd4ZhdV6051OXrQKIlIV1t97ulDLoGkcpwx3
FzEoAlJZqRJxQbzio4YQq45m9uHxUvoKRQlhW50VNw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EMrzW651kMWnrL4iZmHmxByIGm+cfRLEpuXDchNSGkLpaHV+NFx/uImLemPF
4iF85UlHzqgufn6NFPb2Ypd4YT+RyDghgPYpJGzBKV5iaBEgE+ZAwRopI/4C
WbaTKt8t/RtIt/brB7Drpzr/N+i7D4ZIBwQL0GyPELAkpv8w5GQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Y74lxOIoMCkTYeYOojHBRszFk/BMtCnE2lE5XLITvek8rhGMEJr7cnkCDrSY
DVu1vUMYlroOLjfQLmIBT8JOBDeMEIge0m5S1+pa7nWwZ4xjc+VYYCbu3Fkk
mFy0oWyBp1E7UKOXFSnfbWBI396Q41X4h2MxrxMHCe7j0RtY9SclOhJvaX9M
vdwW0WhCBRtL5UtKGvG6yMuD/Fmra+L5VhfDfCo8Jf7ddL05wBKLKW/ILLL/
D9m/8nqOJLBIihjeLWr5LwnEE5b82RoFJ9PcALWzri0ZF0qyvPJ0eFq+eHbl
NJz1SSWkR6farqK3Y/v1GMIWGLfL3fKTwvWnUcLJyWPPV18Iq1RLYu7sEaWI
GtbRMD9VuXWRWivsgcID0Yn8OJgxR6fBQzbAjVjsTWsXB11GiZz/faqaD/UG
q/oYa4bfVUR94EVIZg+qGQFGXeURAynmW9uMF/bdHjJepI8Ja7SsgkCfKDu8
Ni2Kewii/InSoHVf6DFBr5oEbLyaL0UO


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
AP7YBfiddYGJFV87irbJx4N8dgbVmNw7N4kP3IXOQ4lYQpU6ptzTPMRd00GO
Z+kPxPpD7tNMKGRDEtmQlj5d+K72rp3wiWPPkrxAO5UsLRAkgi7MCDdKMkRw
IZLjg/mUTRkOe1C9xXG5zpUPIE6nbt1+uFgVzL0Y2NS96CWYTsA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qykrR31E4TczRKif/hSqzrWynQMI4e0Ts4yjyarVbBFmmQRaxZoZpx0T7oOh
9ZCNtE/Aa0pK2lX4j1ywlLvt80d1Z8O8z6VeXsTqzDHnLolVR3beNRXrcqlb
Z8YB95Jmin+scXwZfZQ7zLFHJ7exSM/yS0r0QM2a1XsKKC7kfr8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13024)
`pragma protect data_block
F3qEOCgfQpFGAXp+hRxkCF6BETSywjSxQZCe46ZdzvziDrV9VU4wEKaUcnVr
uFA0akns37PR7O1eV8h2ehFrPVD/9WbY8MRLU530kZI4id5KGXyLNfiNqZU9
xDj0JuJjJ0AjiY9vM8p8PqiFNMxzxsGjNm4NN6TXdP6jT+7VlyPe+gcf8LnW
Pl1uOXfxcheO0xAhrUhkwsdYnCh8+0iiKnWE9GQh4c7ty2ofnXnbuxhgg8Sa
Cf/D30FF4QFXObyGjJGVICG/7gqJLe1U13Dy84q1WbLcmYbpxIWt4p25C0Sx
PdkwxFx/jbL/c907LkJ3VBUafglHK9j+EDypPy9L0V5Gru+g98FXuA6xZPnM
btlSU8HHd3D2SM/fPv6LcblBfbEYRejARSvrGxpbuVoKwR0bgVpsX956t1W3
4wPryQWq/QezeveGV6bKVfpUJ0h+y04Dpj8SW8+B9zovmp2ajmmsD5MRTBBV
y5itdH0KEeMSZYshpBg5teHjEvzNJ8SeXs1NJ3OdEYU7PQsOyn8fUErdeoBo
uuO3kA/7Qi3KiGusuqF/HsYgyyQMmLCOHLLZP6nHYhm7KpYtm78Zrysbiguq
/IBhMamG+fiD/5kGxp4xVMNiMu7osX9mcvcOS/BQzj6ZhHEYseNzUmoWdEgW
OnSLmIvIHc1UQe4KL8fgpCWzPKSHS3FTEJv65k7Q38eCGXb7s4basDCUJDG4
Qkn0qE2MwvXvcFAtZ+bq5WebKfS3C15FSsnB1GuEG902x1vgBWDNHmnGbSjx
E10OGajbEYkllirzqxpeb54bd469KYD7E7C9Eaw0Yny/yTHfFfBBh9amH9ic
zWHDV9tjiRJUIoWDvpPu5T7Aqxa7bWK+UmacIj1QZ4TBBPUoYVQmBfdpcF59
PmEzw7pD4pKvtyq6Y7CDTkZEGZ7cN+Q4131XO6xLVTXHjKyzzhJ0sPyBysrR
Q+A/Nx0bOZbLlC/44NpQy0Fec1mDbeckg7RuK1fjp/H3kx6YjJocB8uG/VcC
MYbOtt83Xqozy35OgOozZqgOLTjAWYt2bLitCSv6arDsrXveOhXG35yCeOyT
Mfg9QUlkWMgn0U3Hy23aXz4bYPYjpI/+O61cHfxnjT9fB++Ji9P6HdqIYaz5
6CHCuwkJU/5/JyjRjhW9MmvCpGxWvSzXAtro5doFELAdoGZ6SkEEnbEFXj6Q
f6tn4tFDkSxgnS0GV1xBElioy9jJx7OCbrLcdlzzpNesL9lHYFL6CjHCjh8m
rd6xGnO8Mcn0o6P5rC40YISeWJGgX9Uej0IQq1KKLAiCtEtT2Cfx0Qxs0olL
B7D/GPjuT/Dv/N0ZfJlQbTbAVxNaLisYH52IjKd/wFkjBeiIHAxocchakD1J
JyW60DlJy8UOKE0MnZA8n8opqkDLFtkE7Ubhgnhdp0vw1FaU5G4D6+s0NrJw
nL88t2ZsmxGtYbkY2y3eZQXw091d0NK0B//l0laMoKT4bqhfYw9qfdmT89ZG
7C73h5KVTaRw+bViUAbYzfDdRDNi4hH3krQsQRO7tbc3CVWWeFNRyIqlDFle
G/hb1D8FINpmCY19Y7otZqvIosB1jrq0j5VOyTn5WTnpl3GCL0cP49D/E33c
VEWaAYV14SuHAwi6oEGKHEUUlhMY+aXcjf7TZ030y+UFEqGuDuRhAybeNhfk
COAoEVf5JSyYj+6+5SVL/N1y5yT9EUYOvg+9++OPGvVljOJxYwRSJQa+keZO
jVswvsdfxPXSeglkZ/dzMaQ5anGhUizM4HiLdTTVW7c0drhSjbU9B6NCcYiE
4ssI3H3W9AgVbGo3PWHyV6mLcJh4dIYYy34f2X/BI5dONVZbY83H0KcMxbON
fhuQq/+yyuW+y920inas3TFYTBwqakiDleQWZphxDsXOBfYK3YgWkwdnIGpT
3dd8DuhADaHypjz15pUJOq71TAS5ml80W46RSP5smjx5N7BbPHIYddTpOxkc
06g/5vRhXDroKXCr0NUKqPJsJWx03v3iQuDHI21LnyY6ukeuAh+3BGrI1GIo
+Y0CFcxBi2N2P+6Rrl7UW0jtXYmmH2nUuv2/cXRXx8J2lTB6Sni/MhAfktLA
zx5zuFWa9LBRjORlpVeTDFmhjTxC/XwP4ZtD9etcTuK/habeAS+yhoYdQCBl
LZWGgkcv/Qgb1yVy555IHmg0RVbStViV+nnJoUevsJ3baZqE8m1xpZXb0Djq
It1/AD7HGBDlqTNcwNv9n1sXmpiFLk676EK7uMXC2JxW+ES+CZuZnhaDAyGw
pCoMpjB4gsMTIQicpX/JYhWmZmwggK4deBlUeIDBpKbiUR5MJekyCatXJO4a
dDuZn9SxI71AhHiHTDST/KfCfSZk3Hj8C+vBA/vYPobTv967qv9QIeD6WMdK
Blj0Ldc44m8rSgf7E+0wCfRmDhgb5ihTWmMW3be173jweSmAF3Eh9pT1hbtC
8921bAO96saGzXOYcuw8bQQWKcx1QP22926i67GezKWF0b6E/MZLlnYLU22B
pKs2vvVXoxFr5jYITQZUiWQTIWLjrRsXF0PIAWJhgYBD8UAGk1NngJ8zyi+4
LphWOu4g/T06UZXynM71etm4ait937wh/8kRL5N/UPeggt0VzveqZ1+EMf/+
BCzTaLGj/QQfuaUYf51iR1i7+/Zz/aDP8adIjyMZgFzAc1JJfQkDPBJrRZPL
3A0o/Ffk+Z0AUl+1PsJCpKTM5JuI81nJ8t7lgsvV9TydPlMIXvHjefv035O+
qjjL7BKK+PeyN3JxUtqUXjiPLJD/dC4fpmAoa4Qe7eqfa285IbpflaNgvh24
RzbZF+PsJH7jaG9sXhElfADyoBUvdeiKI4Ct2sq2GOc4LuWimbTiYbmebWmK
2XER7Sd09VXDvxWI25BFOx1IR4rTcm6It72poDcS9843fBTAr4zy93EoTDMs
uLjszWSLkljAHmRv0yZk6B7i71liyFQdD9vyj+t4oorrlJPEjHaAghxEh9+x
82cVcfK0RVaYMG/WVqRRglui529sEkK6pmL5oZFJQ2C7yW6jqh37Laslj17F
82geKue8oAfMxoZu2RXzq1qiwXAljPIZl6wz+OG5QwgtkG+CpkzIqkndSkA7
b+4kY8T9AFZP1rX9hHxJ0ZmKDSrsqHSxF0DydHfJECYSRo6JSZb1bVs6BNKQ
xJOm/t6Ww0dMU5QkSLZm3gEI3SU/zC5/Hya0CqVhwDSroMU90F6GQz9yZfgX
sAWluDCp5xeJCSkAhl/sr0qN2QtM64k9ylsfQ2pa2p9J8ox8UYNHYo0iCpw1
1MwtqYpE7mQE58l0YTDoJh/h2m38VAh7j67aHe737IZPpmGAZ44YobH89vsl
2VL9l0zG/du9Fr8+yn1+na6oopRDJitGM8InnlTgNZZ+VpaqAlWHgUzlZ+Fx
s91H+qGWr01jhNykNQgaern8qHJxq1ZN7X8HapjxEhB58JYkVUro6IYL27Fo
rSwupG7eMc0jj29SGwP1hoLmGzoL+wMDgGKIUhn2vUpBUHCE8NE2XE3CXlLB
KCMcSM1VmD5ZBDGBVVToBXPJVGaa7yzdgcBlx0eLReu1V5BsN2cuL8RswFTQ
iCrKuhv+wKde728P56NAviRowDbkCg1xZdjWpozp8Yrhny3FNHDCTlZgjEkS
9nzBGFfwNEKgIys9Mk/FPz5KAjcq7n2QXVSHd4CtyPhyCQ1Abp2G/yT0sFPN
tol020G3dktoZiwTVlFyoNkUX/IL0ErhffGEPsH48xgHzmrxCDeJgsdkYkwT
IvCiYjOMBqvIUQ0ywMmya+udZJduGIkedT9+laIFXBcO+QQdYAvLArxfH6a3
hPe+eZmFkzBn5F9G9XICTFUYz4g7mgJRAlAc83NnEDSdcW5ghuF8KQowTr/I
Bh3LObgvxlJ3M1DsAnf8TBBQxkzbewbTpBthByYAD1zZ+Maoc0Q2+uJNIatk
AV6TEzq2u/0smgX7ePGcQ+vMr4lhhFg7VNHN9gwhgy8h2+UjHHJk6Ae50+GJ
x82TAhiT6VQptw46q5GkyifDrRPg+oiN4falOTCh1WpXDq+1cWLlOO12Hk2i
9d8U6dcE8O8YQTigY0dvl4NCTameM1Ce2tdsw1e9eS6cipHaR6m/KpMrRRMe
Z1fJCy90JjDilOjglVvI9OoCaYzvmwjs55WJEC1s+dGDo1u1qBjpDcrH+c0g
JKLvKXeNggL9bzjDIqIxVLjOG3LrJpRcne2O+wHnawXIxbq0s6DDq+2uIN7L
qdX8auQfp1oUSMWKXQ0vYwZ84Yrx5oEbpdObiS2gzw1CkL/VXBgs+eVo4wyo
+qMbilJEXB3HkOW6jAtourM982ZW9ZUihmbRDiPABbTJUXBjQeDEub9k6Y+N
KHhrCsFO6L2oF15ny6B+RBdzAQimfDhsrPoIesVNmkm1IYejfOh+35axwdDa
NkqRKuK1pki1Zb3WoO4I68Eb9T+XuZ98KjECINR3XYPcVZOOsWXfNySW9e5Z
ozoxzddV7KlJyg4aw+J1Otdc2kK9mC/2qcghgyyFx4iFK9ochgUXAruUmzng
PNwjdNPztN3s6T7BFDbmCoS4cmr49AesKgi0TlGC1dw/b6PszUY3bd15gtMR
PKsXj507RMK3H7YO+DiBC+MfgJgxax1/8NVLXfVX988ErL0B6JLFmHUPZlxG
n4VOcmsXkCN5+4xAPU/ZfL/kh8XDcGQbu3TZlfhJagACU5bQoWbaWcKywmHX
meVSYlOj04uhFcLsD2AnBjJl1g8uY+DWHKz7VVTc+2K6gnIqdYFt2fk0M05U
I/b337YNCt5S/4Z7x1SAb8SGHeoo6QhARzHbsTULE9jB8vqramfD/u7LGIlA
j4/Zbw16P8twqM0oe9XnN7aMCB0KepvNTmI2BRwJ67jrabvoJKMsovvQf/jh
QppGgi5cjn9X/OqVtskKw+1FkzMJyp0l/Mrh/VkLIjI/Lp+tkQL9VjUBPPpR
wSe12RPlGyLBDD0ybhoxkd1IVQxJm1jRJj4LxoPy3e7rh9BLKzaNCs1SWs2N
WD+EDTHl83ip94yruEO36Ye55o8NgEsm5KFEa1Lsfb4HW/zVUt50GfMTpFyy
Zes8f4H430K32gpfA82xNhofxmDkuoxSDyNTmnUs2OpUIhL8zTVVqDTQPfB8
G/p41PpdjLQc/ydQcvEb8xk/wDWcswU7Bno/pOtDXMHdMmGY2Kz9obECgKAM
pPjfhwPEOXr0SH2ZHaGi/TCCTfyrY0a0tyPqcRz1+GKdC5yzFHjxdHfGlJw3
sNpWAYHJRbmh4FKtiPC2TzgcERKqrFQtkRrzYGskC9BSM9BLbukzBWxYDu3k
ZTBe2KH1BmveH7Lrde41GiwSey8m42LKLLBxJ0elzlJSmKpvKG1zlyQtJh85
ald8qaD57TbWlH+0pFNnEr3/6NtseDHf0mkiO2O2PeI+sqpd0DMH15PbjPkX
DVOy0no+v7ER0TLyKdBQYORxAO5MVFcTQFJ4FO+SQethSS+n1uLGlvQmpK0c
ldaafUz9zm0kGeSnRxeY4fQemA54LmonHrjd7nR7bkAQOXqr/gPkC+3u6Wc3
x4sVh3quSUWDGqf+xZVJwSfn1L+etaEOVHbYLelYYCelAt5EjfQ+mGVF36Ym
GLl0PmyxpvsM2L/NNXZlts2/JP6qSLLJflf31MC9bd+Mv31To+jyOQgv38J2
AMZHSRICdXkc4+xfS+L4GbsMN/Zz7OUbBdakKVjsve7qfwVO3/wVcaqtVMuH
Rtg0ZNHtNGP+oT6SyGJacQqlpS/LnasoiKWcgMRpRfD81XtP6FqfDDA3Pwcj
CEwIzXtyeXEzUIapRJxK/Fkh+C9SeRkzfRb/8gwNgdGnpW424Kziy6dRv0xL
/U3332hU/fwkck/+lsjIL87PSlzuqQZEscvGsnXTwxXzr7ny+uunhUID4Wr9
DmxNL9aJSUTzpGAV2V9CqJZlKL9bNPn38jfrU0Dq/g33jFA3tC27zC5yy/UQ
qwvSg/+B2uA+Yd1Rklo+7onnfdxjMXAniKB/ZtfDv2Gu2eFavl4h9hRcpKGA
ysT9oVk0O3XgI8NDD1wzUc00SoxPpShhORHP2M8BoGOoTPJy6ZEW/zH0Jx0b
fS7x+P5slLAFGcB4eCJeLsdEt/TtyS+O3lJhHFjG+CDr9xzF71P1aUdK29DU
Ce63oBpFAnlj9fzJa1KC9OUbzcqrgFA5qFEEA6Fz3jKj8y6hUL/JCX5Ju+/h
TwXUUOPSNpHTsxnIEdMvX8lyzymHBoFG4xbAbjCkEmK8I2MOUBYAHh90UUn3
5IEkQ/JDmGkaploT7Ql4+MSnW7vNYiszixmveHu/vrCE1pSduw2X82KbmLI2
y2zAW4P38Ys4WfMt3cxPtwzgo8kYgEQquPvNgqm9zxNk2NoyqRQibU6boscv
XlPowJWa/Ipovdl7GfbmJezgUP4uIRrYPIRXNneigrGMrE2AIkZkm45xQoIA
iOrgS2l+fPxSkSv5TuCWwWG767p0YvJa7pn03OBA8Q11fvA4qtaXIOoszgtj
9A1JQUuEATqO7z+jrmFfWfcUipNqDX7SUwbCBiuXlp5J3kdLoch6d5XPSg7a
PtNh+zntLhc51b5TyNO3SIF1KxoBoPo3gIneMJFn5btsz3ZzsL9NWwHLU7/I
iGAWJonohCFurbb+6HJ1N92D3xl5QC2Lh6iXe6e9fDWnj9dSxdnCIZToCWcH
k25EQMmaUk9RlogFXaYtqfxcrU+JVjzl7voNhIfvZS2TUt4q+AvJpV7iOBJj
CSwGHyJo4hKresElEII0F9IQD5g8UNAOQzyhDaudSFCWh+SSsuYZz9H9CYc6
5pjzZn15lkXBjE/7mwf1/tsON5/a4Uqm+q5/IjGr0NfZihdHntJNh3exWJ4q
ruat6ocPC7CYnMAkIbQU9I6NRso1DadHfK4n9MgVA1eCBbeKUu8oi1xB6UzA
IA5+47e8MoQ9d2n6vtD/ElMVkcXvN5p92xhhhFYKkyhmWyB+c0obWh5JVFna
N7Ykprp1l1y1gGkL92QuLKDxV4NUCXLveCNxYLiOAdNBTM89eek7bZhlp68C
of5ts6c2Sgt1AXA2VbY6BuFt7a20C+hyQAydxu+0uTz0+UorzSZqXxw+Z2c4
GdSE6Kx/zLq6fFQ5fSaAbVSy4gKEepm5KgoLzQ850O646pOkjkHtp5FCgn7X
APr7zXaKcZoV9nGRBv3H/QLefywHlAGLGtarJbzgL3fn7N+VwSmvnGyPwCFn
ox7gleB++ODGK9wP1rLI8I1DJP6K/6UD5n9+7GULG5PVrIl7XnLJrqSPTlip
Nk4oNqnZZnsWLSuF+/VO6wBMWPvz6RnbfKEM+Xh0ndBjLkKXy5RPUfjwKDsf
dyEXZlQD82mrXUElXscwgLt0wUo5UCF6p8jlDZ5PRS6sCPpDl+0bWApS0Mx/
33rnx9Ha/lCR8I9vrwVtO8o+l357gAR0O7vh1kYE941HdNPEwaiav3dObtZz
nMHx/yE5KCGnW8o4hY72NAPOy+pYZ3fJ0kCJsnRbm4y4xdI/UuseNOQn7vq8
C7RTeFNtWRkniF4CLDLlorcZEnLC8rE8+5LEIw37RUZ5SqZ6FAYAxCevtx02
Bx41jV62UOSlFGUn92BEY8N+IMUi/H1b9BZv7nYti8MrfEOoQ0g0NucVitMV
0NATcWK8QIC373rQ8ZW6Zcn0muXe69F9+VTkvLbcgaLt1i0QBUTrQDKfsiR6
OpqjNFrpOH+m8SdqpKsQkxey/9B+h/6XcVkWjDYd3KkNcZKacK9RPTf6QJfE
Yr7ULojVWTmqT2J8NLk6j8dNqPVdTLnjyExf4sFvlYvO2LjBL0kPyo3Uwvwt
GRMGDg0NIdIpKgBAA4wAwbcuLFhZTkTNP16Ef0zfLBDPkzhGqZ+jyA7LC5oR
U//XMuXMnIEOaRJ2UpY97mD7qkqgLGenFbEzX9zyXyxK+VZKfpA/WiZzc4fd
MlGKSOq9FznqvdSL5yLKLyiWEJpki2xDmgis2JvbZmcNhPPV/IYZoxK+Fb/v
totfYNmqxky9ztSQM+CRILutnRep/0WkMNOoXGvoGvP1I8/FDvOQr1bRASpm
13c13ITs9QxkJBpqeASSSadtWt+v3yVG4S4FEOxvRxsCCAkbhG5SWMjOgaA4
1SPGUfvu9MSluJzXxQHJwkiPCk/7UdrBJc1I1NTsIFA064nj8GzqJ9XmwBey
vKd9uLnEiw7LBFm+EVrJ+E1cmI8xqHpHd9okJm8HwHNTwrVB1xdBuk9UyQLa
ZjA2ur/Tj76fEU8whxomatWrFMukBvJpxG9E43Xb5AW6E9aXhtYpvOIqdxhY
0YFtoDCRNEdycLilFXz0PZaINoYJLIpBgZBLv2WYFx7Ij1bcpoVY2vwhp7CQ
oFX/AIWKvRjM3NRtkycg8HLnJ7Ipeh4OqRsny5/Qwa1mD1qjTVsaY6IV+Kd4
/kPyf8nOgFQQDzPRBGMgFHjtuh9fGLoiDLK95tA4b2IZZ/dCqgesPB0pmD+S
B4EAHAfp+xfodXS2NFveM7Qym1I2lmqucoddZOgMSmp/xNbJn0w7g/I14RKz
6fIamaGMXePYUAlSjxKcTRJlz6MBRjAvQVMgyR1+/Po68Apzd8PZa4/NKWi9
JhVHc6DtlAwgv7ClEqGAII61yA5K1Tj0496ccbOtUOVSCuSddGEe7jkV38WU
qmwGng2MExdyf3GWSFmZi+HkvyCE4MHf6CRy6BsLrMTs0iCCfu7V8Bg3Aqoh
rTujIlugEgN4fxjQgPI6mbqGtEQLgFy3ewEAuJ4dUwTbw/ZhkPyQQEdm76ri
p3FnkizuON2HvfOWAKKc2zNUOvq5nvu5A6BBT6n1dF80k7wO3j84pb9zvpOP
t/Ua43mWiTlxpYK0FlkGHM1oFahokKSCX/NZs4kplpiJoi9RiHCVaR+cSiKI
NNyOAAwQDBuB4/nIZuTojWlwmryRhsY0N2bXTbGJFshdP1vhpYWH6upYZw6k
Al9MCJfEkf+XdOw29qNk3uCoLd6JHL/AdjKPcG4adY5LcK/YUBLcewd93Dw8
6FQxjIWU2D8oiwb82k4sWuSF+H1ThUyUFOvJCcrhtVNwRWmeZvvTrQpdF+wI
fCLdsBmSvJPInyUA3xwI2gSVNMu3DC4aLZA7EOVxn7kIE7MJodmi0bsr+i05
YRQE3JVZTqY/u1sAp0uTj7KS2FRIsNfKY5vs8mexNjC2/IzgwqxxFZyrNoxt
qiDO+evWPOeFrGCslT2CdNSmXRJ+kifNKh+m/wpE1XW9lJERj6pRjMy7PXgE
ByiXU+jga96wt2ULY908ZUDmPA11tGzxNF2PYPpSdT8g6twxcc/rGHBXmflq
fcwrVzTRAo8ouRlGjTeBpWKWg5ngBRQ5rsyxzNMGC/vcz/fAew5XDCUOiW5/
c2EvWELuPLQZXB32luhDaHy7Rm4iceoaYgcuYfB2C+3n8MRAg7vi1pGR+OhX
NSNgLNGvxAasY1SQhFEo+HF8ohbMxVrMcIRC5sDx0lY7O8kOw2IAjLjVzEF0
IsrnaICqv7qRtqc/O8ddRVn8HecnU+SJ9/G2r/v/BvI3egryU2cdXpnAD5v1
bd+0UeuDKSuHdEtV0FihsUpkRzolN82pVg7j9/FKoFLpQ6c2e0CiD1UFEqPC
c43+hOxkKYen1EjLlzHcDqcAr4MnI/OsUpTtdHrilo5Sobx6cjfdfc8Fx6jM
wTotMs7x0HhHepO216AE9oyYtyyrx2jAiEh0gyMd51rW3cc3wVQNDIt/iF0z
68CxJkzm/jY2KY3Wycn/UBaVV8iOxJHKmTxFZLwBjRhGl8dyTjo2f+DG+P6b
kCiRfPcUxRDRoLGMHLnqrfFMqS+jvE5jNi7aC88DzQDN7lDhsulLdMDhHhga
lCRo1PKp60lP8d5cEMQjwsd9jj+6pD7ZjThjy4IJk5D0xjuCoWqNck510Z68
y/99GSjILwLTJppsvt63a/G8jgN6eC5WjcCG2RZhsaELuQZFXItCR1z23oAd
VS2ykT/9Y9cv6Ad2w513iFYjzYEivfOxT108lTPuaRyOU1yRy+VKxKJTUQZ/
TJPGva04OrNXKuZnI/Dq1ZIN7hRbFiJm5KD5KUHMZx/ypftr9xuRrIMdOBiB
na/1JQ4rLc0CW5WKFihMihxWoDO54L2x77AXw4dmML643M0nfaD7Sg59icaW
bi5jDiEN7/eNozniyHZY6gatNv9CL9hnpFO/IEoeSdEimll8Kd6jqMME3LyR
rXQy0/ofX+llTzbDslo1+BGInlB7L+pO6fehaGn81eoNfqpny2YI1z68EYZK
rcMnlRdLhwiiBKyPfkIQUOgz5NOtXMxB4bidv7cS7b/qpV2iS8rEYIGCUNOA
xyc02YrHhVWmNLT80R8FTpsToQkxaBuLUTox+bkb8YNvlEPWtODaUZ0vFKHd
btIS4c7LUX6//0fw+3Y9StadFD9gqV8Lq93OJmn6cF/MPwMShK6Z8ZFVAZgI
MHW1F6miYipaFakHCN9IyGz832EEo/K+Yqsocoh/UO7aGTEHRlzuAAExR4zZ
QGWUuhKoYO/5zEsD+CEHZ+IXkdN2OqswQEFXiks40BU7GtbTl8u9RG/Iik3j
cNkuFry5xVraP60X1Z2KwpaOO/b2HeNvKWLKjzyzG1fb6DcIqwTTxgHOJLGL
qKgUoKVUckNh6jKQ2lM3MFR3zmC1tfFeLRm/a7nDT+UbwjaEA9DYNrkUmPWH
Q6+SGR/AV/DSla7jlaaFQe1vHFTv83Z0ZUl6MotUnx1bZ4Ir8USIPBwaKKVn
AZn1YGgydhf9o6IovW7ZJwJErr9SSPGSzIe1rV/AbJ4uL6W7W9fmD7/78RJT
Ha9rhIVtNKaJ5GhteSJukY50dP+KT44ot328KqjMLlMxAJotFCZYVxWV/5SE
zLRAvC9E0C5VoDN31R6pWV8/7X11ayRfMqSRgnuMUbVcnYAGhHKFwY6juOmf
9S0ut1mR6EPiMTIMQlI9j6PlJDmOQOyS+4MX8OFgiirZ5GUMQzjieY3Qv086
HlCEvUiEG09dj1yFcdZCQFOapIdvix09gLPsCz2wNYGPNuHgmOwz6ESlCyBr
7kfD4LzdEPPaDVlW3EMmDqSDE8xgEo1kDA7eNIGN+X+TNPifZHgdCFJV9iOk
wjcnW4BELjTOJjKBzuykXY/GeKipKP6UxfYfe+QSfJuKnM4Gkyw1KB3P77It
rAjDqa9E3BSpE7zhnknTb1anr7ehlLcD0qHuAxC6Zte+8XMk5m4aKOKK+ugX
pHdYAWe5ZN/znZe9UiGMnpCL++2Kz8V/o1xsWk/COs5DOHa94JWWFr5kpeV9
EX3f8BBX2qtlCZ/cOSkFvL3aUS5V502wGNzSt9UQzRTVxvgageCB4QOPEK5d
I/OGx0+viV4NWcZELQbfAdc/On3KVxPD/u5y8rgZP4JkI4qRjK2R4gwP6xZR
tsMEPCDr+kfpZPrx/8wVZrxOTke71gK6SUk2Ha5cAbpcNUHSQwUD6Fnvq5Ws
OGiLs5lqGSBhNvxlwvAgajYniG5DBp3GdiFnXXPHHcZbBO0U6sCMSRWfTGW3
3/R8mwLHhAlCZbDDX4gmqVMw9u46vvTU5QmIVGMzl/1Lvq7+RuL36r6E5ZGE
4dQgj6kSMz4jp4a7v5ZkP7i4cFqi4b2gXFr+C9ZXEHqxkyupIdHGjLs2NVX7
US6wqSHDKAhX0OimZ6LmmbEwHP/ea9ixkz0UeH+jPE4r6BqpPhFnLZn6TCsU
RdBJfgzcTj5P93S/JGb1XNW0Q2yLujh/HXDh+95hpqRnM/cgZEpOiQDZIU8w
TaFQdiVjyO71t8oGWeKGy9jBvQ7MEbUCG2+oJIH30yOiEZkmdIN/PD8Ebhrc
LXEKT2l5OzFmFfgN82OoiZpjGdHEYRgrvwqtw01hJMmrQpGA/rTlRlX+xL+Q
5FGmnb9IWS5UztJHB3I0r3PUScJ9cUUv0RiFe+Hlheyk4W81wgnryguWteKP
T9JnT9yVLraxpUAzROctjwyt0ouxGNd5PBtznyOS5s74bIazgEEhaflIqeDn
lxPwcMQaYL5/mCIxS9ii/iNlxqy5ISzf8NSjTKuD+ouqgpUTu3IWu9FC9pdi
cIutXCBwYI2KjxTFmsGPVuSxHXx543POOQDS71bPDkEpr/nBIZxut9xOjH2i
hq91rT/WH5jq6C0PRH4D32XLETBNLKf3ftibGcc0dgp0xR9PY6pLhPYd2u+N
XEtvlaEta3OGNOBhZYFws0FUpP2wNjReYT90PvPAjiwCkB0XpF36igHQZl6y
1Xd49KJPp19McUiF8FgUClCj4oVmoAk+sCTcPoHqd3GkWRrfmPNsCU0vgw0J
yjmYcR1IoksQmoL8jCFib9sIyHC05294RAPvt9d/VFofnbbvEKL78OiQnnMT
a3Uvs9tGrqpAPtpE58vGrQaOKVdvusxmXfrlS31nWwhM7ZB4VkRJw7J1RM/v
NlphZamYWin/7+JGRcngrZvse6P1g0IEzA6iBIUaPnb3eC2giO+JdA7Feu1v
66fEOWwaZJsz87wjBNvmhgd4j/OiuMdRrqLG8zj+nMLYUuefl1Q8Y0mh5cW6
YDIdqezhQtfAvFe+SITbVWxRl478CgJNVKaHYFP53YVIEv9Wrr2mveYS/MGm
zj6qKtnq1Eqhh9yS7M3AtXHRmYmeQH9bj3W6d/srIOeO9O5SVA3oJAH7lyF7
XzOxfQvp+8UZma6/PL+6X+ULQ/N2MXyqn8VbQ2CU28WSHyqXhi71ls1Eyvp4
VrGK2c2TmGZiCOSMPek6S7Q3fGahF5Sytzw5vBSrrzPPDcmCE9rc9r4kou/k
R/Nm4gZv/s1xIkGavTXxL6ozt0qmL4pDLOYqEOC/ynYZaiqq8aoWtrHwQtZx
e6IAsnFcH6jmDSjr7F0+rP1fnXlpOG9NXHjFSUU5ezNeRIc6k226lypsJrmk
B7omtX4fn6CBCKa+oB6F1aIzqCDrYhKgMmJb94cp+4ToSu2d0aU20VkfT3s7
Uiav3tcmx8pdCTaGZUyxpRdk8hyPdYf6BoCl/nOHcD7wDMbplK32B/Xv6hwI
HzecP9rBoCVrqk/zwlqzYYGl16dAufOn2JP3oxOtcgm5+KnzSz4G1CvNwhRs
s43iWNXpXle1Fd8t3dgeL8RYbLdvL8ob57BReeVM19hpI7MK+b1Kzg0v0Lrz
hv8pfXcyiltAKMQm/Oq6qkvShSxa6fPnxiG6qf3CIb5MLYcpzWZiXzOWSBKf
Gd+lyr+011dV6kcEtlBH3WwTaUXmA+l5Gx7kbMP1jpfPHhTfoxv8ZeUOu1BX
4lZwELnrhDKFA37js6On5b0GLI8Fs4RHHjfbR0sH4atw1rCWfmZ9Zg+6JzdU
ClWvg2Phv3X7MUojr6y+G2iyJtB34YJ0xvkncyVtgo23xbsfm4b3/j0T2Acj
wxSsy1tLmw0prEGcc9/xB0sln52TvcNODZKV8lLgwrTaleScrfVUEudpzlWT
E5x6YcvfJo3DkoI/4OroYvP2F+mM1C1/s4W37WGTTgtZGsvT9SSB6i3FpECi
+ZWsLYs/2v6ZU8TEzKcPRlYRm5cBFwpQRSW5CnUw40biG5ayGgAep4JMVpMm
lSb/fte3WoCFnxQOJFvntP2L40Hf+Hpk6jqd//gd0qezCqKfrxCR/ofHEbAJ
91VBs6qGUe6KO8czsjX+nQu0aW4I19Q0aZMn2SycbCRWD3begIuhfDmGovnN
y82YwJnLjAXTt+aGigKn/mqA1sUoMEFz83Nhp957XyR7snEcNU4yORYXCuFL
Xn0dEmukKtCOGi4LW48NFRPb8lV4Pu7JLxYADNjSmUCoEc3JZICXYvvKLGhB
Rm0HEwEJf2cucLlinB7caIVMGJIAV4WF3rq0BY4bVVskulxXvFg5121eyvF/
yAlAonbjmYhW0UTEyUFv2H8T9kaQOyzqSd67JXyv74Ww0sGSlBJ7VlY1lJ7p
xd/SocZ4Xlp1/R0l5VZAkzBw/5KlXUPTPZW0S/PDaW4dYz33dNr4qoBPrKaq
MF+BSP8fr3SgDgwwSEXPKpIBlPW0vGXwnNNgFOLqnEi7tOTOx7lH4wMH1DJm
Fc6+hHJTXj9lwxZ4hLFSzQQrMXqFIHXQhOnpr6MxBG67hipc46+QNZwbrtE5
2/majP+5kyR+9B/uc4WlD3e/XoBx7n1H2K6Z06v3/Z4W7Tfliopqu1zg2S6m
tVYC1t6Cs0Q3/bR9NP6GFf0PUbmN3CxSjR+NA8bF20P3jHjXjmuZ6+Wgu39y
dQdc39VxgPKswlAgUj1xw7UPDyEXlKvhi+RrE/07gyGT9flDVEKDYsbAXzYo
autDR0K1hyCCSB54fL7jWPteD7re2DE2sEKofWfhG49q+6w6ycTy6AKGkqV/
Dwg8+HhQvgliVpl/jZCHaANUdCUzThhuoDqmiClDwdnZmjId1WoSlKkrlFez
JKDr0i6H88f6aHxq+Et3pPH6tX/vOlV23BwTn0BK1Lg4oujUyzETyNyjCtuZ
9zwtRLVkFHnLHjZNPQlsylSa6Pth03Jg88tM6wIBbzuODz0G/RlTh+ViXChJ
p2Pn9SxOM8ANsyde7b1fKvOtpYW5YFltP4C4zGJG2dcR9jtCVMxa8BhlOqvl
ez60Oq+PDRvm42YcMce1jjCmPbtpbbg9PNUZ1i4mKTxeDZ4NYjXrSqnAxDOw
cNG4sau5jUDASdOsFbAhhX6V6dXVNTU/SD48B6x9i0ilDvK5wF/EZ5kV5j0G
Oe3xkMmGYqAllJ+qL3SI+FZEiFXXQB1vLvcsMftyXJ6HcZuPhJp+dyQxHQD0
WiaFOiM/41fkzhe3OAnmoXE7go2g2432cUti9S3AqJQdhBHmdsD5fsp3TMMk
duH5nGMREXSv0eOHNyyXH7MeWI4f+sp4GSA1C6w8ROWZD3daEG2Z7IxCDgys
esBeSTdUB397d/NJrx8dIGuiaxuzSyC45dMeqNd+9Zxn8W6bby/BO4g+ZYEH
Mv+t7nPObK7zvRVxW564Yp16ndel3lq6aI6WUHkCv3jXfXhqfirX0WkdaD1G
t0+m+fg35238XaGpuUbjOZToS04fHKP71nBKiC6uBkdOBx74eqQN5lndY808
C9tL+Ns5OYeNUXilnkgHXaqFbQPCcI84XOvwK16Dr0vxwWfu2sgsBSb9XC8X
il0UnrN2pBzmg7p6J/9ZnIDotSnJqkuR0VcH9yNMO9dc/S3SNfA6rvsUcsLt
KCm3VrL6L5ZjlFrsdk48PsVXbFKbV71HyXIXKyF9r7uhevt4HXxQ5ulTKIBd
yJamyH9jYcTpQXzND9U7bx+q7Ygbf9AU93n4JY0eCangz1/Zzl8wkL9v9wCW
qkjY1+Y0dQm/G8TfnzPWMjXV4GaBVVt7soOmxVoKCECyzVdTZ19GTjJT5ljG
AZ2RbR1qLLDjvCGfhsOOkxOWQiseH8X4iKsO5i1LaFh8eogGlMhM3vA/njsm
o7wue/3F8IErDiMBD230RMsUfSr9xcNW+t7XhMjfHFDfja6bp6DVV72hMS0b
4sKEXNyr0z2XLCrgKo7ng/7Ppbg2zK8enNRceZrRa44Qj6+uH3VFMWlbY3ZE
rEgX7DM8ZEns625HVA9YUBbagVdn+70RO4Q2R1QWY6TJsqAftuyXoL79xGIh
8gm9jB+0rA69Z54MK+9SGMfvXA/0c81HqBJG8l8Kx8F1cXeVyfMjcRcPTChr
LAc4ZmWy+9hs4rn3pXomuaPZVkv5KUp4TPD8LEsVtGclooo1Db/ZOrajioaR
rkABL1PjMtlLvGpQCU7P+LnHBTFN0NKaGusHKGb3EE9FTO6LjaV8fcJ48wjo
yt8wCp6vA21fjLig8NmSlLWMrDMGBf7Q5JUUMg0AdjgP1eJEc2CfPaghXxyK
0vrWAYl7aGWYzighY+TETGdemRO8OrCbTKItMrAt7tvSNe63pmKB1V2jdXjq
UjWpCRV/PDVOX5nBkeBIwfnx/EWp/XyBrGlO9WIUBXIgQY/fV1tlLVWnoF/6
keteOLibdyVf2VzDLDnjwB4lZAuDzrpjRYF08QV8wuvBWSk4wUcDmRYJzH6L
p/xUI6Dq1D8qBvS80e7qVhrY0X8CwYDqxVlHtUUxyq9N2xaSxuzDknYL9FQq
84NHjJmOgdXyRr2DEjM50rGp+/sEaZZmX4vEANyACf/xkZVbjzr0x1behYNc
O5j4YoK5eKsm4B26TYrCf5mQi5R/KL6n+rMjVesWaU8ef48TBRNUwiu2kY1M
8IeNgKug42DuxSOdE06KpKzQntaoAQswNXrwXdEVtU+b8D2VSLGza1Jw/C0p
W8/lxR96GcBM+W7/rjWqEx7tGeqh389u4RgmBrLTF6+/3bfSQR1XStDWKwqP
UcLZT0re40uBsRbu2kVRE/7Y4GZXNoqs7f/2p7uWDD8ym0ILsI/NGKZ6ozyD
IDkzdz2PRHCXhwA8ecdBQQQ4jYsz6NXGwW4IWqAxspxqn9vIKEPiFKr7k/to
CGQnUlx+FkIeSFS43XFvdRzEb1gB81JNCPabVL43i3U0DGIfizno5aBh1FsF
yUUazmCcLHtUZIJOyWSmVPmIJ826xz7YGJMBaHgE21uLjxSVc7MHY7beykFp
K3QYiwXZFkTlQEuLdY4K9iQoe0ZTy6T6q1/YAgXbifDXZ0JjHqCrOStfYVrN
bj9X4td2QxnMBp9WUKYsKnXM9fBAlZemUYEa6pqPnN49qyIo8hJnXOKjispK
HadeFzqOCzPuC9nrjk0Bn6doTomsXMu0Mgp0f0Ti9mDK2GafKbucU1etCCbi
H0TisQbSaiWzfD3F2CgN42e/wWHLKEbPzsjFEBb+4OjfZ55QwPl91L8VheBl
TKfBYlkkjadtfTwiQUflgZTG30Ze5j3Ss286txlxZ+383nXLpI1gFF14tEih
37X9M5j/PGHzrxb8lh3doc4s+UwNE+Y/XXNN/8WMo3rgzPLHE+C85jCyqUWV
KUEsUZz18Gsb9v5dSO616GcbxdImEzLmAVBC89X8lqOwSi4Qm7zubvsXNZsi
dvvWp7ktkr/8KQ0Fk3fW4lg6DX0tnuKs+mb1LA9VUMHSUXDemfOmWKWGIkr4
GaK7qbP/jeXcoyDMeDYPaiXkiUAywQmWjZltHQZWPv2syM0msdj8GBXBhcac
M+ReJrZF1o3zJn6+0PdeWaGo8FGJ56sPYPxWBxk6ouDYbD5sRVK626pJwm3/
gK4WsDNvBqrxEsa+SCRB1zdZWtAJQ1EIZdhW6FnCJ6lWaYuiNxQ6qUY5J88W
ZeA0W9ibUx0dq6A03v8JwGR8AlVHrXQdmF3gGKuDPc/iSAf4ja0xcIxuooHB
23jUvj+UMiedTz9UBgQ1xgJuyQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mnvsK2EezCxvIql5TE8xXpjdAG5hofRiNay5KjXZeTOBx8FpZPY/P4aAqFvDKr5OgNSg/t7f/s6Qm+rt4t4iMMzPEGqxGNT3cpAXe/YpWxEeF8FCun8pOVkLP5J6pleB0ftelH+nV6mCRh9j+HrSkSItFuVIgIfU4beDub8vs5m2fyzfTznXkDzD/pL1wPaEah77ZmEme1r9awG48FG4p7VZSHfqHBsQGM7GwOzg4s8RJb9rpJF60Eu8aZePYxFvLPMb7dXVVXyfdNEXLjpnmfFmemQQMuVJEdX6qjzyhi5IUT3/pxnn48IlDePO2QVOM+5iaqFBIig/Hwp9vELEJY3ltp0EfUHCxzq+5PkjPQNFdwug924ZFz/5FIwE8XOrPZi6/RAw8z6YAIXcdI2vdkspMon9Cg2asK4JXaDaomcDEJIdjuy3elBGDiQmsc8Sw7BfjmEoZw4ql1kQXIpK4xLCavPmACzTRObA7k5AhIklBG6JFXk9c+ZJ+6whlvp8J4YsdxFpDcDyZw+zgl3ZisgSEVe8ZaHSYJibJK7oRQbtFEF+k9yWPB1muNSI99kaltrwscZV433/KmLUQjIKPzdi8kf5665etGm8zGtb3P2QZiJ57Dt1iqTJ687ExP7rLSm9E3Zdy2s1v3xXGZzMg3JNrSaEDk2SrXIMgECIloqaQUJ25eWUN/k2JDz26BmqcNhClnDIiikkON/NA0jB75z2xjJEPaX/giYZ+tkNM2NYiP5QeclR4S9WRG2JskMhNPG2zufzjYbcHrTm91MltN"
`endif