//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ps9TldPun/Y5o++H5+AanFzyVlRYZRXwyMM5+hmastUFAf5BY3l++C15weM0
tGX3DUgKcHHXesE3jPx4zKQoC4o5fq2yypPq8pK3amNGwDFStGTYfZ9oE6Dy
bLUGIBvgVBivm760M/u2ttCpvi4B3cJOiW172dSxr6C7orbJI9otNT48jLXv
jvl71UMTgVbn2QONGhraonoP0Dx7UbjCuvmW4/46+Z7JDgRUb9cSg0mp6AY1
+dv6nd0gmOI0Pol2bchTeAKCVDHNsqkyDt3qsJKBgE80abWAU3H9bDFG3sFo
vQG8j15nQgecEojofJwbOhuHuOhOo6S0rYgNVSxCvw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f8WfpoKVc4AuqwDdk5iw/bEjS3MennaVPj6iWq2aJZRBOSjIG256U61yrHtQ
QRfmVkyPKPzU4pmTvklKFh/TSO1VLW8vp2EBIpGZbg1844wS+uFS0W9LkYdk
T69Bt+zAnMgV7rLk6iJfkX+cK4CgYS+v8shAB2KUXRPVnfdT1bf2Po/quBsW
LlrRkEfxG1AMgpS5ZHB35B30yb6gBZWG/BPhC1wvBZmioM+ncxUZZgrqjyEl
3K356SlfGRTFma8j8ONNAqNYWib0YEM96pksBNVjySy/nVT76Z7dD5N6HcEz
yo7BAOiE2qCYeLFimaxk7GS8n7DTh454LgZDNh77VQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
KyxFzGVndAlPe02SKtMbSfaiLG5Y1ZhjnDelwSvY8x0LeU/9fqtw/rTmqDe0
bxhH3XIGE7raDVM8eIurtaQ8X2LIBoxX8GbUp2S7pIFcOXqAe8NqBeas6a8D
Kv39qt2C5Wd8EKlck1CgkwQZnE+0BQBv8XrxMpzVbPrwH4N+2nV/oUSN5beg
c7f04nyUL2EOMuYt0pFt5kN6zGqoATFuqKPvHcMLSstn4sByz4ZxpfrzO6YE
S03F22U+FcmjySTXQQrHO1u0Zhrtmr8q8XSn5nGxOiTpZehVP37I2qDMN2W3
yxkPsjBrWW49uVLk2aJGq0o8FR/eqnYXRJ9cF8ok2g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mPwKKsZhfJaB5zHA2wRWAgJ4OaqXadSJA6/rersJGrmaPvAJBnrbeWycNI8u
8Om0SuZKMCVrUQTesuc8GZ5v2NpYYh/FPtHFFEYEvWMRyi1jJ3gtQpEI6E/y
uHK6AFHkNvI1i3mx008E91XCayOSbmT8dcDYPKsWiR5ojc/qVHE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Cm1tV+bZgEOyexm3BkT6D5jp1HTSDE72Fnx2R09SeNhXlyT5M5NvaFIpAZ+S
UwYmL3S1YeiGFDw9Ydko84miEWDSm3wxXee0Urgcw31pMFY+PkiUkbyhOGrL
cedG77QeSAKmj2VIIb2A2i2IkpEX6bDmeaAueKnaZPCDDAPoMU0SwyjxRDIm
F2BpCMbahCWLQ6ZIzH9gXu1jMW4tBA6Qd0eihirsk8b+bI4GNs0vVcG0DytW
sdy+ey0rrO8mimQ0GartifeKZesYmyN3HOUjOVk57mUyFtU1POX5um2riHhX
Ct3/OJUc41JVJ7RBE9CxRvSFEn3g6WcMceA2F2X8C+I+tbeWuRIgKHm7yNFV
AEoC3/EpVlLyOa+4BY2Amsd0XamlnhuQVH1WyXWSupkjXGWQnVpz/fROp+aZ
LvlOzZ2USgpC4AwfR14zLYNAuWt6twcGr83Hneuiuzu2jprnLk6+gaCkOnvm
O8cPYYTDRuty8lMM185xz1tX4CsC2Ch1


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NKeMxt7XWYug/LlfYG0XpgXVVe+WNorHoG84xK+Ko2+p6hEnqNrWFkuAb5Mt
GVvTsoMXJQqdATmRyRIvyVyGxIbwY7MYfUUHL1jxmGmLoK3VS2PlMDmaHM2l
mrxfS5DKCXIUw+Mh1Rdnfw0J1dYG5FbcxFMqrg8R2dbjFoLDUh4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fhx/dgmO902fVMfpP4bvzVulHT2+GFDIjMYbHLTGUHXg7PZ4gLykt9SR4Mfj
Le7SrpQyMAAA3nRRlXE9wHGRRMa8/PT9ABrIAWoMqBBayPTBKEjh1ejhb79f
XyrmtcJzSjrYfQrNLdVYjhljupYWHMEfl5d6lsQTAu4jSNQXJ5k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4608)
`pragma protect data_block
7ofFylx3dUhYI0o/U/kh0VJ+tzx7rgqoudWZQUs5b90K78Up35z2fdSEwc3P
Q/tS3IXq6s/y25ixD7PybcrSTOTr3NjITS5l+IoiEucp5DubYi6NJSd1/MR8
vl1jaM7sDhNgz5ARcIOf7sYg08W5zVvTltrACk90cuTeCyMNiQ75ql7JkqWi
US+9vwfUEnvolDSxipZq9BmIKdem0XwpUwp7wdYopZSel3LAX0Hwgsv3E+IE
tPkdSnTOLaGNju4lvdVbLGGABuL2QCZtAw/OTYXyeF9wQb+f4nG09lH907mc
LyHR9nLQfanbDDPxcoU4/8RUvAIcwLkNox5wCnHWR1FJY5zzPx2kEjMD3uce
88DizN2HkrhSdLiuAj1XhSHhFo4N5GFWEcwpfpW9RO/WPpb8N9uuFIL2o7/U
yW+52Sj6gkuX6Gay7TH5wXsf/LV6p+bouSy1zEQ/RpjIZUgC+GGM2eKWrP2f
XyJujiCYp7sYtXa088d2/gclMMQcXcqtRZyY7Om0MsEHxBKtMdsymLTWO6S6
dG6CegFMS+hUpt3yK7sedGX4acbPjQ9UJdOPVdtkOQTu0nKIPHjbfbk2Nvun
RUWodrwnxpA4vTtnxkIrgOFC7Yva1V4hoRzxTb7ZpaNA6YcfJpoUSEU6HaEh
GBkUuvb9mis2ah0ONFZ44pbMvPvdsk1QN3zTUH0OfbMoOVcaTbIQxO5c1I5m
d0ltN8OVKBLRM1RiNvt/cdNSTqEauCTj6QEqR15UuErMNGIlaS8wjBFv5SPD
veAFO+kA0h1Yb9kJdXYGx20kX3Cj0f4tYG+MJolL/efoR8m/rTidUT0rY2Wg
kQbQhVVUHZWQ0GcOiAuPnV3Eq0WpM9vW4wn+6KOdGwYW1kYzhluSYO0aWG1m
ywffJpMH5iq9umn7IVQ3HxJSKtHt4lO1cw6QXY6CHD+V5bgQqPwY+TTBgtGD
c1bMMRy7syE90XrWpCTC+3oIpfppUvN1q3rGD6fsG5uacBffStPENZBxF0tX
7MROMHYTIDTirlLqa2kIM9wB/VaX1qRXRoZRPnRaPXqerPosTFHqNecSkUF8
XsIUGkDQJb03uSlZQ+QYdhOPyGkwjwbqR9RcQzWPMZWVPVEx9d8Okx0MjYRM
GncI8MqkX3760xWwNtxdDAsn20Jttz70D3B6XXnLnH+ihY34KrXIkB9B4kdT
/EkKFdaRoKv8XoNyuZKSxcIyXcaM4x7DyaGwY/QacJpNSWpFfEZ3YzwndVCU
CjMFGygfFFYFVICp8LEswycoqgSMYRxiF8Zq+64FLQXNk4MRAe1xkyB3O5EW
lGSvXIl6lWK+li+6h87IESEb+lAj+9R1MK8yxE99xulrRbmjLJtfmnBoRKfH
MCeGronwRqyr8gXPSeopEOt0uWz9/PF4EDnUnQ3mkt4CKOz34F5r1PhYzzDD
q+lU2Nq68DfM4LwVczSOiHr9flqmUK6FdTnTRzRj6+vf2sHQnToZiwarvV+I
dYyp8ceWtywNzmZ69jfty8yM6o/k7Xt57cwQ7CkpRxKacz6JyD0pgnsTRP+7
NKaz/jXzqkUHpi0Y0lv/WhQO8WHh5DIpWizqB9tG8Usg05uPu8Kn0ARyo1QR
6iWVT1odcta4FnS/+aSgOgDdLuIbToUtioUzyDQfqjVibk/YHZbNhaayUzJU
kb//heD43RPXM9xRgO4UCvKG+msCZ6LzLm0a5qCwn8mqlSTqDp74HvKmWP4Y
0FUE5RH+b5uqmY44INImz3KDjnk6cE8ym0yLEBajlcWd0vvZe1CqXmBpCp/K
ghSZJ9sGO+0ipQ+ujk4mFiOztLL6BrhvaxjMgZlOCVoqOUQMYOUo9BO4zCb5
97bc57+uAuT7pCDDvTJhl9dINga56dnxhKbizxr1YEv/pnLsIG9Tz21q1xXf
4KbmbBJAS9XV+ohjEaBwreo3lM4c8psVQ9y/ZOvYSorBamg6G3BOO4kgpmO7
8gOd2zee41n5I4iMTYehVcl+889pxehMBdDUEtcNTtQcggwgxTrTHMy651D5
jDIVxo71OpLn5UhLuBLXKaXvxtad8WPft9vXaSIo4pDXxfyQ4GuS5sY8wZZZ
oWWDs3BYvAPOiZhOfHuh+XD1Wr7qKLRZmJQ9fEYih1IlvHq2pywYkRCWngnY
Ef+QLQgXVG3hEwiSzavtkEfH4mSPvryKvwFIZitSVMao1zt3/rk5tWIem6gi
RwWRg5pWU8GrlkgZuNahtDtoKOi0Paf+T/SW9YpGe/lLwA13bHHTthTYjpBQ
KXbRXkWSKH6YJGmDmDt2QkypNonvyMhXzDLY6si8vFtb+z6feyjEhmjp71TO
0N6cAaICgvfd0OEmVreHwQgYH9MLwVfqvx24nq7JtEDyczLzHgvxbemOU/KW
Tm0xYa2zR4GvfdG1z4CpVgfsRpLP0DddCubQTscKGvH1TETabHCzpJ5VowBi
wiZB6HOP4cX8jWg+V8qfd33U1x6AFhWPqBGgdY3emppcBoC086J2sC+IySIM
hz8ZUQ6mCJzWQbpvjxYmjZiPtY/1cqKtDJhkV7ODM/m1L/ENtxGCmNgKMe41
qI3UCsIDymfUZFy9yXtFSaTMZi1SFqcMDL7N2ejIbU2V8clmxWEq3Ejo/DC4
QNGbcB64QYvf4RFNbwJrnSJNnTQ05QVMkoJ6omyILRDv0Xfc1v9K2MLwllp/
RdNCWt9mseIr61zXaUM7KWbsHZvYrgQkzSyq9TlXzPmdcWLIOk/5Bn3D9ePp
tbdCkf/UVJlBerbLAJFxVWo/oV/ZPIBH/zT19nOgBTICWUcP6mKMEc5mbqvx
fh+qn7rresb9ma6J3IdwYqMnwWyWCbXesoWRt0Nm7/FmEZxQOxCPd6oRMd6Z
sSNIWaRsstUDRD0Jh4pUO09VQt6D3ZhlDIe4smtEysBNGu0vDjLglxre4+Vk
QRr/69dvkp/RY2jBOTfnPW+wxXTtxsa93+KWM2eH+gwDiU61edy5NgnT1WNd
gtSUQlUwGgB79QakVFR0PZZd7q9WH+JyyWlrdj/Aas1Ds7KgZ8itajdP+tPd
gsCrJnGzb8++Qc2QIWFkCo0zb/EPt+rRjlbufcaNZ2dRo1ZVoCTSi6igmbnj
xxNXWXXMvm0hVzQ/3mkTZIzJ1NiXwXYDxelA5tj6yAh4eegdGfSSr+UV9BmG
1iy8jjUlSzWYeDD3ega971MawcBzfEnqJDE80DlzVhII6y83vzbbeZB0dGKh
v1r0mmPOB8awksxYZnSGZpTmaa/kOhIzXnJ/h30Bv+2U07J6V8JfatLgy0kl
6xRW/KqSLK1EWIFMwNy48UH0rBLgh0hP4hna4gQxa2DMecEmrzTQBHrMTHdp
dWGQMjPj35477LDVp1yXpvt4n3eY7ncmX2vJ3TlcZSOVhUK050GYjX9lDsl7
egWCBc3Bc4dz0OpvATkScxh5IlQuHmZYZZUpCyMfwkI89fSNY6fKFvZvhcD+
OlozEoGmzBcp5fqYrC5clv6Cvso6t0WOH0p2xm6rmR5EWBRy5uojvgSnzzhX
255nerE/fjMGlTned88sYXRu19IE5oGITpW6c4mTUx6kDeiFoCr9IyYnC1oi
Z44fZnvZBk5gd7pNkRNXQTe3RQsk5PS4+z/LwqdmiIIT0iaPX2eYrKbtiRuJ
Rs1uoHFcwaDNYPl5BJgEBtiKJRNCK6OhHg3vMcmo63fO+cWI+FzH1wXibyoR
ZWK0B2h+J+/6uw5oZ34UGVhfAWe2S1F3Re9ov9QwNefc/o36pcSKeSLcbSXi
pOlp01mPoEwVeJcnnapmAJOxe0g6GMuNZo1GCeHNEBkc7xh77+aw73F9cKFL
e1DUIbwcnoKgJqAqB1pPSVcOvndhAI25q4zEe2bV36lX5POtDOCflKiVXgE2
JBskPBz4QnlXQSG6FTXXIyBaAabG01drfRwFPPD08cA4ppJuL2P0X/a/jMsF
KaCOQXa8oGU4DC8G/EnQoMTVYcA+zg50W8QuHbyCh91xBQ0/voyORl5Vv97A
S66K4YQ8brnQUg0/UY92bVBoAbqTMRje+uK4rJacei3r0uMvZRml6FL9UnxE
R5OJ5G3Mx2Ql4wpdtKM5y8EZ/2hm4Uio95ibOhaZj6bAa0kVEl7i93UOGPhz
KkPKA7aPPglEVr2Xcm7ZkzDrTnxCfujmGC/OwA0qqNdE7Iaq0I0kehbmZl8r
DAiicDNRwEWDSxyV3LMtg4NdksfJ7+wJ+vYzFvZdXqtPcPsF+aJtDl8MUXDf
lvFt4EMA+nejaAuKOcavqD/MGtBBq1/B6dkzLOtWYlRXsltqEdFwZum7J+0g
hEMRsCK5R6DgrBwc4vaM35G9JvG4YUPntyU9h6LNBl3FNiVw4Es/r4lovOiN
h0IHfhGF5JxcKN6QuG0t5ZMH5U49i9+U9zh+nEDU17ZFqniZAuENUGuYFLQd
kceH/7tixmRnOYZkyIGfqTivlmP8Q8MbC18zDgEb7K1Mk0TINxjIkVVa2B4y
PaUAjC6OOQ2FeSKxmA2ULfCv77uvQ8h0zMQh48m+/BNzmhdbWFZbExHUQ9bz
SuugBtbqbVBv91rh8mjXE75g/+rbDryhoKxwlNgLifC5B5z6dSY8foxEnof3
aDXK9tBiTZjNTCjgWcJu6JSdbuIcVQeSlJj1gDQmC5aMuhCCXAy2JnQ0Gye8
rgnlNusNktDpLaRrpMwUOGsrfuffa9BpdYcWlEhKkmoJ6ZhLpi7pqsX60Duq
meoO070NM4tiDx2I+1JcYLJjUBhOqGoNufPd2u0WtpsK29cipU0OlduqDBLL
DBsXbBYauh2y3IGB2p6fvVyepkvDeemL05N2k75V1W9v/yPAyYjlSDGRhNZb
A2MaylKqcKivTAr340KbE2128Hkcm0z2RIqpPOIxROP24U6BhiSS4lfiphAB
deal+HXQCJ/IgpzVBppIXtPQYwNl4BixaBZUKJQWqKXAg2BpJ2r39WAxgy86
vS+dNprDcEgkrgQehLrUTzT+9/IzrgZeQ/GIy2XpWCeVb8KK0Az9lQXHDxpX
IeFM2jPaYtY+AJhQS+4D+8lX40xKbnXhTuI6CL6ANzSDUg9tM67jqbN+EzCQ
mKZBeF6sSwm+NdHUubP9WHPQyYjoU3dqSBYZb6N2j1Fvb7x3tucfN4kfFrsD
9+F4kbKD6VaV9W0llxRGDNZ4jYKYUMimMvs1x5/d2z1dsYiwy67ifo1aJf9E
wUW5cqJx064SYH8eIx4iDPLsCvGEaJrQJof2C1qN7LKMxbtKveU4c48XmJWx
mJzSYdsy1PU3nfE6VCdWbmbbCxnzGzcC5iBYPZdn1sc6F1pNuEv0ZzCfqSDY
7SNgwKPi1YH9LQ2ITSrU89q88zqcxiC4eCf0ktLWO88SDKoFpifuI/RGxSa2
NGRZAJgfq/JpV3VUAaifM45j58sX7hatEGSJUYvS61MkMsvWrC2Am1QzKD48
1abNKa8wHl+inTkWymKffMqtWrydSmUU/gxt8kbe35kqGdzdMwDQKypvYJL0
OeyOIUFNmNHt3TCf2HI2qtuOZZAwiSZFDKDfiY5ASqd1BRvGIgB8DfqIjikF
xUIRs3sb20PKHAx2ePph/mUKF1/OR3R1K+p7kPuGgbdyNc7xM6CPoS6Z9n/B
czBOZwtmZlx0T49KdSgvkPluQYQ91ACmJlw9bGAqfpAlWkNhn450PCuNNaFG
8xcIFdlgLdSjbRkfT7/sd5QXX+9BFMD6RIInpOLMsKPbUw5HWcRYOi+22IiW
8WrZBae1Cbfr/Y3w4yd/RtBYLGybtqk4mYHaSnzoGUonWkLEWh0zSjQh3Zz1
dyysA8AZXAxfGim7guKTxIcD4pl28S7g0bQwCYRo7TGbxreqd0OtrblY5At8
l7CkKwmRQsBRCPJEyvPiNJIQZtRn9sqdr7IeSyslyd7j4CQB0RwM2Hb1JzOu
L+XMg9N9TVVINcTxvrqAg/MF1/y+/aRGenWna2KnOHHO8lK5C7gVEjJ8mfWW
ppeqqiYknfmxhqk610dI8h+c46zLNy3cYGaiQIqEsfRn19SxFv1jqAV6Ftn7
JBkReFAxZxCPUhXEViKOFjr1lg8uaqzNg/hfcMQZLaVU614VQrAXMun7XbMY
A1bHM0EW3Iwf+oQ+9K5U1rvg

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mzT8TNfU353DrNXWaGGCO3KULk52v6xuZ0NscBvQ0NcHYj5gel2QFMJm+Nqfw6GqDBUUAvl4wC8p4tWDageYU79wclpdVPzNnx6rgFeetXazulVZ4AYkF3+4ay2Sak3V0pD7X51idXod9uUnbaYNjnJoml2S4fFX1ThVNtQhRRdUhoY03gai00PosnJhRMaJLE6UyQ5YUk47pj7rpqknybJn+ilCmWdiE5tOWBQlC9DUBXCkMAOTVaExXN4Er/n0Sx+f1wiJP4s9/InLzBnT4gn0ZsmwW7aLwe+8jg/EP/wGDRhEQoMgYul+kAhF22/M1yYLBb2iEmTQ2Y0/rfKyM+uDvwJ7xJOPxmXoK3u2esMC0unxjpVYVuX2NBGu5OCod2tEyxO25HFZiZYHin0jFeEFO0D0IP9o2pKxUn0U2vYsat8LqOfv8zYyrSlnAictDqI0i1WTKaZ/pJ8hjf8Q079ovStAkuFsQH6QGKPhFr4KRIK5kfzZJ6eP5wTFQd7l78flM3CzOkk420NZbmE5Ixzh2bKfcvdOfWt8bqyRP2minJKieY7GfSXt2YDk4JfJdgBcSHc2NEm7KLKkro1lCSmhjidlBzLYsoGYRshAP8f+c8RBO1IYnj1GyVakcDEpcLN1CAIW8g88cttCZq2awry0xqqUaHkyY6WZ1oxX0imTBRlxA8egqiDHdb984425GxEP5eUUPpZDni6rtNkTdqrVAXGeOS6FWp1ySzR2r2CxwnfxTeHcmFs6B6zK229NQDluynmmORl2io6GG+p2b8"
`endif