//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mUYCdSVuR/yy+r2bfCdaUcbP7jkRDBi+UKPK+0YsGOa06mxb25GsIxrOuh35
K6ko5IjsG2XyUTCz8ux7DlHf59Fk4Rgi7yJkLeyTB4+GAXIwLYICjnTmOfuQ
Hke1VuxxoQ0LvAKkafV0QwdyPLKFl66ddscoLw79+biYaP8ma+dXo4ihRy3G
g8cYDD1bHBL8oDcFIEniPsKmkFH0Bgpaq7tFJkFuzwDrmfTWz/2S7QdgslSj
nrt1fWaFmPVbKFcPeUjlNYO3v4Vfw/u0JYN4XANtHlc0n9M2w4F7d3Hr8S82
uKLl9GgCAjeWaBDkF6iD2mG7hFIlqwpfPRVBZ6JOSA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
o/9wjeHwKimoSEb30qc+MDqQlD90Ah8WKdIKnaMrHqW7jSywBMAlhXs1WXsL
OIfOecIM7Ob9OaJAd0xZJTekFUmpmtbo9AmXFlKrjqQ3LuZNTHhKw81ftaOn
+OrF4w7YB5lc7oqHRFjkxCajwCrVP4egSr7OogCpMCiZqJAXJwkvSoofgdjw
9csj/1jzNuS9XyynnJhXdc0pviWcb3+XUyWkoYfGF9n/knhV5JyaTOBJY+y9
qjBugf1OTYVRSrU6JuNYN3Jvj+4BAUMoI6/J1QbWHBv7vzk/b2MdtQbGfzgA
9AwJMLpNIzTGpFyDDzTzYO/EMSw2zTG2gJMRlFmG/Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
X7BHmzIMAA7ekiVqieKWStF2rbvhn3s0w+mJNk56yuqWfQ16cUDT0Zum6kav
ongTXka88cfKeRePT700Ht4UhdHyxfp7RudpLYazZ+LW1f3WnTgvIR3QAPXO
9vzANRuqVMqSaXyfUln2eL+UBM9iSU32hgTG/1NO8T5EaH8WNq0srN5QywfK
Evm+/HAAjHEfODiMkt9IPlyKQl5Vz5SskuSIFi3FYANTd0/X8nHY2qjp9oeL
Z31/Vf6bKROLdOHz+r2V69nj8c/AegXdisyzBfs0li1PkypPsyoPVumCddCQ
RYz1wbeYBdU8G8/QRck2iAWkE4X+aA+KYLSbz4+L2g==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ELqTLjX0XdSyF0vtVvK9uZoBqv2nAlQVg8QeLCQopGpgatZIa//397Vhq6GN
IflRJTdSGYytxOUYUpfq/Pxb8av9hVyaFd4bCDVYTpr1hwXRWcvy3YqdrmxY
G8oA/DaZgz7bx7NS7NTr5yinj57Bsb/ZjrvPenJB5OVBLPcy5Fo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OSHIQJylN0a6Q8xBaoqPGMeBduY7Iw+xLSmpl7p5ijEypRU+IDkuHOWlY+PV
6bD7ry8TJTuOmxlIBGaf1BNUpnNyR90lKVv0dvMxhMMhKvzilwo3srSa+bpN
6KRKBaxO5EDTp+Bcq/sQ95mNRaL2HrhuvyUzZVrVSnerB2XzlPntDbKQiMGo
2/otaFaEyHOsJ+O3v+hw9ym4//QAFDe2Zu0oRbZk5xSzOeYEw2f8mVu08ayK
XSBNBYPocp3qB3a0ZyiUAoCx5aoUgFx79Z28WOBXpRiZHYTnL8PeedekwDJo
/dpHhF63Q5Rc/QjoLM29f64tCPIHO8d9TI9bZHxtZEDThzONSDvR36JBINmT
67je7mEbF/bs1k2eb17ZKs/efF3MytvM4NYNngCWQodDltVHqFNbDuuSkitQ
teQcbF2M9AG4OGsk/LUqs65CyUguQWD+P/Dw5xe96apkRQiZ36USoqy7zdZ5
LuP/xMgM3PIzsYk3rXI0a/5Yq4aSViA3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
P5CrBgcIs7FfEoIvhJoqrNcaTbb25Vh6zyhVoseY3EA90oy+KHrFXpFcs5nu
12Ak9AVec/e3NGVQbFhfttHuu+wyUQFuJqT2rT4hiK6wcgXD2Md4et0kJ3Cg
2051n6k6XQDzMjie+hrRbYL6/2JXtT3p7YdOHwWJ7xRxMchz208=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UOYtmitoxAa8wbQAjE6dFjB6T5kMLBA5xgL9jqcC8gaMtjNsnBZ0FChKKX/I
nFIv2K0JHN8Hky9+45wmXuheaR83pFDFvWZrG33b2CwI71R6PhN9DfY4fl4L
ku1h0vAo2RxcjhVif52kBKuO7LBmkVv0aW9siqOeBjcGWWbV97Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7312)
`pragma protect data_block
e1tsZ6GQyrW6+VDMULMGzrBBuZm1GR8Zp89EYyTTu0ml/rAPui7i65aopjrw
Rjksi+QW433jD+qBXRD4zusnC5lUtulaN3CWbm4YPGXQU8POKw7jJehq9L7g
1Lpf3xeRBLoSZqwxx2NmBePLcHHPgiAWJ2aqB70n9h6FgFEgszQdvTH1x4rx
mkzDpGZN5eNtFyf0fojcvOdDEVEkcucq1seTFyfrLULiesAw0fDJu3AkEJuX
NWI0rrWk6Ou3UtQrFI2GrU+A/DpCMayP41GbhmV1A3eI8P4FrRSr671i2lp0
VWdphol5NcFSOjwks4vR3uquaHkp5fZ3lnwiuGnGOaNb7dk8CGq8/HycZT2O
YjvtyP5JQ2dFyBB5o8o+ihiss89XOPC6j0A+U8fa3kPtlJnm/eYslZZMNYdY
X9D/fJnswP1tvQHVVpl1YPyP5IhAEDTYBGEC3jMfAx4D3SLHmaRxpkXF7TeR
2XO1va1GLAgsXC7CE1USq81aEfVyJ7aWhPqWjttgW3q7TFMRpbLIBzwfkR+/
+97+jc4FRTMI3MqYce3PC0WKBenor6O75uKotuR659QP/k9XPpu+Z92WLf3/
4YPwVXD3GpEH6cR76RsEDvQHD2JfjF4DIxLwVtw64d4hR+cqOPkpQmNMBUCv
VISTvBVMPS+GdHodwDpBPXdb70+chLvwRDiyhbBvfQZSAat1UO1hRpnHxcQj
JIVRd3JQByp3/3JnvqIhPUxD7hmK8EPqYKyAP2W3hRoxjPm1kBwYsz7CFIyH
KPuWrRLRH+KRe4/V8iWbUTvZqgz7FMT6TOabw4Bk2WQgtYA6gdVG/oKDcOUC
5Nlilzh/RzlAfSYnGOznBHiIfjwdvCAAeObkf+5i7h11jpsYJnKncxPOP8oY
SQX8NkCWr1QJ3Nb2eTvIWsmjzKSflvRN5QU8ZhC8cg9isAo2QYlpvixRvMvv
FRyySxnF/A3mb+Q6J9Bo7hqcATOK1D45DCk4WdzQc/F8rKPJihgrx/gIDJt4
w5IgIgob9hcJ3g57cunB89kwzrDGRmoOXm/4A5oyiVaPxxBob3MaftS7Y6qr
GnBgaZEG0uEoflv9EsyJFoWCXPKC6xU4AEPx7o58R44DN8GRDrmfkisr2pq5
U38oq1BVdq4vs+tsitBgvhMfE6GzQRxoeK/y+RI8uqY8ASM4FWu3RReLfVjJ
mcOe2pgp8MHsooR90l8EbSfRR3jVo8fS8BFflEj0IJhDcIJ/detgtn8VIcxb
Ap66VauacUXQxJzRuMU2mx7TmTrF3Bmr4wl3ReH/OVH7Xp4cyipero1AenMz
2v21sZxlzdQwPucdx6QtlpDKHkAc3mj2bf96seE6sbnZOuT9NmWy4YfOa/Kq
BunSklR+8+ndKFzHhkPhNqe9+vrsgTwOyothLuQwrDm2qKVJUAuMks7NGERL
6bQUFmMnIKzmPRZWWfULXVrapcPt4axZ3Su3+hdCmFco4t0qeNw91T1pDs+6
C1RLdTaDBX7N6n6IYKQ+mr6bwzz7IDhRgJD7j5FAacNBNnQqwEr27MptBtHw
8urb3LdRhAeW7NT7Kq9Uy6JG+K5FJTbeFUc+oIeTBXmxvasg5Ott0Eq54A0e
oKWIFGfNX9SnavupjnI03oH7g2jkR/mj8WInc2gcthE1p+3m1gAPSJPYVqsN
0pgsML7gYP2irME4OAwJitxEEDYZ8KPVkVllBiS1kkbDxEWYAXaBE4Vi7f9w
He1qyKkrRF7TSh87tSiUbBfuRoGDu+WYR7J2ZT3Vq0LPPvw/lPMN3Exn6gV4
XoauqZ08wH2rFp4anMi47rX/pGyVrvduXp8Tf6LmBhYH3Td7/sJJCBuphM1K
NTFrQaARvJlSQ5kon80g/nrRivagtncyEYKVb5v6KTN+7oRPh+ztVnwh3mxL
6iy0hRw5vm54VExFscNjlxonz4UVgC5vE9mwu+NZPiBeLShiDA5e1dorgpyJ
gCMf+zf1IvQS9HDe8QI8pE6slK2mCpugsI17sBvdPKccO6qhvHj6AAkpd1mj
cKjFeNlqdmgcmujStAUjWthZIYAGkUEV+jUlAstwQTJYqKG974n+EIxaxsRM
PYOjx4jeeodiKZLWBjW+YbwWw9y4O2HI2uQCBmRvnGTheKr+ohYVRR10su9P
yYUtSFqI0i9+FpDCZMq0ilNtbJAvv2iifDkdctv+WAdUa9eb2v3VpVoGsl2j
X+sjUIo2wi9O4r4d6RQ0kbZI/WvfW41bPUH2w41nKnyOnctvzyytPIXISCc0
Kf2HhvzL3iykXSyI+jkOeYxjv1RzTbE9LckfqBmM+vuC1kJL26/A5QtodOHI
oV+AIp5rkimhF4zMjk2oqUqtdEIuICKnRLfAhvsLyJoi+BCLp+kDedouSzCq
5OQp1eyj9GkhmSvlMjjjCwZ2orOOd/t3JcsKR0UTX+Z5JceMjCAV3tWdJFmV
nPdshQajw+O5QDiMZPdELYYex5t1SpGOXVd9k+hB0s5oi0dGfyJtiB6iCF6M
hqnKKT4NJDy0H3t9MJs8pG822S2bMY6//lQLOZUILMYjCh4lObNXHxf4rZBt
IaM6dZBDE7cBtT9/Mge+0EJe7T7JXM1eriCy3ckMfbZ2ikYpyBgpk7olNkxg
zGCShCGRfSVDBRWsu0b8U/LlVvPT28BwQrqVYP9YsZ3AYwgJIC7w5QJvgNf+
QWPmLaKmwC4Zf1mhJ/jD75LLBz+y9aO7xFA+pMhCfGukV10pBkXoTcRGFyKc
fwEflRl7u2pdHW+0/XguGyEvqGXj8K9aR812CTAcKwNCPAxDNZoYEt0a8+q0
cnK4GPu5f1i2jL+F/0SgCgu3klYEn2s92hC1qHzZv9XpoUHwgQVZksGA9R3J
DhKjLkdTPNZGwZGTSbvN469R+nnNBLE+kBjqLXITn9PUroOvnss5aipnYJlc
OemMJxrU/RzJKyHVF8yvKUAEwE3q+lfbCxsr3booRCUb/YvvacWbeMQoEAgd
lf+8wx+NTk05pQRGytGPXQWOzA91BRKtEeYt9fwsBgMb/a15GGyuDfFjHLbb
p8jg8WDYeYFZIM8O73fgbq3bpGjJIpGps8MpMRyWsLajiOsZZbMgCP4lV9il
ezjUCQpsSr64vt8PzzG/x1b0RRYxtiCNMEQaqKS96xQngtslW7KFQjsQ6lqg
TOsdjdr0/5oh+2MBKmrxaOoeWfL1GHbxjdDIC1vC8HfroTZdHfvEKfs77ORU
SLsxNUDIHCGZd3cjYekiFva8EOK8oi2s/+PTWMANw4JUqBzoSmWYLzxFHbIC
K3rHztPDQGYLm9WrHAICBDFbmVEoBsCL1/2MvDcegse2OxYMD0iIOGH98MMY
ODNHzYzL9PCOKOvC2Omb+9PrIdIu/6CM+FuRsNML7dd59RyY1AZuzyGUnMQJ
mMbKkK1I5W8Jxeynwi06RRFpbe7RHdMVmUic/r1ppgrkRD9iZ8eoNVmHYHnC
BJ8L1wcIcmnrwDaqmTAVaSCQxD9n9PxbgxpGcZacgc22YbYD5jWIZaRXOp0i
9KE0epsaQ0lgItjXL3tgSIF1/MvpcibXZOhIWvqyVvhynI+6uskzoaL+LXRO
AUIeejNOTRPnyJF2Bmedw4comXmbmOSb8Gi4jN+SCF1tlgjbgv4p88EKWgex
9YeTpK2PLs1YnIkZXke4tAZB0sWD8/oDNr08tDiEls9YHbIY01LJPH2240+Y
7iZI5xaATo1qMaRZ4YdYYKBuxZ8ai71ieydJXMY45JjrOgPGoXZCBlo2mf9M
pH48AcZgu6LTxXHjUvC6uSw3omWzrYQhvLCp40g0mwQQCKl4fSILESNmlErP
Wev5Tn0U3z4iDn+FP3WXChM1oiun7oT/YsGABETeFzLj8BYbGqMHv+nWE+sF
gXflGriJITZ5yM+HlFWdHAbwpJKDUHdyl2cAi/joNQWkYQImfezfadN0ThAa
rjjKAuQ95UGMFcauNyZPDHQeutfKMMgceVcL0DgTeA50zHEZzqFI6C/DCgFj
/5GrQTXn0JzuF4ZmB3GeZZAoP0Fk26VB7ZXX/M0eXL3l4yjiWHBZJ2socb1U
+FLLFFAew5yDm/j3vYr/Rs/XkbdJgIu7i1/Kiany7B6WHljsoqtwJsmH/NWU
Q2dktI4afEqEOAERi+5OiPzeV7e2EjiY4Gj2Ug804aQRUe2o985Ir5/6Leq2
Geh0keAsz2RMgRNo/SIW20dfYJmJmH4m5Wafhn7RTOc/dD2+aZNOr5v0AA1O
QNfjsH/JJyfIcpm2nfVJrMkfsiLxnDdEXdZx8uSZhffCysg4LSqiwiVg0bZJ
waviShoVWGA/EsO+hWzzaDRyVIJNw9JT8MWBUMVrL+9dfvy9lwmmhNQgz6at
/mhKqOLDEIoXIQ/56IR6rf8sBtCeLoz3tIGMKDtGwWlC0aGTosRbQ0BfiBK9
Lw5Uj5OiBPSF1r65pZ7Y1raI4wc5w2CxruPtFbSeU8LBXXvV8a+SBN9XKCDo
HaZ3coTNKSQ7FTihGoUXYSS1MKCXWJo4L6hmQWr5CLYX/64spo7NwKgZGxwQ
7tLIFenAKXjHrsklj+lgW/aKaf4kRgmPrhrnTx6KgrZuWi9naol6ldnKElSr
PZ7JQQCZdX7xp61Sk/9BfTvitqcdNPnDPR36rVK8rswP1NCW3ghsrXTPvCcf
Xew7TBBvCkX8kT/cHfs3mfKzJ+A4kFCoCiHKd0S01wjYOm1gHRBqR963MKY5
S1u9gx4njMVb8XUxSna8721ufUIB6VEu4FasuGB3DyMqIrXQPTg4rtw9gJET
fbAlhmkAf1mhWWNn32EuSIs3s0Zm+aXewFwVe4LlbT8NEovY5qlRjdLGJgtx
rYzY+98u2kFKGVUei6l7Ul2VYHyP1mGVBoX7aMUkTe0uBDUF3J1ui8RInDR/
u5k3tDifWnvWnR+4fdHp5AO/vLYrCEaPZtPaA2OXJZdqVhdylYCDGwPU4LAP
OVaPSG6LKPc2aktYQD1Fj58KNU/CfuedUDZJKvxLb3l7Ud/AEx5fUFE/0IVm
MlSClQeWjaHeyi+aamflEgK+y+6uQSF41TwBUsmSBM7MsODVaA1nGmdRirdh
darI5CHCoYDO++z/1w9kO/asBldEoJwFRIifywzpSvdMsUvttoIya4BJMGSI
SFCUg6pi/18FMpMnXd2SmOsSVYMoLZtlpk4BdBCn/kVMUJ3X/cqd/LBS84QA
lz5Ps68R6ddvVKbHZZeppiTRUWYkPnT6B5LmpIMdL+12ESeujcna+zb2CaV0
85/GBRG0TknULTeb6lNR5eSWURNFU8SspvxXg1my1+VUEkThZ25yG3bVCLle
dD+HocwPoyrFiixB04ssfTWolM4z/lYKgzLQVsc6R+YDdatZTiFMh6jh613O
anV3Y5nTLP5oqkk/yHLwoyaEup0NnQiBICfvjbVAtTpXEOej9i/Q5nXCKYZH
Mr9W3vNs271vxFH1USGWY3Xr0A7MZzQkomUEy7l0UcXP9AOtTzXEB884i5hg
Rfdi/jYvQwLgHjvRCRXJxjkJWByEgYB5lfdxlfx3F+qDbW83LqPO/NK7y7mu
C8NT1Nqizb6ySZBmSUIKC7lIPRZFsJOs3BzsrEwtlVdJwG4ethMnOU8X8s8+
LjkoMCWxZ6WIykTQXs7t+ZoXdrkVQ7VNujOjdITA0PaWCWXCFpaYcYSMIHuH
Rt9uLabu4CO0JERhUcgr1Ry9TFp17NyCp5GvY9b0lxXb2gwGr0fW31EmmdKR
e5HxSwtbU2VnqQGhIvybVl2igclFbuv194CWb7UZNbiWjqPb9kDkmoR5SoZW
F5s4i8KFq0nsxKOtjQdpY57X10p/TQWWOEz+lb4TphtA+8tJgPcNtCi/oShE
NkdCio7jcVkyhBT8rjbDIZQ2hQlVXpzJzWEunfEztCiBcHD1fjnLLJEonfUO
mhnOyMRwYL5edhhaDp/z9K230GeeRuVKYFDC1bEZy5lNVonFUPVFWaN0tvGG
QXfdyW5kVtX5o1NEYA0Db/T8hnnJlCvWLV32Oe+V5tg/+d/4hT3qvRkSRDD4
u7JhbPlr4k7TX1csWXiX+1vf6kiKwyDKStwIoT+RL0soRhT0WFsJwdJIrzgQ
pCAvsPOUVKO0NUGE7VMyDQeV3AwT5xWCe5oaCRdjem8chDaDgL7gXT2F+3sG
6HdQT+Z7j8j1ZiAQtpHq2qWDHwpVlHQHGhO0eknxSWDd16MadbxqQ7nZBNd0
L1UZOKY7DgOMQDwhljLI9FL+m0PICvvuVDWWI1+c40j42b1E4lktE23bq6d/
F2xOAveJrWH9H2iihriYb23WkpNJBeK7FkiEkVeJYKTx1RCv2jfplXm9PAHH
CyEUyOftWvvDV5aAWBDYM1uecxe+ZDywA5cevHLTvNeuVjkASJ3ZmyVlQ5x8
a6DRRmqSECJVxfu1dqjgbLboM1t5RFWZxscJTkN3FbOxDD06PeWm0OCQjFNn
eZ7/b/R0aVww54IaNQOXnfKld9nPDDJyreP4tz/YRAymDxrXj4E9OuGf/QWS
YE2NGphR6gZq6GH21J6IJnjD9BrLkwkvZlC3b7lmj2N0sfPHg0Jxok724qKZ
4FVLJElgEpnchapy9oFH8z9RNGSEi/f9/xwjN1Iw1EnQjyUheU1CKuNzfpTI
2X3RGldvBkHRWcbL6zqHrDAtlvNFD2ptuJAg4jJ164JVwoXDZsGtRlCcDnSX
g1/WAlYp4wJsz1KXiRRTI3VjiQPeWAJdFpNjAyS3eQBdUKZtb9eyHlTs0L0k
V3oLZY/IB56ygm4gVc0hW7b4mfLSPS276hdXxAc43/DfECYg4GPpNmlNvwyS
gFMgWGdj/CZ/ZafpV7QT+x9Jv2OCBD0N3CIewAuMJiGDyGxMH0Rs5i4kkQfd
spt/VV0GRj9qdLQEhNUG6ozIVt1q1/Htmw42ewmHVo6hA6ffRP/Jk4AzcXIR
EfrfXRO5i7ZKhc5H6VurBJz2LK93SORhe5CgCPRRHUlnO84E7DS0BSBEaCcl
qzTBpVR3LBN9+7/QC3NVv7jqepR70BWCI4bOm8EUELey1cbiL6tFxTI7m/8F
RTkKGiga4LiLnPhP6nGllfvoWzN8uuYiYjJu8eZIA0v4Ef/B+bTg3g/fEjZS
mEfdzx40yyaIKuMdUcRXNe79B6xE0D/6DYngDy6SFpE1+gMlCfgt9y/msQ8a
ys1bEN85XJVc8fFJO+zf+jAa0luvQm2SIUxx2KhTygeI1JrJD4L55/tqP3zO
V3sI/YWqLoJvoNzEdF/WG7K4oG+maZuyxmmQne96httjvsl+52iwNbTGDsqD
3PJiwUwHpJEbpP4bqlNMvzlXQy3nIxO7rJYCuJRU0g7+D4QelyL5PDKJoa8K
YNCjZS2MhmEPQWn4nFJ4Jhn6/6PN19JKarZHWCzWKkUk935z4w3NxpUgCQsa
cxEUW4fS7l3v4A0vo3lkj5o6/QO7wRuZBFwg31BdccgZPo+i08oiDvd3l8U7
/8ASraI7wwe6324DGuV66k3L1Me1sXp7n8Dch6vyqnjy+1BZGjXeoYTecJEq
fDbIWGU4jNA6l9Bd6BH/pqJKPRNgnUideiaWaWpw8hyKhcfQBhoui8hHHkOj
sSucxbgkTNQR36sNHlIWCVkK3IksOWtxJH717B/EvYzAsdYQ17ivW9fmZN2b
LVWVhn3SZg+13W+ruRlMchFgL4fDmgzTvm/7pb1BL+Jxpg43jmtz/igg5PjK
2uliMFDyceMNwRfL4U2oqa3ArVY6CvkdLTnDHRTtD9N4bBz56g1wmi3GZZ+0
SCqV1PIif6d49N81fQYaIqmmrpFgSPIlwSsO8W3eYdIc/4G7CyDiTTpC4oh9
avJOzhdvtIR8o7p+uTBt0ZLZHi4hxoDFSIOoY8d7CUWCJuKxpWfs+I7D9BeT
9z5lswYapSDnzsmRCQXP+HfJ7Wjudiv3gGpp+WpKRKGvp+jtNN/wI2iAj9mt
9CQ7UVX0Ou0CmU+bjB8BgCo1wuCmWrDhrc2Cm5wuGZ9MBY20tYPMiKK/jlUN
5n1dHLz2dpZAr3JfpF9tOecU2RqfE6zXGlp2PeuWs/7g+sE+gMcVrsLQFexK
dlqQJ2BSkO0T8fdgBduHpc6d9D/QVyG5YaU7KlkUSCxG3cgKu4QbpyuEbCWx
OEJtjT2/OmRCWQakypjdp2unFDYFttcrb+TaRH1yvdSn6KIkPmxGx8OB1jZp
WHlqKQ2Vtce58gUFdyLpuNdDnNFlEVZ7MykdFSfYCsmTpvIcy42VMXFXTeCd
ARGyPIxVfP3W0vQ3DIqt1xUot8O1MrVZpoTe6iZiqK//O1dfUWwBNnipgiR6
qyvihI6pXWnsItPJPBZqnZEHRC+Gu2n5w2e9UsKz8tFJzMCGSRsOsSnPW9HY
jXGi7Jh6jjaNPRcGyAFZljgq/ZscIgq52f4h0QdusGCBIhIY+3pVUMscYCsS
GUmzO/40G394HX/G2w8wA1CFwsJNA353H3YB53mck10WqFfJ8R39ETh4tlQ4
EZpxrQSSl+Pj5HYpyOIYnTCscS9wy6UjP9OTPmaWcZ3O0WRVDzP431QsWpXk
yj5Tbp7oCedG1uruV7QUOfU7JkmeNDuXhE87bC8cuBlSwn9LKaNmTPmnZDzb
eBbF7jLmX/DnTOFP4eiot+LNZpmiOe9+qkpJHvivSatuJbJLAP49xH+9REYk
ym99FaN66/zyrIY5hikRaCYoyv+hA4dqOvFxOsP+oT9cddGsY8MPwFkC+d3X
Va5R8kYd0RQsN3txDMxWM6ckLRWEZdo8EVrQrOuM/q9aF1Oru7MgggarLedb
UtO4JBVVCBq1j3g9c0WQ1qWMl/AeZ+3bxh3Y1RTiHjK35lwX/vuEujbBFYPt
W3PSD+e0vqmb7NhYX2uhAohHib06Cfs0gajZTN7zUqLmJw+vO72KaHnvknFF
ybcDk77wPaqGuGovGw89eUmCMHr0izJyQtW8XEQqEb2O71vmSPMpXi+j8zBk
p8oYe9rosrBZ6rrd/XHyBdAJere/IWVBMA1l62rlzGwrhi1SI1QHoGBgyKEF
PWtfO1SIXlZ70vBHABYXFoje8VFWjTXSFZilZAwPFCS0b+knHx5KEOXcIK2A
kHe3XHw1yMlWDI7BqAqLk2VuTnLcA5djbttlUoYBMHyL9FUjIpm7RbGZytRE
bMgPldjjnH7hQGjrkq1kEnDvW0uStQ1idA7NeMSPgvmMcUGHlUsOlcUvMI9C
OFJAKg2+fxUUW5SZtGEddZcUsEkRI/CswsYF2Ekq+Lr5lsFFzDvflrESuQiL
4hLFJCxrZtu3IayBVoYmJvYfxUdlRmAc5EyRq/wL5oxdCuXlC+MgWdBI0JZS
lnUsDyVjN6qgpyqoHDflOdMn0ZofVONEFcDD6RMFlecdYGSOvI1DUOeFdd+E
jHDGgMy6FUIMiK2b1NCr2zFydIJkpEQI+TEUSb3hoBaijlANFjzzxWhNwB2y
brBn/VJYskib0GxHXe+hlFhPsDY0b17YBWHO4OlxVqQ56cWHPGOeNp06BUKa
HWmXeKMo+HFCjxUkNEuMj0heqXaRQCaXAGovoN+YbE0xxDlle7l5jcXyV7yR
kzQKz7UrINl68Aquefc4BAKj9SvomfY6lCGapU/DP/clct2B8s5GXGpO0Evx
HDQshSJkCI7uFnIsrdwsg94oUrerTBKmjDKwmfUbCKjzhymq0P1RBPNKX6/1
zejP6I1r2t3+9c7lYD0gpGxLeMK3EQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "gqdj+Bhjqx1HIOvoRxnndmXZrw8O9IOJiBLHVL9y+7sADYqabq9i6IcqVqNsa3CsQ0qSvYbfOz3APXiqixHGu7F3PgZxyjQknIVBXaeoMGiZ1HLO9UaTqGJxU2WzoxHLvZ95I5TvNXGX/l8fuH3ngQIev6fsulB3eaVDwyMKby/JQ1XzpW/++wuu8//SJfOA0pFsYNjEqfw/KQAeoqM4XvAn4+PdlvtnN/wQuueTZPk6KP9og4iaWDuDtbfnqEvgaTbnVXR8FNseiIB0eT1ehoj9sSF6z3RKLb/fuYF0cvR7Ir80eNey3SCka1WXRyblpns57nCehL8DoRub93uN8Sloemqv4EFsOGzqpTIl7UOBsG83EAjA2wmS5O2aoepa8rWzslJKX5JltRvjR+KCsI1l8cHTrbOuYkowhtQ83GE4Mv3rpX/YKOYYaxFjYvP0rHFmCJEWveWSZG4DDI6XtQUeDXAKY3MXbx7xLTbtJgK7b9ZkjXtTLhQMIZlYCCFyP+Zb556+idbUqeecNwrWZ2If28dHNJFdo8sg92LLigb33ubgh5mOIB/D0JcHMKjNR5MTOerB+rMcnqYRcMsM+RJmIsnbSqISIJf5MyoCB9C3/ocpy9Ffxdvin5KBS/FwqKAzVuuVLWRwxHqgs3XMBzcHm0LbT+xHixkKs8ji6NqucKtdoAcghKSRfYK026zHP1nQs2Q6814e84LD8HlvZvZLkCAEpXRa5ojZpiWzBXLN+lvmiXMBc65EjLa/npPliwM9BS9CZYQFlfjx3IvFfpi3qTHPtFRds7CsPlD0L4McLxV5YjpPOJlquM7IHTyZXwRJmrVIb0OXnpL7QXyAW+uiPaPqCPu/Hm/KtOAq9I51lf3BGuOmwZBAqt+SD3UTzIZiP7aT3dOc74tVaeWrhiJ2OOaxlP3Pxj156DfwPTki2WP2VdYHBDvXAt4lvE+u0ymlRwl+ZcftyM/K4qz2emY+U7bKKc3/s5jDJoq2gkkURX3t3ccnZopK1bacJJR+"
`endif