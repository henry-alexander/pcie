// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RYhDmDmo8vSxvau1Ass4u8CA25/dkh8PwOPIc7UkA69bSCGuK58AnSnemd85
7f8Bam0F0fweasCZJgWy+fTrcjJ/Hda+vCrWZPyIqlp2ftDZz+39l/+t7ZnT
7LnVz9K+Jo+ceENR9kkUJpc6NWy7vySR7bqHGR+sSkRtM4V9vWfXo5yTTrY7
bJrBICDjMg4M0xPnGuKjeBhFJNq5zdRttuoUpkwkdAsF8v/rjuLPVFGKMv9C
vmJOFFC4NCCMGudJU7bBIu+re3/n7lurECOnM+XOm7fVVUK8436Z+tloKy7H
JPVoLWY1wsLOcuqd9Y7j0nEfsI5UgPaSdw/JOZdMJw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
f9KlE6tUK2dcpE8vScgBrY9TZQ2tRXhMzTBLwVvo+KDMD4GRglogsU5+0pub
Naup7w/ZA+fiL2IrwLAsr6Fwh0A53oryN5i3XCca4mJr/Cwjj7VrCoyyI+PO
c+zaMg8v9dbXvYbApHdQw5T54mIn8VNW5IuVtsoFzslptWi7qiwI4FfQTj7H
iFiXRVOSJLsQEqkO/3Fbs8BsRlHaTaZEOOHfY+K6bpG0tesQPrITkmOJAi2w
IqE4nPyZGaUez2EN7KmSO+hbrVu3+Sybdy7GME0rXZn7Lh5tt/nbWc4EObIC
NvPgRhiExw3cIv2gScj81l5Hjrqhb1kRuLwAQaQ8Gw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
aAJrZESm/zDWvRC0ms+dA/EpXugTQF41hIs4HiTl1le6XKOibCkXdNPMpmtE
6KvO9D0pqzUjc90gENAEdeEyBkIjlGrMgc5Lpvb3pyqPEG6UN5zDiuzi9lqG
6I9FptVS5Yd2T2rMD4/M3oXq7z3VQAY6/kslCngHzQmtYkkmNy5XZdzO4SJn
j8RfIYrCRuHgXMZwyok8dDy1XUEQWCcQaWHMEl/77CvY8+xZH81+M+aO2PCB
+Gio6wLweaZqG59hbMavZ9GSikR/q4UkALTn/q78iEr8uEEz3c9fjcoKDHPn
CQ6lecB5VbLv7OArauki/YBl/zzAypMHBjwTJPmZ2w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pElFVBx4vkKnpcN+UynU+j9bBbj8MfTmW1d0Y+vYYwU+YRfGvPQ9/USrIQ1O
AqpdRaZZIi0orUzRQyGcTTxeUsyEsKIiL14OHzQrhRRSP5+G6Ak/d9sxwY32
fm7RkcHDyD+Qx/JfIcDHR7yueI36J0aYXcYJY5+0KKxdxneHp8c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
EBovLn6R9dhU0LJ7DilrRpNmZqULwaSJZGt2HpF9Q0Aczmv9yeUf94GdJIlG
bYWZPCgjNmrB9ksQBpRoVXThfUFmMCtobE9A92d9HMue3aEmKKQhsQU5aN6z
GmfzpDL7bMDjEpUAM60Fs+QZTv6snL+kY/NB9wY95L08Txjy5PH3PkoTOI5e
Voqpgoy4RgFOB0N81/jv3gEvIVrXWK8rOI2+ZGq11YH0sXq0kA3AawrqsJw8
RPzDxHylTC0H6/pewiZGIP+fDZjoJDuHCSs/fa2KwDG64lllgHOzsOaJgAVw
Kbv63T9wxUhCFmKWgxjfx+i6Gv7GRaB0aCtnQJ16rOHa/Bm/+xWKrCMZu3yU
xS8BucFGZSo7FNlOnKtlN0HOIk5i+XHPg8VaQV69UoUaf4LxGMtWgdWEDLog
acDk+kV8TsBlndBoG+bNr0fPWc32jyTMM1rNsqX8klh630NH/LTw9tKJmLGq
iQhrxdK2xq4IWs+ROYSyZWp6u6Gs6Xvp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lZrqHn4+/NPPQ/kvhLYFPIVbX69aqMU+1AA336WlXt93/cWlyNsGkDnxm88g
MNKLIEciA/Vjnitzot5h8Ikou440jcyNPYY5UaOLNHtjHhtGS+g9/vyhaVXK
ERNqeRMTCN4lRHofo1ogyFddS06yzfANubLixVJCm5Igefb3R5Y=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gWBQ71zfEfrFKv4R3RX2xmd6BZyWzawhl1jsorOILz4bLXJhJv/FLx5dvw5l
WnIcSxtPeNJEglQJ14goc//C/DtE4V9q+UJqVvwLUD8ma9CondG7lPvlxL7+
l5sKbxIa3W6ngzlkKumIH4EoLqILST4bIfHgK0YLBSHT4OAN39o=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 16592)
`pragma protect data_block
0fJ/3pFB01NF42QaJwhKat9c4rCsPWDNNhvgfJbAqY1DAH8UOkgB8V+6tIAp
KXP5ri+ZTtxK9ldVFl7GuXlF/jQBq2ps013v9bJkWl6SFKkTtCzcYKmy90Bk
pgTNivfsJKvgzuOLV/opljvthggf3JJCCUywKT9x9Rui8oUQP8ZckJGbksqY
kmgfI/JLE2qyv2B8YsEMrioVRXjVaexc0BUi917+O3jpRHkVvvM4WTm/un5s
gmiVknNKwqDyOhxWDFxjQTN2kUZ6Att3JzGZOBJuF10AXAdcpcNdKfpqTgOK
nrjBm3z/nQw52O/xcnrJLaCPjSIAOp2BeHjyBx+RY8PwjS7GXwcdrkcqtAr5
9ZyKJfTo7R6QolhgJI2NHGMDz0iD9Hl28zVqpc5facowj/fwEZg6VKEqNsUa
ZpysLgQC2w24BYn89ZN5mbuNpAZjfc/2wh8ldz4BY4lH00JaKTc8Shsjdpd9
vdrpTh0W/BySAkxMIgkKJKKaBZg/Scb8kiKwiYQmXLHF9k8OY0BCrVC+dalu
A07x31E66388Jp1ieN2GqSi4EZFF+TKocQGuEW3vZrCXwbiZ+hvrZthUwDhu
7Ojn+VOM4+Jg4tlVTSBmC/3wqDqN3F+0ksy0mvsIDtOVu53TGVooxdo92P0S
yFXYZrCjE1Iq9AST1cQcJcheUFY7VAV1HQfZcKcdppHyNt2+LMXN0mak2fR6
qN1SlGjKkB3V9jfHAFSPYJi9cE0C1jGHJ/ddoXzeeTyf2hi9Jzs8Ua9qrCLV
mpZVs0dvyL52/mfq6r5LPesPJ6WhZRWr70ujvlSQfG/10L/TDNNVrkvs2pEl
/H0qfLPxzCRI3L7iYiXo16o6mHGykLsE9j0jxFT+DgpYuV5PGBdTkRm3gQIE
Ci0tmo8uUvDq3n7LcWF8m7bi/yyQXATe7uRkkOD5fVr8pJPZdWjyKerr2F5M
Bxcw3lnMa6vET0VkczFd0UXWwEa3vqXWn8CHgrnTVTHRUuTDtmJ0H8r8UQdn
GO/M0a9yZo+KCN08KrjSjrurzYKMqZZ9K1Zlv7Z2yTk9fJTChKbCEDVz87Zb
sABFsiWo2/PjSHfxuryRPdYD0S2RLjP3lpWK9UqibGE0K6EJZi9pNMNWaBW+
q249tIGjyUEHfLDoip4miM6MN3nxxkHdjMUNm9u+7Ki3yVzMU90a2OOcSK/e
4HffTPZbLsbL7M0cJRbwPDEhiIzIwLDv1exVbI3USurNvbsiKtTE8QRbBKDE
sf2pXZJAGZHqr8zrgAvjJHXDx5idTvWjXaMkfyAL2/TZlytaiNbuAGvJrkiz
xxHf7lb4muSVtBNxMM04In86jJoB8g+jMTko6k8mr8xwTAcG5VnkpmbcE0CV
zZOwHFHokFF89gtUuTon8b9FRBKKVRDVYbDkZ2YTFTZNXHRT8cmj196sms7E
rGZE83iqvho7oKXXEDyAZ6LB8qWGTxfY3pJjSrbyMNDUZA2xG+XrZpIXbjoW
FhO5ynbjMjZvXVCt8aVQ83yRNrkVgEzUThwrYG0EE+v8834uzj8rNds9G9q1
sAytAy9JQuNXk3R4X8nAD7OkzFpjiiqeu8rA+6lgmVJYVKGMJJqxoNBdKFxn
2677XjdfRaU142loYp9uFx22Sqcwt5Mnw4WztKj+oM0odoMRi18Q5FlbpjTk
tJMS+iU77clKIUOUBjPE6bGL6RcTFw5nebPGley/2Yg4VZZlgwv76zfAI2z8
530aIe5ZVIZHUSKxLxZquwYMeRdRCegF26WXjxpC0A9VpI9z7u7r1MM5Rs9L
9c6lbIJDx8TTPC35dDC4hq5Vs6ZuLEiLC6x6EpGQ1Tkp2R05/OLUNFQC2fr+
rUNfGp8n7U1qnYm0q+NV1kGZ6jKTvrxf8vBdEis8w3A4fK3oJBnvLhBMh3UV
Gmd1W2CAiM6QEfmzx9QY4zBX0AvHa+R3VnDMVxHqx2uJmU5UHL2TaL9GSLSb
MxtcSAiIoQWRbOF2X9Y26S5pD8uETGenwlRTdWWxekc5nl/MOqfT3pueMPMU
JCkvnme/4avs9w7zXfDEf4/0eEqeGR2fj/BBsj/hH4Tie6aSG1ZNxFQfDMcJ
QdlSwpk6VX8c96jF1mhuQhZBT8wjtxFlz0VYj6cTHAtN9hIQaeq8eLKg2U5u
gyVeIYC/VPUOZ0St+qD5c2iaGqud+HEhcIaeprY9gpXNSQTmOoiQM+G+kVCz
vRxk9alDrzB0eC1vN2sJrL0aioOwZYglh19JZHuK5Oqj7447ucaA71HhOXlx
fD/oUhUFCAbow7/vmnKwHNnq7UdSD0WW0CKJdezfsdYDlhT1c0sz0a+5b30D
0lOCLeNdOQXKbqPznuCc7LzsmpXS+72A556AZU7Yi50xchjVAVrjlWnTZE/x
xxwBsIqHR47jFDJFewmlQbj8qB0O0PrAwMle+SGc3/Cm6+k2IRJqWadcNF9o
f14OVNwpIJWdRRZyj62YMfgOQc7vKiKwu0vJ/2Bd0UCzztvGTCIVyHyGrFdb
CqbEhjX+HPfiRHCMnyJdCRtK1boi+ouqaLWcsuJ97HcRjEuqTx4FEsCreSJU
sHIj6+QVGg55vUyqFdYzyDhTdNHBqhDvsm7osVqGYQytazHyUzGfYtLFP+bR
bgWWt5x24Uhl50aTd4fBp/v9W9oef2pABSzCw5nADcmbpZPvVX3I/Yd02IQh
GyhEdF/Ifx1/SOPrznQ/XdDqDUIkUePsd6w0cJrj7kP8wDGXnPZANKeQZcPb
EGnaTyf1+7rf6FnzBMHlgf9RrL7xViI1NkjZo/Y5ZV67OAJyjUh++sbuX3Ae
Si5VLXsPLZOYr+Q2wgvSj0AS5RsCrIQS28+wr4txu5V4mLucTu0R9eSRUVXC
4S/biPhCBx+zawLxYbVKUGDfvHqN5XK/MJ1Kr8HqUyXsXSOeziQoK+0EH/R3
nA+VBW/t8ANkufWAOcw7aQm2xZyd95/PlPpb5tx6gWbqYJwNvSADO6k6lxOi
IJmTyxK3MeU2G/PnGT6A8NZaEQ44WqoqqxbEWsMwhEt8HS5/a1g23L8/841P
bVp+5pDhvhlUumfpCZgQE+ZOcEvB33tvlsHjuhi4E49zcsDbMhEe/3m6tqUK
t0QJ6hpz9eovAY/TFne2J8A3LNd3prpG9vR8nQBmYILfJS+lmXKJzFPoOdyX
Ml4GOkdyIJhbQCtU2jDpTTaowYDVUY7Pl744GQA3t+GLdc8+hQIhG6wln0zc
ONuQGCr2QkNNt8bzvCYxjBx6+IG5SD95tbtePlkMMHlDk1mV3KhZs9vDz1iA
midNKLfjQp236Uqno3yzTzO1+UbBy2+rr7HZIkgXFj6CkN0WFiBZdFe840a4
Y7LhQveNepOLckOetqj/nfqgmNqPBOBpvADXIaghgklf1hwm+Xe8ASoEWkwk
AbZZI405ozegs53/Zk3YTJM79GXwHura+ELdKUXExas4QMSz8JGBvLcfkczU
/RJuR03QO9vpKfmjsPs+xfyw/y9dEjEUmh1VdgcTlN52/na9Ik+sGac5HJ9C
qPIfEK/xJJqvk0wMvVoADROl1svkACha9fdDa9r2XbPSJU4Uc7CsYQLzQlQV
IygWIf6imfqSAkVv4zy5lmtq8CRblj314EGzjHF9qt8U8Mk8MMkt5fDzCW5I
TEKx95IumeO8qL6zJ6PYPLVpQyylQ6qeNKJp6BC/G8h04QC6EzX5+EkQ42LL
FmKnnTl1b+BRI2RQq32vP7B1zDAZCaJk/OoudM1iLPY/MS0dcI9VUr4qF8A5
XdeL3DpeAJ1jZ5r0wQPhtI/abY3zi0K9Yz0lHe06qIq8Kk2pN+gr+K648VDs
odXmOa72H3RXH42h/O5Ri1lE1XBpdxd06HbM59sy0fQsO2JBUhZVmlqAme4N
odvYv22bq+49Ldm5xU0XdUA5RlLo1ICQKD5wKOC5RdH9REu1th/FiJcxmzx8
wYxdWW1mom6G8CgNQzlIUUtgTySkmoiYXkBTvCUTtmXi8IfTpPCcj0Twyhqj
Y1IUYd6FP69dOC8gwpp0QMfkMStRw++55zD0kTy7JXwSpJ0k0fUDqGWM6qqp
eaIgYwss5ZAoKTarpg3GwAg0BSGEHwgW2snwt/29ikLSGv/yHeXzuwyzsuVi
4vhfFtjEX68ueQp0wGXrSp78mi2HFgVximFYDc0HawO+1Mr5SYR8hPX2JmxD
eV7HWFMLiTRHLDZcltv16HLEKFUmeEe07D9gZagGquvUV8NYkqEizWWTleAk
uVuneXDszu9FL60TBzvNdI0O8TEt6XMUtSxMdm6qqMrkr+T+P1d7pmJdyZuo
9qjA37ST8K5+Vs6nnW9urfIUNaHNw1f0tEnpQNraNdiFijA6KXKeWH8x8k42
UIVyNM7Wae9C4h/qVSUv4QDLh7tTEO7lOloGz8GviTLJg1jkCRN/6R4nlJM2
gnRIlK1OXioZfb66X6PISrDaQ3xQmPWNOgwgVFmRsTVW6uvWET5XysRbjQt1
iqh8v88LcB8KqTcXhirTknCmw4diDbOzTMyL3SA5iYXOqWL6NKz/zvfkIk3h
wsilbq+wPnbS8CO4ZdYNuB8UlxHazcxW22fciUD15fxlrDG6NFJtSsNjuB2y
lLCpQ9OgqIGSNCfs0dmmdRcQ9gcD6tUxglNKo0LV04ZX7e7tyXbmfC+9Q4AG
kJRzQK5k0MaUNjn7Jj/fBP5W+zhb9lthxKPCRaanTF2JfR5h1by//w3eD9L7
1hqqxyWH+1OVQhfYRB9Zd7LzYLKUm54JvniukRaGarE4vjqTpbbtGk/tDB2J
CoOs/+xBKr2tGMxKssrTxsHpayYW/klEwevaNRGU5W3nHwFOWCVfvBJK0ISM
+XjCHrGUZzzuaPZhzU6sOie7qd16BxnGCoKveyNPbzl8wZQzIfH9dKL+67W/
tYvl26KcrQXUwurrU/cgsCsjygUYXfigO+b96Hxb6BONZvia+Q9ncOPGwLQC
BFdLeg/raFL5h9+YZAdV6iXt+cfpgGAY+EOcr1qw+qd++VBbhiyX99tBW6fI
KTliKT+AMJPi3A4vOkVgqxcc0PpPlsUgTZe4i/zwlrQ78/5jFQHLo6iNTQO0
k/e4sgtE6RP2JofMifTuWYGBYAendJi/FONYuevAbR1wGqEFKxQ36lM3oIXY
qOiuhkqQf4ZpcJ8H8J60nAVD+/6QGuUcVo0EN6pSjyYqo6/Y5My6r++wE6S3
ujoUmg3QTlM8AqTpCD7irwYJPXsypGpeIoq6cjZ/g7X7z65ZCVBrL6khB1YT
9biH82vicoeUpT/NZRTVriZTe1ms+FBhNxb+e7LfPX5FT3NH8JoFKHCAN3Tb
iPGMRUJs7pyvfR5TO1DjIwEEtJotZjOfY4HRZzPLnG8ji2Ut74FxmsRZa8XW
qQXDuF7BtugGAojDcyBZf7zaFmLceEhULTJ672WFkH3W1mkasomHkrgCIjpy
79lLwJ2L7vLOq9FRIqvArogS1DymFnyhgu3rfZwkDvq1aXS3dEuEhZQcfRWe
2qF52X90GjokZpwpLH7HdjtBjkkrI8BXi9x+07dGG3FQ6ZLMRY0Hwc9MH195
AT1lNro1h98VU62e2cgw+3aLKPUqsreM8Tw9HjJv517s46u6+zK221Ted+GA
qgta7TlulTxtd80LdpHKjF3GV3ovI+EWfAM1cZ6O4NMccXCzePopCHbOsggI
U/px0syWi2VW9sSuqZc7i6YVyo+0y3/q0ITDQPRZb/WbKoZhdJTiO5RTryz5
kaUebcBAHWJA3r2pZVf62oegsf/IBZjHdKwQX1XBUUskJ16rT/xjER87uI3O
VZDdVoRECNipIANaBA4286d6UymyelcKkOXfZgtrEfZe2M4lW/BXdA334Ept
8tDg3fJN8uZqiDVeyLe9hW78R2rq2kc8j78K19NHZZ0t49Xf5HEkW7z0JnPi
W7EXTU/QaqMvdehiDch9RucYfWyFEGth+lMvBUpUSIfbtxKMkoNA8q/tBRPv
HqPbk02Q2HgTKfhXTCUQ26co76trX/nM9VdMKDt/ixREn7QKF9GmyGxvgjI9
vo6yteQZZ3yZUvrJ+3DQWm1f81RHXJhWWKidRzSXvpM+8CWxGBvOtF5J9C9I
RAqZjIjoKxPhPMbHhB+6XnbnUWbqd7uAQILCaYkWUIXhWVQk4igMs+mk1HVR
EY1/Pvkv6+JmOYej+Z8cByThk0LpDAAWwfP88exxuDR3HT181VamUjVb1Dbq
Be6524YZtgy7t//LV7KwjmUHW3Kl90fNSFH8rCWo4IF0kmy+JmBvOhwefzlp
swcwwrf07pAr3+LNdGhjat2qGlt7G562trQJICjs03DQVvR751/K960/EUi0
Q37IgE1rVdWfFftRgGbXAx3IE9IU79/gAFquXdEolIwPk21ZNsBVWmepokPF
m52kOQQD+8vD2BufXyfNWQqOTEQoxVZuzTTDHmK5t8nL2nKJgKe8HGxEF3U3
nq8XANmvyDn2LGqzJDGI810aLQZnNAgy+B01H340HvxzDD+ocCm1Vb/zHMCj
gOiLO44azmitx9T0nYbmxBvUf1Q75sMgsgpYGgScjae4tozqIpWvt1hZSi8J
z5yiTk28h2q611w0gtaY7WZ843prBBRYmZeKHHHIafW9xk6n/chWkFjWd7Ju
TrN3PyW9ji9VJsaX80m2FQjXD/sOXvzHkfZfrEiQ4YxhSvV6YwD4E90C+xZm
gqPqGTrX9rt0CrKxFEtnldK+WZISiJBcPi3G9x5xYCFWCNApI0ngON5LaY2n
AePFrfVcyMwuZCntXWu+6Eb6FGzHcJoSRzuztyizh+V7V7IRo9+wdQogPQrv
ZjQX2jEbClem3zYzkiaGT9OoFGTp7ghjGXQAt0Ogckp9DbI/0250D6+dWokK
vz90/TI96jYpXZB4Rn5Axw788u7qDn4uUu6WS4INORDC8qZ+LOB2o1S1Qmeg
XKTLyAaF941iiMLqq2I3JDDd5UJB8GAvfMJG5Fnf+OvclYs6jjM9+8QL20eu
unVfBxk868GPw2sziSbqu3rZ6CCqgdEBvUt12HiibHbAjO/LGyinT8F+Yvpo
C8k8X86zY1TCYlUD5wIZw9Bi7urLhBB9Ne1qebbnvwzKeWUKfb0yIyj9oebo
+/7CH6x8hDtR6eDTzqj2bw0Cugs3WKC6sFl+egFqKeGpm4wlWcyPSC7nSCdX
X+EeEU24niB8WJ5unNEZYBF+KIpvBrw5J2yKnFS5xQBd/1/XTiuvmHDhvrl0
4aX5qg1tSkOp09Ca8Y/UWm2yRuijbPIkqmoNUQ29EfVcOUGMRlxc+EN27C8t
DIuW/48hpX7DT6QaOaA/iT44WYJcZHY/nWwRMTvDFMCtgv1hZ4sFgHvoPjfl
MWHRA43IC9wvNClKp5EboIB6E3PTELclfQV+6WjDn8EWJ/JBeSfbzWUlJ1Sy
hC/b4/t3XHgiMWHpTVMDlqytKv+HQi4wfJq+W727qRBtIFp0H/Wjk2lyiEsG
PUmOoY8m/KDVxrJMphebrlVosfxsGyog5pp2LYuU7skCHwuzEDw4islxNPu3
ZBO5LRL6c62LOKQdRxlrruE7Ce5zbWvM7AXaisl0D/3rpRi9FsZqvgkAKnCV
Nvg0/o2o0V4Fg96Ko8TUj85WD1oUndl8JoqhM25Fg3cFQt3lkFqD+Peqin+E
AYQAEhnoqHbTPagZkZP0p2dcEAQ70IIkUQYortaDCzvE09FJ3uAliLkcv5CH
tHFFeGsNte870h/9s9ue7aFSC9sEwIheNGANS6q1ezgVhIzgErMJggN3qw4u
wayXx+ze8mNrJhtQqsI7UeyvZqRUvzXDSwLBIS7699TPjNbV9Bi+DoFRahl3
8I8vWZ3iPGMi295I3+sp3Zw96BUitJGXutLohEVQ4lV/YypoTfm0v3XKMM/G
SnjZofFOQdJt10sUGLt9rmvTZ+0iHg30AfTRdvSSndONQIR+Q6gS0V+Qhcxv
Je6FilcsSHu5v/oj+Mdyd8gFMeH3eLDOrFA0X/nvIpYTx2NMhlkdOcj3bc/A
/HOZnngpsFmsBZrk+psSWlElWCJ+Kdb4So4SdctOoN93oNO6AlcEQ2F6WOL/
cxrBK/N1QhBi9Js5Zxk72UilIQMnUtsdEGU5OQVqmtZwEMb48lYPXND2tyuv
ABAw1hvvXW2I0RHKgxLVOpq7NcoOcHgptx6LlxszQvATiPuOW0xbTve8zsLL
/KUOE3zrmX/9/DSeBl2mKAy0G+w7bAKZtzUndBazjdH1rMfF7BebNjQGEZa4
WyC+e25/8pO4bYKKK2GzJd073Hh4IZIoIc7dDy8il+sB15JnerP8UmTnn9U6
TGoCwI3vMzc84WG+kjYRbeHsAYeSCtLkYzrwSpBzKAQ43DLO0vVRGfNCoTvP
6xpSDCyGTYeI3GMTM6IPC4xSnE7J1KpCKFUL9vTtQtZVpydYqJwVWyhzWtAG
4gWjM3kNjQobtbc+EwuoeKxBbjASLzVws4zgJWuLR9O2NISabNGZHUw62Das
b/Qbzlh09J1njo/j2AvDSI+875pb64Tb2v3Qtyam+BJqmq/NZ0bFg3w3wqa0
mTfq+e2s9XDD5MZVW/LKCZSJ2Rnbn+oJ46sRceC9cD7XIv2RGWKhsPZZsEF3
mhQXpA76SgvCkgJAB9BDr1E7dmJgQMuC3fXcTDraErg7HzHt9KgOcH3fkuu8
toLKsfmUmr/YYRNczfuvCSEq4ejXVrXJJgGnZY9Pe1fJgkMwZ10Gi8xi6VgY
pj92oZVs7N2Tb+TmHwzYPoCUtTgumQsOyiwqWmuoz5JOYgEk9ggJeB9RcxSZ
UcHHC7vyKKaRGs0rb70m1MlpP+iINCnnMmiRXg+mTwb3jlwFa43DGHi3xvk4
5NiHLTQb3nyqRAfuFDHGFwE+svyHGW0Yn0J//la+n55aTYOjHD+65RqKUXpV
YgXtpbxClQfS1auK06Lve61p7koOONBm7yMyQ7QvGYHC5e1ELMd6rbru185Y
ATCwZTaBwkyYyFqBfGaCGKxBhoWwXvZgl1HSkKkQYUWHGQoD2cVg/poYdxly
Hdtu14K6toJIMXKbEXpJZn+biDQ2XNxURy3kl1s590X3sujSsuk5PqWwJCr9
qGICicpBmxb7QeZvGC8iuYZ1dCQnECZKoBFu9dewfZ4KMQdNoRFqTeJwycUc
XLSctymv3ICcqOLD37z+yZJDbqTk2W2VNbIgoXl9OLPzX75a6I38u1Ig0LHs
t1iNojzgs+BBI5bo3kB/mNKA4jwt2gqPsInkgogoRuHly5vTu2hyy1dJF+gK
kn4W09+WqNQHjHs1mByoppMQ+BsN/RC5dxAb/L7qqF9txNmJ7Jrptt+slclL
NmZ7V7vmFk/Od8/jHt3hRJ3/WPUDradVPGi4nLF3+EZUV74zUxEJb6ifWORx
bLjphXoml02vQ45mUXx06YErAvOaN6xrhUFzaywWEoD5hIeNPKvKiMGeZTMP
E8dvFdT6yQwxd7/v2U71Ay9wQWyelZN1zVXbTvBPHvV9tq3Fc2N4sXRk6jmp
/D4XcHIcacMGZt0tAw44ia/BczJyTVfkMRH2gJNkc7ba5fGtxCaFMgMmqp01
vHhymyMQeETCRBbVekYTsoi9riceILqUjF4dXCp8bn0rfnGzeWcQpWONwpKv
8hOF/QAMOLpsoH7k+iNTGrlq8x6UCgMFrdOWlykJgIQVvOvhH/L2FTbaPV2Q
tao6+dui0QVbsYTiGYpmUb5q7SHnT5cLb149hWesUGPKmBpTUmw0SVejRN6j
pZypFSkjSpRVQLYRsshawgI0FHpzEp34lGGtNwANnH63e5+rAZ9maE95cuoo
iFh4rn7rqAejJWmxALIgEIL+RwN2blQ7LYemOYwmlTpi1iAYy+B2l6lgeLVt
vNcs/VByrl7LCslYxAhyWj6ALZqXmY35ogzAzI92wAbkhtS+10VLhwsyGEU5
0yOyR0mcpGIW9Fzm4gCFzfAW6Py30xgx4fGlbKQKod+SIZidAkzoyXHrjiv4
Z3/VM531JF+jN37EXeBZCUlwtid9GcR4GQYZTUpJTK7mf86neTDdKbZ3z/Nq
PEAdxRb11WXj3THyxjVjAtTBfraWqpz82sjPw7w5BwgkjBH+/7GW5+0xnhw1
Myg+X6lVTrDvJ9ZnT2uAc9S+5p1ZVdW7I/uSWz1zqpG3eEkIk4UhgjSZ9cjJ
fB0aO20zCuLMXZMjjBCPVEG4uMlhjD+QI9rXcmxCtW6U/tFNv1Dtj59wxov0
Cwt0GydgrZJkzMI0pMhLe0bzSQAV240ewvHeqglWAqV8sxOBhZz+A0IXtpgn
3fEcdJJElJ3sjShW+yURGUBWDsyTAE2qD8Hyria6Dfl8KjA47Kj5s7SmTtgj
SzzsTfCoayNXCgFmCvTzPQiiPt+35x5PeX13YnsLCFyYgDNHnG2GFTTzcdPH
HbcJgpIIz2R6bcZHCs354SYSzZQFmBwM5+lUXiH+JfqMa5Xybd7aSJXyw/32
OGFJEoqPx5f+inGAoPbYffDpaf2T5NYkd6YFMhPAWLswtP7NE47fetpw9Fqc
Fd5KGG+GE1RznUxgolwVC/8ygOe2QWnGWF2VPSid5bBUL7ufB73sCe4vmNIk
EmtblpKVOuGmwCC6hk4e9bQiyPSr9ZigOLGODAILmau5YyCjIWj8+iSLCNWy
/vUA5Bk3GUyemrhTvmrzmmwIny5uANXf/gFvbHRTk19CJASjmSFVgvXZlG9o
sIElVxfQaemsbG3qUciGOtzXrOOOra3H3W+eCktZ7/wIfd8pD6RoBS26Ts9d
cpq0ij1tOJ5QaSsD+zklw+Y4OjT+nEpaybWd8smQDXMyKjfbSPw3Nj2ZlG6B
AdbSBoUhOicevqPhWYUqBzBXfiVc1QYX/vYwVkNZYTYwGSt6YCGQCJkxlVLY
JXgwcctAkcJ8zFNGaALuITsacW27PWjuSYk/NhP9c9i5G595PRDuOt3gP+fh
dTuKEkRkZwVE0Zg+atDk3kVbgdb0L1iaCEAO9cAzF/pejKFoIj/+3a/C8z60
gRLod6kSpvI9g2ASs4g2G746Nz8uJQ1kmhXPzSfwmqvx4YLudi3IhvKGphNv
QwZumphHDP9CyOBj9as1dq3qa9uECb3DdclNNqeEQZF23lF06hsLSVxgOL2Q
5Ckr0wqGMDl9M9a+Upcy1h1X3O6H3VYOYgWRVXuUxKGTvvXJUVPNJr0UBBuV
ADSB5GfaHaTaGIoVtnzczcqbx49X+EAtXK/MkiOVymiE4RUBvYCXmB3xO7WN
svFhckw5iYWMin1aHYtZTabiXgXkfeajW7L5G9G5tdIJX4nlzppxKYov/SXS
NA2QudWdgrBWUdIL3XB5miJmwmkJnjTO3gjr2Ly9zC4ml+XXsfddX2qkLLXL
kFeWf83Ij1JMGQeI66jtel7ZDOLqRzVGm0TeZl06oU6jeQ6kZ7ZlPdFiKhYJ
Qj+s0UknWqnTnUOSmTrHXh90wY1iwmg7MEWiiKFHQ35CBHlqOIhWILhPl6IC
r2MEN1GvzzE2QFifhVs/q9PutV95b/qCcAtkifURKRtNnRyRE+1ZpbQRwHox
JiaXnAOHxxBeNrYVtWIcjDAG1PRY2hD8HVGmrheySvRwEmtpm7YxVTjhmb6k
p3sVpO/1layYA2FfAfBP8WG200HWoXTGn2C4ZdCvB8DTjsAfi6y0n7F+Mwtt
q7MYwZxd/p2OaBQ7KsfpYHjN6OKcNa/jul3aJc8MCF0aAiZrpC9LNs3K9aaq
1fuXfQnSJs9dfn2F3oUSyqxxqyDjIPh136OkfA+uOE8HHjC6wp9KjnuyGar/
2zUwMZJqI03o3z7wgC7UZp7eYdkF5TlA2DIwcIPKDfTGw0Iwir06NteKiHFQ
EE1ovkoS38x5xJflWUymoNsoxRF/1TQIntvpknY1zjvNBShDwPd1hi8ztceJ
LzafEkN0IYWzs/oBKGBSo6LtMy956V6SOInK031xKpQi+BqH+IkOMh8Rrg7j
BWyKsAmkbh+Jt/0aK6kIREX9Uguekl/QqLqkpAiXcSG3fCkAmhOIfriGGoLN
UlqR7LHvbDm1A8CY3za4aIHXM3N5W3VMyddNH44saK739rcK1Pn9QIuSXciZ
NvWwv362siNtIfv/ITObtSjyblp6Jrr5O7g5mH64AGQ28ggQq6W4b2+Neqbc
ebOHqEYInG4ZdQ2k9ql7kNa1sQPRNJ16UumxjiH3j0IBYV/tfe+nSlSAXbwB
+Qm/aOEF/CePp4YMJddlBlR9ah+b2RMIajs3u4yyYoQpWrZ5Fi23FsHYBFLW
Tho9tX6WNir6lXd2M5VCfBGkg9UjHG16LXhpA9Wj1Rhyj58CSbNQFuicDaow
Bt8QMKiHWhM4kquWNX2zRl5gtvh4JCXV21/do+lWLL2LssKy2G3h+56zEybd
VWTQJmVeqAARzGc4GlN1jEFsc5VTb/APzIuPQjX4HDmJKPWmCoygFNoB5azb
6R6f6lkCEkk3Yuu09HrwWXHdOAWWhZ9uMsORnvh6KNdaFLAI01dtzwgAGse6
rylNR8CENBYXXO4ct+h24IXA2v6EveXCHk/V8hGp91IVYai6g/QP0pavqw2/
hYMnHJT/W+Y8nTcMdVSWZaF3u8Qu3k9+kkNm7vAPMCBnky40tU+crmJBY1qL
7sXS9UGeItOfTeF0FlONOpy+xqEtsciAXTFPzMAkM2BNfa74PNShFVR7950f
pTu3YtTI3eDqjhgUc/6vnsWMVco8f+CPDdJIIoSRSKO4ruA9IHMZai2MGzqN
QVGV+J8B4PZFTrt16WhYgkNFbHKOY5jZVhFhdSnRfNXV6awO0TmAGEYbUHug
UTma06fRw6qoJ0i8EW7gOPi+xoI+A75ecj6ZuebLv2uAGS2bPQzE/MG/JqFO
8BIDLmUCcp3DKvtPyGmAzXeEtaXgdPr6GBJ0iQUAo2oY1haxBbQzan7tNytw
1wyYYH57gLI1ZDvTBisNaEHTbP42E/JmOA0NrP70A9Yz6+lfjNXAXm8ibVls
E6P8psEaD3pMDIiYFNW+vD8slPz+8kZw8vbadM8qoDdpMatv0PB0okfvfpy/
STWCmHfNNRQZ66Kri6eeFcSk8ZRayhpgSVnbiZHiv3ayg7CxA8+3v8cpYJ84
h6Hk+6B26UOoTeGfSDCMsS//WeohItWgg19qdmodyBtz2AD5kpLG3a+zY7YO
A4DShVyysMs3evmdcOq1F22V4dNvdfYAAlWFBvg4IwnZxU+7ar/e0cGGbHaW
lMOA2MeYZoGEwK+C9KKkLr/QJ0sO9a04UFOwFqm/dPYDzj2xJNTpQP0jHn2B
OZyy7ZG0ba4XiClRUNTnPmC72rv/g1JP5Z14joxmgmiIn5IvbfmQjnPyDtgq
NplWcrSkI0768MZ8XkstV214d5Klte8JgL8Kyen1qkm0F5C/faz75+5xMr8c
gcxgiLqaIQ55biuNGKQQqVDJDhChiqRSEjkopKrAc2075stAXc9S2Exfxfb2
H1Iu1sEGIXppWx/VcUJy1INiZkkF6grHCSBOYvG1bwHvvMKr71KVMuY28egN
8tZ+7UJwXkbOZku0he8AWckXTTHlL7X7zYW4Bect1rUZ8eLOSVa4KzHP+ITz
LKFGeW9FWakWnqJGIPssANz0htx+yx26tFecdJw2iBsdgP/CZSeQuxXOU79J
HrQZjVH6oT1zf5bFNNO35nDBOll/x3n3AC8ogoFb/eyOVsWWNmHG87dmLTLu
nI3PfrBB1BA0llbPODuRTutVj4Sme4C44ZX0cY1OjBcWwfDwZVcRZ8FeLnlE
4tNEnw74F79XBaNTErZJEudQqIv6MXWoqfeGecYyRN4UiMDhUIRNgPNN3Ynx
cvxFpH84KO4/bZCAHbgGSJSH7meTB8Ma1SThzzFeQG/tV8vN4cmDV5foYBHa
42Y8vDMsyeyPOxHXqod1pfLpr64s3xHF0DjT3v9MBM4tZG1Ep4EvcubVt079
0/2+ux2/jG8yo3fQUVdoP1PLmkUwIQFtPBkqah7aGWnrcwzyYmKKxE5lNwh3
jzgd4ld8qDfEK7v0J8fx0UleDgHCr1fZ9QP+v8QzOEOMOYzeZaqbUv/STYYE
3rqNlu7bOZYt0pnnpUhkQ3O3S+/fSv4Pl8ZOIGFRIUDjNl+3oJAkeCdN4w69
13ZVOO+mV9M9TcgTkE+w8kB61nwN2+M072kneJEXiDVXwOx46BeUyWnP4qGQ
rozwBd4LYhiKrsCzmulEG34RxN/kWPeVcrNVTXufpHgoC78Dr9KtkYpAcNX5
Vh01sPiuWZi7gfkQcBiVGdfKmvwMvH76SW09VeamiI2R0K+eVwatbSGFjuqz
KY+50dRterHbE/WPMAQBxrsxFj0t0kMGH9k37vjsQeLWVZuqJ+OelcwwllHh
BigXIu3jyZ3WY/ys1kTQJsdQ2AFYlXHJiK+mpFWSCRXPp9Hth3fx8w0z+puT
RrsY3dxskXVaYK2+4ERwFYBRy7WdvtZvasMtE6UPXbIWNzqsE7DQ92ME5+HE
ECW+UcruFF9GDtISGeHwrbU1V/KKzIVfY+6W920cri61Arf93yTuAh0VBN1y
/Zng9L51mXr49ogAYKLF0kORVGUOBEyo0b43V9hVOtZcq//sEjW/T8BLwTV1
mVmuPWYNT8N2r7LCbUrZON5+LbAPrAxdZ/wv0qjbpmqL+Z4TGxtau+AH3wOR
bhigt9dvSG6KbblxfhK+4+OH593z5Kjgdr2rdRp2unJFj/J9n72LCLA3IgFg
KyppuCENeMuvorVjR0mck3BTsjvwiidZ9VwWS4YOXet2skhx7GHFaIBcqy6c
9TFwG72hox9r6+AWl3r1a0sRiW8EGEyhEgB6vKopP0Zybg3SFPGImBKx/f1l
XdCq/q8tfbyzVyLeWeali2VOKPws92SNU01P0Z8PcIXl6cZe41bc5I72Sz+t
ZBNdDj3Iz/pwqoxxWWtJFjB1bogMwzLmUmsWYbtqRrft9jiTnPH6sSwgyMJO
8lD+CZTKyI4ZbWNeBObviTnW/EsyY026l9qOJMGgfbdSWqRR5bxs+X/74cpc
lJm/bkYu3VNUSps42y8cabJPnOPykkr0vDuCQWooQP11ljui+FtBxtrAIMzO
84hvBk4hc47TQAuwSxJw1mUmVtHERof70fmyrwT/qyWchc49w21rxQW77lj8
uoa+CdB2FsioNdBN/pEOrKv+N4RDf0k6DXVbwCUSnDA7kNXmlLq2pA2LdIPP
P7LSArxOiNSrAcQA+vXxQDFPVhbEsRHU+5w/hmaxsd9ykB2AjgBR3BQN6kBx
QsJAttaymqceDohdPc5EpWW9Ax9xY084P0CrilAH+STO+qBfZ1oevyT3TUBy
w9tNwqWl+X89S3f/diUvKwT8Z8gb7YDO6cxH12W4qs0ohpISgYWxbwoWtAFH
uTF8dlOvny7LjSMKcdqpaXdNYjhp6Da4Pld8fU+LsVoY2apg0GS3aabPYzBN
k04DN01j7pEROhHHxhPZshRzGQI3SDu20XrFTpOPHBMODMtTm1/twdX4LfRF
bBUITKKyh7p3D9BdSFHZE/3ct6juj+NhDhs7LpqCp30WhF/PU3L+v525HFdc
IMst2JF6JI+B5ksO8MHUZ7Dk+F+ZmvJF+nw1jHLbv1UK2T/ipS0O3q2Fbnu3
vaLGaL1HcFnf1nLVZZuRgBQEu1D206OCiDbZ/aOrCIOD7gi4lvYKbJlG1y7C
vyNIoHbAmJjVuRd6FPKv8rAKFRniK03Ag/7jW2NEZCEDuiUdatoGajkecuE8
grYcBTt3AXhWitYqbBr87xteJuquPqdW79ABT1gEDCUWoJa5QaBLhSMHZu1L
boL/pcvosekpjHW5ekRWMz9zWDI8AQIHapIFgt+xTQeJdiyBlR49ErT8zT9R
kn2zRpMsL4HBvvxcckjhtqM2l5xgkAa4CsWlf+hpe8SgKwCG45jDynWHLfUC
LUPvSiUg8w5xPGmA3SzzzWadLwIceBkEz2fy9cAUd9cAUhj9GNaBSVVOSzpN
RHxK9gG/+DyWShbjwWnkB8F1SSthjjaTwA6vd7eP9LZPnFe/+rQwcsUToAG+
I5iigvntK4y0yC0boOG9mve5U0/0wt2XVI8dN0opL57zNotfA51OKFof5xPB
GjBftuMSIEWmWG4P9ADBA6ZUpEVFZ5ohKjvN5BzxqRO6dwLByGHVr7rJ3xTD
uL9aat8sRLYm2jvcFSM7nXBWS1KfjSvNu9sKJVbE5Ixge5mdcy2S9xD5wewE
kc+vCr/Z98NCSgOigI3/RjSbMw+eLwr2eS58tESpGzC3TSTl4sPkV38SCAKF
L+U1m1nBRAeBC6VSSklMMTdZ8xhysxNFrg7OGm0OA1eXczBzpIwz++A95Rvf
8Aoy190S6y76/CTZXSdIUVTkg/QS+DHCnCMqqV+oW5354AdGqzYRaPpVaqdl
H1NqZhFc3Jhw6xvlN9Yi733Ul3CG4MSh4B+PEzxMcZHOtlGY8mXajGdl3RbP
AC4Ez0bbJsDRrcpk5mqVOiwbZcUx+x6K1h4H/6ZmZwnGdUwP7ORCMXo/ZbcX
Pev8XSb0dvFtVnVyE6YnM2Vk2wJAohDHH9uYWHrJKhkPrJNViFNrgb7c8T81
GDOgdV0K7oZXLWDDPsV4rmS7DSRo/A+MxERunBJrhA0RAphneNzN9zDDIH9O
uaEz8Ik9l5JYKaTu4h5U4rTKY8r/wYpyokQSR9pFrNeoeUfHoUjnGpjdRUH/
kcI10800b4GdleuKWqFd1aIQXzZ8eBsQzin9IsHRQT6kzs/GcMWKPbI+ipYK
SGSd73h0MD1yo1nAKq9vkx9ImpC55zqDGhYt5LPSY9SOqEP2yKE3BX+axBhR
i7Df6M3qZDhWPRnyFXN17bpxqe/+W6g70TihJhua2sADoMXmXiGm6EYAO0PZ
woLISLMclTcdCZf1xJr2KPWk6Djnf2GPYM5qQDFMS3fjwKyUwpgq0lny4U4j
SwFuzEZ+jbsVtbV++N/8Z/Xztyiwv1cA9BqJeC73xfRjBY6r/x4itN/o5Wtr
8jykFXY8RWBCzSGc8JGZLHVtKgoZpASAUMM5oC6jDOqubmhzeSvatG1CVQfF
8q815r8VY3EudNz/BbJNQUG55irD2aL1hct5Pg99Cl6pbRo405zlLJSn4xxQ
8oXdGK3zcnsmiSlctMoHDRXpVBAuXEqvQ4cDxYz6Tzr0hWeAoUYv9Zr1Ec6z
bXCz/pOM6KC7q1vLyDgQF5K0/lAsl9wHLYYI3sOl+wWra3w3y5vMP4l950Xc
f8esQMuuP7ssI1LaRSca0uXWDpETb6XKuBcGbbF+u+s92AXHDPaRLSPty/c7
AWaWYLrIWDycfS3NQ9XvkfXZ6M4WZuNE9EcCU5NikjVjP9AAH9lLuo8pPXrh
il0WT9IbVOL7WP9U/NeoIGr8AlALdluSDKv/FiXS18R5ZLjPRtX576AeBZj5
IqVIgu3BIOfiJsyZMt9I98Lva2iETuISWnkhbjtf5aM7T5aolpC2wy0n+Thn
xhSYI0wnhkWYNvUQ1NRlGxMD359jekwzYU20WUgVMykABXaoLVFVjIjfOYIc
BuHdVRhnvo2wZqM/zFvXUhCCsFNMsUd1zskQL3/QK3Sx7KRTyZ5io1aAYBfe
2Zh5um1hTlw+V5ZlZi5dK20dIf0+2toCwKwJov+Vb1Wtcl1untT94EFIIAlV
E2O0JljVzx9AGrkLcPoEeupLBOJflir0odzhd9svMKC51WCiAL5H23+X7BXN
QJw6whITXIryxGrU2CcxIrAU0IWN0rUmHhTK2OtuME0E+Lbklq5FZ3voylvt
o2m4SuQoGt6cRBjYvKuH4vdmh2ho0JqJSrL5AaRf7bBJmOyhP0kDXHG2LKAU
Y2kIe5HvWJg7aO14v/y8CQIU9tT3cRacXbhkdVjSxofFh0rlQniQBauzQnKu
vXceUjDSixoM3IePdpudqI9n5dsDy0lgxhxaSQD3E7orgLeeKO/lkrEzPXHK
OwuamyGbzSzufBGLSBZ/E68BDbXmZUpStXrJMQz1S8hROV4IUbQQjzaAkiTy
svCO3X7xIQDf9f4p/nuR21obrp9lSgOhVn7gUXM4Lv+0MwNBdqUiNY0Wq4Zv
dYW2q7fw/OEx1RNwoWEDRUWIOB563Eu2KEvhlmSU1T2HnczdI3wk40Ay+SRE
XzQ/8Gx+bZBqv8WQ+XCxNchTj518VbCK2EZSdGlzWkBoc+tqDCjaEjzObKOR
sSNK7iBKWSiP5w1a8VXBpxn2CWrUknq49Tr1rkWVjEK9mOEnVLsAv0L+7P7h
JK9sFdL7Exen+wNZaYUFbUIuqF0GpAuriGGeBboteFnCFmgjnX39S7iIMWLC
FxXk7+y2+JAApn7D+B1kt9vr2vtoKyUmqpH6Ut1nz1Ai+A39s4i4cj5k0SXh
zgzCYHTqfEXzaIxhddkF5L5U+bK5a8rpFe4igL+TWqFdAoza9XL0N+KRGytv
nuBN3ZdMFN9YigDDjtDA5eWNCy4S3Wf0FEQJarJUupgrCDAlzeM2ufIxTgqs
UM8qRzSfyZYx1Y4bKyxm87iQMpf893pot/lCag787+DFYOYpCWJSULNqgv6X
V2jQuUtqUHhMpXNWngF1CIv9rT5jgLKCvVdg1vAd1+UDzRoCZM8QZbnqcaSo
DBOH2+l2Ose5KjfgloyEQ9+cO5tRfqmp2AdqJYFmdvRTDoKpv9TOcukEyZzM
SiUN5ntWUVzS5m/S9M+8uFI27xDIl7JdrIPoW2Wzxj8PV5PUncF09YMlZy+x
ODKs3zXL/oybj2zC2dTxMmrrgopgqo6Xk92cmtvc0rg/yeI3U7V08kgdSPCi
oQu9ULUPm0dCzRTVT8zt7CL66n6cxa8cXHVtdGV3FQZoJ+r6A2GfndZ8g8Zw
QJUzT4cwVlTuB+CBFPRwy5zeodCnPSV0DICixIgvT/R1+LYv0E/zK5c6mly9
ezgLEbpgHnNEpsN6ULCB89M5DbvT8c+f/mO3ax8AGZ7y4Erewv65Uq4+EoUH
5ueOdn6VEw3NAowgF7mlaV3nwVhXz/fmIlseGq8ZqpEAmAXKfn4ncC133IcH
QpNXTUNxTchFziwyyTQiBHJ+fGviDeXnytR9LP6/wiz+UuLBogSz9QRz71S0
aJKO4LKYYygvxvC/dcC+XHnjCKr33QVEn2LY9zjwokD+O1FuRfj6Iy3S/KTi
KWZBz++sf2Fyzg02rMPDzILs/aXUzdl/CuB+5eDWafvHy/Fo1OEGvjM4ppjS
7dKKY7lYnKYob3IebcJ7yzgKyF6SzmWHS+SaJBSZC1TtfW4teINk8q1jtV61
/na/6jrkVAFjwCj5Sm5OIqgxIJVYGSqovvwdG8kY0Fr4seW2vJ/RK7lNMO1M
MkFueTad4skdBob7xJBq2chnv/5xzcKr21zitUIUXPWH5phSfP1BkQi08GB8
+iVsA527z5MRwnklqrDo07Hizlxs2zqpeiTKqO+LB8UraMb9a5T5n/3lM5oU
dnSMMJZswLvHDUD7euxwehdamjoR6zYfIn//nCJ93SAiPufr5Afr6Ufi19sE
tZ9oSiwVLTtgBhhAqXuMwBYE+E7pJk0QRRhokmUwmv4i7nsGTGk88AZfvXIw
jhiN1HngM0uzadghpUUt/PzIn3DSm16SqkgigOyyKyJy+Vpb/e02ppPAyg9Q
rCPL8M8y3DzM0l4rglsgxfPC2DdZ+bkZDqMXuL7EguAkCA2+YeMCWo0Nf8gk
pyP4bhx20Kfs7a5PQTXx2PnXIQ/3Knn8uTmOTHK1vHJOElNe8PXO8zVN6xn0
IfqrK9gwqRHMuJCcStjTEhdVwnuH2+nHaGzvki3cmq78gSLRyYXakixRrvow
sJcGc1KIzhOpKfzR2YbgWbw2MBj+L1sCGw6b34dM0fEEay/cDHOqewKmynZ8
1s/btcrU8r35JQkxIBHUSegiX7eJbQyW7OICZjGhMUGx+nGNautHAOf8R8na
T3iyZcTBIeseJ1XfTxwyvS2kSBG1ZOIpqJ6mFAcZezEjj/F5mLRWIPv+eYpI
LF0idiU0xGR0imOvMEmliPDDrhzXjhcge3gYVWtXy0uEPkHllN3NPeIWjP60
N/vMIiKvyRRioaFKT2b7MGJAJSvFNadzQspB+JQChYION2J2kEnLx+2Yy6qt
Px1t0YJ/AAj7B7y66cjOTPOvRFVPj0Qpoo6eX6usPedwCWXpu/KkTcsENO+r
vydAAa+iMjBzqQtn9k9+0q9pdhYOO4V3yaHk8O1WzCwKZVTJfz/ErSKaWNrO
CkdrjP/w+E7QKfhvu2h4Jel1AJ1I/Jhjxakvj1dBLGumtvzRqZNVwpExTmZB
6fEMaTCVSwFRPBE2wnUce8TOeVCEKEgmh0RPgte5Use9XQDkcTyjs4qkjq0f
LbHPW+SwJNpQ1ul89QNd2h6ozXJeQJN4xJqp3j3OUGUlgsuUJbeMQ/2sLgQq
fzLJkLbEfvTzZmfCr3WoI71d81n/ykoqnYt5my1sRVpjImtTqcCTK5/8tltM
ltLRnKhiQVsRhu26w9VMrGolNb2qHX4u4yGx1ugF3kmeghbBUcyVk5XzgZME
z0oelOHPGZ8kSVaQ16Gsqb8HbJ3j9xwmbCJ5l6UQC2mXmnTFCtI+rpy7qRQR
1QcYAWZWSOWIwnvWS5+DMM3fitcWI6M7wWTx/WceygT5NCR6wTgcv00su42l
42neemhmlG+H2/4RFaqcQcoLGXufTdJweKollaBpMSEHbBI6rA3aPXbywHeU
qG8xfgeIs82w5lwAuxcaNR8BffNGHm5TpESmm2UkmKEZSZAe/cpT8d4yykbw
ThuQxNvkkw2tJ67mLIloKai/GvRFMsmqaZKjfM9n4YrT8CTKRUY6KShXqsme
dohScBPk2aC2nUuXSYaO+KI/6Wm+TLPe79aKv+RTugwCrgk7opGcPua8zUHP
kxLiQER6NSrCvMYECgY9qqLAXKzLfPUwm3WXmJV5JnLHsVCNVvdC8dU9JuVx
6LHo3TMHM32sTIJgumjtwcUELc5oSoopQN6czVBxjDNV2Ikn7PKIuIVRw4Wg
aufkB0U+O6xd8cDPG7ox1CMCQM13+6hkGHJahUi8wJRCldpa4vDv9iBazXTM
Lk9eI+FI1pnP7M5CN8aHvR8FXcHTTUQ//cowUK9pnEVaALN1oEDFOs4bdCaR
brQ3S+7fanWO1rnBK06NYd3kzcdw2/mjS3dJmMvXr/0xEld8nCUL+O7Yfdw6
giwmpPktVtLdl/fBLIDqJ7INb6g2TRwFeJYJdPzxAY2hOZxnqiViyHNlU9+f
hOnbE5tCTTC7Y8J6awtDDNjQc7yjIxV2HLw+oIIS1DaVh0p25chLZC0Qz7c1
iSxQXe3a7W2vvjZ/8CLb62q1VrfZU67AuOKCMJtq8MOEpRJH8CaZXaFvXlL9
naM8oRASUWVzdeOedBjAqq93YFKGNUd1VyM4D5/0Vh6V6rOzdj1pmVbmZx4A
nuVrfWAbFZ28A3YJtbPrVwQ8p5THFljRacyEl2rF/g5saLxvDJd5qJ0CBwlp
fkZOlE21+2CLEwJHQX9VGqlH7LDcTXa1C6EprtfTMr364hvb/Elq8eAKJiTp
TElNc7UoTmFScsjZvLCbuQAPbLNpck+p0n5HGdfCeyzIW0XoRn+KCuQexMBl
yzt6JSdrFtA/858uneaMbQ3TzysvDNgbrTKXrGPwzJ+bCexamQOwO4JOPmXm
ZZaEh2Um5BR1SeN4VQ318CN0TdooSOVIfD8RbjuwOyxiVSp6cOtcX4VTidg4
hkATOfLM6tq/YAt0YxykkhwqtVC1cuzKPden1pFOLfteVNJ4zBHX6JOyx2XS
I3V70+lAlDdCeGkjs2evlw3anm5sIt7C4vv+JySsvsQM5ye8b7CDkz8yWtZq
WeZ29Uml1hXW6PjVUM8f2xSSX16cT0g9NnzC2/Gq9/S/ry2cH/MFalHfOIAC
kxwcvGSdAwfRKGMk4kgojCYA8vc8p35QZaevVrrpoNCGcvIKrIdwDvhRZyQS
9eq3J/pMBrpRKr/D9l2Ao6b68vhAZMQmA6J5i0EJDu7hYHMhWA6yoFJ5ybVf
+55wz1Lp3mTS/nZefFcOlffXqnfolcCccfw7Gl88ahc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3GV03+MSyUartPEZ2SuzWQqG/W8KTpN1ZxnnE1u8CcBMPET6V8ny8jo7+An+ODb4evixzfaW9rW88mK/5s/N5Px5qCR6Dz2Bq/0v/UsCZZ//Ekjg1eP11HLySd2BVAL5WmQgJA/q/1hTkZ5xOPeJ29mIROCujseQ3L2MoqCGtBKvrmaNR4KMvw3jvd35nZgOMr6jA+PAXMWY6UCUBNbwKS6ZSCQucRGBiSBDVsf6aXPhWqixdNnXVxmQPbhpxpP6asVHbvOvSdp5ShFNRirYH0QKpru95vtBlUIKS1kKJfdt2pSrqY/ajQrJOBm/o4TsCqt1HT+xWIBguQHDZAGXr0cqAY9oXN1aPTR5+/FRsrpsglYcWS58CVAJz8Y1jIci25McIhtUSEDuKEYDKkrwVZn9BgYBqULH/SMe9juteMac4LrHvISqNYhmI7CR+tH4M2F4dSANspnizkPn6pPkj5uOktD0jmTOrcnrXxL9B5RFbXd0Le0whfVoTNAPvnqmSzf1/lAABQa9pyFdqZ/YU9VuhopfzaIlLv3AagQhy7avsq5aMOUF4UqYPWVWhr/qpSZfAtp7q3Lb69NlZ3WdiC5gspHtm5/hVuwI2mVhpE/hbPOMriLTYUeUaYbGKhA7lCmJI/PzOAeoCUHIEskO7LSrOm8fU2ga5hqz44JUppcIGyKKIgeBtkxJA5hJK7aqWrUiGN3d3PffiDjufcACv1uVwFxLovCXlEQdkM7IDxaZC7zuvWXU6hKXnNuVYxy6cUX4YiSiGNOov2YYcFDLwBo"
`endif