// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fSt4tx0Zgo+FUZfCHaDoszfShJp21s5wRdwWB08WfaEX/7XktZ2b2mrfEv/e
RtMrpimZsN5pxn2v3Ex0hsWkWK32C95ykkMfaw3G2jz0HGg/+b51EZs1GozP
FIXCbeGScBJhw598hY3UqMF0c7937ib7Y6fwPf/l9YCaiMwEsRSsF/es2pex
nK1NPNbYtsI9oEjg6bWxy2H9SZuatK5E/aGoknVaRiB2K7Fw8WtXSeyJGtIW
KeaybPDSxxhk7WTJmB1nTaPj9wfXioG9ITOQJCKAzyR+zlDTWzOP4SzSK1o5
hW7Sf7MbOVts2kQlSW71ZGXMnERpzWFX4tQyftwIGw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kghbSI7orF6EYdqGFdbnyjyQAjLk+vusxxtRklstO0tqAZfoT/MSTx7uAKjR
FemAIfxOCbStow0QQ4L14NV+Y+wJkuVREVb5/h1VUCcztgPq9OV1gKZUK2Uo
3NWbnk5wiqWoBfeDI4U0aqENgnJcl2AysNJR7SwNyXtnPk3e5eWqLtkPUnQ5
vBVtZW5ulbXcrdEOjPiNUGvkX5bOuYJ7yo7KcuX0pZutWc29OqdXAiUHGs+k
2QDNZev+qg8OlZA5Azntt7qCwG9mPujZow98YoIKCcvdEDfcmSRjcRE1leQQ
gvWp3PMzpu5XhOfeR97K6NpVKRxNyM8t06WcpyVFSw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c39c3CklQrpgrPhr/Ua9IboZad665VSmsvHGKDhmyAC91ugKjWYNXU04vvgg
kuyTUY+RklDctMdmrJbYoDIdBK6T/1eVwtvm8lxcqel3gCXuF1CH0h8BZoTb
7odHs2ErReYRbCTWxqndVwvEybGyBBcVWlDSu7z0Kw8p2RH7GL81tE37YI20
AUoY1vqIpM7cqhtxY7/vx8MwLVRIZ1oaFe49OWDtsAEGo9irx6EloCb2dZ0L
I69A8hURQastaB9bz+ZcBW7CFRvHVXgDr0zdnx/pPB4gjsfXW1RrJff5CJbd
ax8PLLBcu9UqQ8rzZWw7bVVJPKA6JGjSje0cZJeCCw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Hc0jiT5ieolH8FgqcpXgOV6DCnQrO1tr10CW0+ouo7abWuOp7q13nptvee+S
1KMbqFDlIr2WilB8TsAU6woD6LWFvV8XMu/tcWikSo1yKGjbfaEXOo2GH79H
Acl6jg7U3h2ldOw4itKuTVm2cWGEHUGcd5sNyCLZI458L7PmP4k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qsL8HPtFl7qFxNPY5Lz57SoodFNuucnJ4VDEwxALn2VI2RLwrVa8DTwPSJVX
4Ii49tL2++GljoU1ncTlM5J6rLvWIXHBFc/WK7lU3LWQwqhV6gdFK/OBOief
qM/iXYfDvZugrtAjxCqoE/ipN6KmT4Fo7d88aWfKr00A5FVJH0HDa+NrYSlS
0R6x6MobD7wHRCYzxHlEv4XLKvfljVRHTXFDmNnQ0FNF/jyiiEkqBOOwha4F
mUGOJPCWk3rL+l9Ug06NChuenY4summASgkhq/tl1gsnO8kncpguckPGfrbc
Bv5GEYQYndWXlLcu+rAcilTyCLM75KBvxIaC4LzQbPqPxXAHIMcgHbv1xW6j
nVjRjK+zFIYLwpfZqcSBdIZ6IGaX7FF9bUZ+XPL5+LOHn2EuZY7zK31B38DT
AOZeYsEyM/dbWAbH/LW4SHQbF21/xufeZSvdRNyd+kBLeB6dzXF3GEA2XyBy
SueWUeQceIhKhuheFpSBener+ckKQP6+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RMYlJy27Q5omXWXEHRBxLts+wwk1rHPYRFSY56Mpq2+nl0038F2zvUJCKFBG
OLI7F7FLCCR676SLABWuO2yTd16nRQIjJI5egbFK38jWLOmCvEFC9tN2DhUR
JgDXOdEOLQNPNr5Kp6v7vNqOVbVVR5sJiqDp1TqKdC1DCjk8Hec=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pJW+dsBuR5B8dsGZZtAxFDhecmY0Grw+fFh6sW1RMGHqEhdj7ER/aVf+dkkt
3qvOd0l2EaKnFqpgWBMlYyz2R0lxq25WI6XfIHpQMG7JuKYSl2+D4x7Hh3l0
LB6MAn7xI9uqx5Fbqn2Sh6Clfe12Lf7ZhVai4YoYpueQyCIPrGg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46368)
`pragma protect data_block
uK/iz0gCKlzoUa+XUDPE2ZYhO7i/v9RQW0yNQ9vV0xflQDR4FqMd1MmHd0sR
Ub3w/4SJUluz2IBigEFBrnOtXjp2VUX1aXYu7BuyHSzmO+K4Czv8PxOKELUX
d/EK5IfeRNgo/U2bmuxx77r+sh92N+OiYpkuuWtyNqBTFEt9aPYdK+uuHKta
ShiEVGpqlPQA5pFK2r9XKzF57WdzVDrRQJg/TW/h+r5XN8Szp/NhWTt9xGBZ
g9oJuj7Es2KAWvNJgSiHTr+zy+GVLIzYnXa4xd3wyrMDTdqSLI2XM7hACweP
Vs75jARU9P+ZFVR6lKwqJ86dWqOTGXhO7YxALxrLqvGVIpZD5oUVR+N9WmIA
fRRbA/OUJGCpPqnsnTeKxIYpE9QsSj/eXZxKiFJykXKb4r/j+9uTXG/oXhPC
gDfoAKIaRA5l1Mjn66LQvT2u80wT6VW157E4CuMdeQjMI562t6/3GfFPORqB
e7Repw1iFs/N4t29N9v+scw/Heqe7Nsr/5AbcoqduiPxmKqXc77qcSqNhsmP
HHOfATbeUj2PZIVDUKTkbls/h71/wpEVxVONOs5Ea6p2RGGifSyTBzQGpfs6
R6GZmQcvyhxnqkpgJE0qlwiY9Ou1GWNNCzIFNceL6RyrSWjyL7OV4rXJrTFW
Js05QCyao82JCDn/TQAZ/nkC007ffNBsk+x5I1Ci7NpVmuQVv0b5YBpegUKi
2VWdkKC7ybIKelF9vYQHNeMNbXWtXWi0S1cbxQYNoMycJWaVNYR1Wobp3K2d
6bfV627KZXkgapnGwLNQvjhnAMWIko2iqK8iw6ZWvy6KYy0OUwkR775mxgT2
s46yf7XyMvCpZvbGxvfiOtNCfV2PnDethAT+kYsahnuPmEeyTAom+0fSNJt3
Eh1koJylBoecq7UmH/b6eELnRbT/RY+rVMvZkIWkafXuckCT+xxZGY7b4/BF
w1lj/XoTvWwRfpJ++fW8aRz1AvVrj197JnsRxJLh+sB1gVy7R/Bf779OllOH
kSl/h7BWksHIRmfqst7LYzgtZm7xc8Rl9OCN8hH6oxk/o9iPITfka2+UEUHs
HEBH1VB66sCl9DAN/EKqw5cz0wLavcMrANBXbEgLk62gJDcRYaZ5n9DPaUd7
IGA++ZCxysdgRVhEK5VFaew9O90ZZ/v6j6tjn4h5tCW4CM9lvUV9BX7EEa3S
/nSrDJUWddNjUa4bjmFa+kGpEMl2yy1Gv4nvvqx/M8kINJWWUQPX8bZ85qQ7
lLLAUivGVKlOev4qrok5tMS5hYUdQna++Eutuq2oD4q8kz4HkFUvyTTWRjkm
LxNsRuDpCA1oIUcOlSX8feR6aP/GdosNBNuuXsWwjvrZH9ejzRp4EjRm28/O
Jz45hCePwYRayB6mBdg6W9lXraiIy4NP2wegK+NzSbEXwGR3eSlQ7O94B3MB
3oXmtbGF4SiVn0CEsg/L7Quvrvmeb1J60e0boGNS1LQEJVjnK0FJhH+rm3Qd
cmUtxqihyF1bDoo4yBPHlO8dPXiKWZLVn/H0FCQU8na/YxUranYISIMlLBUY
cXgJ28FVsS76Hgx+W6DQKGAIyW9GjtjXeUTZOqnhozS1EQUTJLdZqMhn8q+2
7rbZQzdwVLDlXgsNWZyu0oJboxIouMtY7DkKM/+Jyf1IfmIWZY/HZbaMFaZj
ZlU0jP481nM7vSLzaRPk+YOPD9k6+VdMYHz3VsN/xP/ZUnG3SIibpxqPINUD
8vFYrN0Ki5GbCu7rESkhNPkqfkWUf30905rra2//dNAgnzpe0BmJ87BdgHkI
qefMIuS3HO/aQqs3/vji1juIRHDXx5Iw10rl/oc7bV2pVTi1BCz2n+xhDcd9
7BlBW/1+OxsNJBgLdQP2E7oQRtniGSrwSx1jK7lpkkt1YSO5nCpIzK7lLryW
op5nTkXj3ykXt8iBhK0B9fs8cMKXW9IW2koyYltQPZnH6PYMT0N+dEnJhsZw
w5IXvaMIJUmDewRTJaCkOHkpoLaQVnwh6C69FZkrKqFnc8cVlN8oLNDNs9z+
snM4cpxVYTOurXCjA4u/HMc9S9x3FRRVkNLbdh6ySR+ZQCx9xhRGBW34Tb4u
84jf/gS18GMlPXD5FHDnM/rSriF0dLH1ytKspcludTzEu2Vsbw7/vCOxV1b6
s9f8ljmLLHMvi//aJ1JEzPmEArF9zBHODtGFZh/IQMI+G1A2TMAUr+/5e+Dy
ULzrwk8L2/hafg83wOvlcW/7W4yrzxcOAESlXqfKCLrnRbF/KZK9xwqKhmbG
BQLXcKNl7NB5ngCYYoBHB3lSs+lcFdsCSMyG6MBoRHGPHAwfUarf2iSODEbM
EifLIeicrz48RYDNO2QuKL/BB5sBSOMaGkDfcLXc6iqmsST5+dAI8myXNQCX
cFu/+wCoQ6L7I3jMbhnjJuedODzojnDROAhxTWcSPI2GUBA16TR/PFd/MKXy
oToqpnpUnEvT+0qIW+Rkr/LCtl4CFgHAKn14lwXKjxtiVdR+6gJQuEoSMPUt
4yTeRktWdmBXHYsZrsycDmXgzc3p6DGZ7t8Ga/Gwk6698W8LuPPSdaypH5/l
90Wn4KHy70BHlqBev1lVwJy5eWOVqWgQAAMRa/yiixtkWMhfr/owUVRKmQTg
byY81a3naJMX42zVaxEVCnj6/UgVVQo+Bm3G1+zPl7GLYNLM1qlQZDLUGzIe
5V5MeNlSD9EZIMxS/un/V4CeDxDvMF5DLcp8deLVaeSsIicDrKuFxb1LkSCa
9lV6gMrKkLTFQIc3ycWlirS5YcHRs8MNMfiPAOAQdNqpYNjkPKHULKVl/5n6
X/PCgIm9dfQdgxYVZuQKbzyLcmh6RbuVauMa8v3X5AZ+JB8tAqSKZJ13ZtAp
kHGH91aoTWsmGwlDbSyo3P0mshUoj27Vq8fAGqnHg6wecHTdJ0pBbAearJcs
UCUjJYxDgMJnS9PG27E0XBOiDOyMC6ecLCWUmR7QeGkYhfcK+imqKpUZA9bk
VnZEvUZLwt/WLa6Lk2JvocqfI5KnGVEimhacgbMHKVw8RkkOJ/J83wsb6WA5
ikvOHlzTrbG59/CQDuz0bwPoe0WmOphYscMcoqH6iS80RgvEWdFDDA8nGPXZ
uJmm96C/ipOpR/5xOxMKacveMw71qmeBmO3ZzruVI7mBpCzAXFCvIWmOxs+U
dJ01EBQ7/6RZnRRgQ+dxtsm5F0XCzWmYpS1YU15qBX1f9trThjq3YlypWerJ
QkS8f3cNjzquUq4iXNqkwZgE2QSk1CzaE420apEwt7shMR9Ae4dZjIgWHHCl
leM7pgYZUfr2Z8iRh9M4UE+VAkUmAvHi1+4kDMHb5hTFjDLk4t+ZihuWXGAj
Sf+p4+wkas/yl9EXUFcTbN2NHga8qHksHjvOuPwZxwRwdl+qx8FFXRPK+36d
l6Q/FFXEKOj5Tdn5DCeXE8Ik4tcQxtmnVYf5KFcmmlXyB+O5Fwt0/iO5q9/Q
nyLIfgOLbFRyOsnrWqLIK16yD+NJdIHiKrwtdZx6G6AieLTdWt9eUgkOgWrg
TmqqNIsw28XJPAQQCkCz9005wmyvFDRkJRIVH3w5eIPQm6037Nazxs6BoCe+
2ygJ2AqYuePGiX7QSMAcRBe7/bNtKtdPqq2mhmG3KzzNYfpoCToo1FdhSyJB
RjevfiKoL/Kje6c8JBA/1W9NEZKwa2LtRtx/Q89Uff7AbgFejcNHnFD1603T
npWVxyUmLIHdz2IIsqj5L/0xhycQ6YTP1g9opSF3Orr6RqAmtIHyNYMop1YJ
k445iUP45TOaTFsVM3K7ev3ejxDof2fWc1+tyUEYaCb2oJJ3QbTH4iireuDm
yIHVmwZPy5kkQpl/vMccR9ncQJb4bNkl9qPQgs755euwHs/B8DlKnyn9fW9B
+KaXIeSxXp3D6k4vicgzoZb+mU1pW8r1hvr1HbneNNCNeykZyrHDoMXsSuXQ
KBKQKroQ1uEFza0dumkiN8L9fTTm8GKBcIywdmXJ5ZznbUySIXFPyJVLqLmB
l3B+FoR/YmiqdGx/SVkS8qVrZ8IhsI3NKnDl5uKt56vNcoS5sA0CMCMLVhgx
x7+VwdWeIbO+FRwqWXV7f90MPW4UpQCVAjWKtUrB43SeuIikIqmUiI/7s7lz
v/dHfwiKHpLsY1GBlTLM/AqqqPOBykECYYPBCEZI5VVoWq9x21PukNdUx7qV
IgDH05gpPz2/CTEOAAICLRDaYdrfIiK9Tz2qooYBzElQT5z9Q4ZCfvYbWz6o
kmkqNY1pOO24dfMrOQnDnS1gKokK2NdotXVxcUBJ7dud7RUDCasZn/Pex/6v
DMWrp/rADUj6GjppDWYADOeFkusW6MGsES+PfumI+9aMWqHE5HG8iIeA5nuX
YB+AEI24CEun95gcHT6aY9aWfxGh2CCizWKZ/wEn7Nf50uYbsI8u/Ku+jEIA
hOOKxzQ7ehw4zKY3uAG6kD33cDUP5C/3KjlEmuh2IHI+3GGrYaJZe9vOFkKm
ldq4TvCi/pJrf3srnfuLuzKKCLlyR2vRS4ZlR/pBcb8Ca22AZ3fx0x9pilHM
01QCAuOwHzeFPAw4v90kRyZt3VPr/oJPZgF8EoxY8yWLsNEUlT8+TILQdLoL
1Wn4KphXLA6mYZwlNhCEtnK7QZ6wXDkfYvqeKk9mMkVRDby99FThKDOMKrX4
B0HdcO22GGj1efJcfP0oMBC57aio5iFSqy6x/JFlDFEFXAnbbHN5RTXDj8O9
QA2J6FtXykaC+zs+QNAmOQ3aT9EskODohH4bj8aoO6w+ji18lAFQshAC3384
3v2+TGy9A1AhX8xDllYCK493iQIOXLAlOMZZPoYUT/dS1l7kKDGURPlgMZJ7
ZCuh4J2zFtnJ32EWHpcUM9L60gduYVq36Itjp7aJ0KHpxT1/9SJlJxnuJK1T
5cNKoah4Y9FaoBHXPdB9mHJKTy9qd3IJuZsWkNly018rNC6FGXyGWaAmkKIk
di4RFgXGheERcsqNZHQWLysU0MrtYn/bsd+BTb3X6vKPj7OcHVJQKdML1/O8
Gqm+medYp6UMd1Hhzg1SwHGcZ/4+4xcslilp/VOIoqf3gz+ZGcbcehZ+eKQ2
VEGIf8nkK0QKW5Vmwieog4gDS8F7BZGDWfvHtKNVhL1wMuZ/QlyDUy3peAUS
4jqAGe03ZiWmi9ZLhPUUHzZOC+kYrFMgXZPnfkX9V1VrQdva4wz3Gnt+90cK
KwUqZbvc04T9aZvx6P3Xdht9O8sNTZPI5lKSDZrlSSJEvF7Ou8JqdsU++Dht
NFh5eQEb7SomxlSBdb6t4DntcSPufsHDNKEat6ch/bsJFhGm5UZ1Evv4zFJi
VGr86nz2nmMhWap4aDTlvE1U/y887Q6JPGRzeWQJMOg3aZzhXTTBdplbwxp9
V320Zrn1O7RNi5FRL4aE8Jfj5fd0IJ9mFyPE0c7wOBNANfjHDTfhfrXoPLIY
7/o/CSpAKmi/6OpzfGvIdcoBHGP0RrnNK3+GpiuVyO96fVcIYs8XokLsRpBA
vkKgT+W25B9fAh3iAOBo4citcNB8AhtW8aQhPqBcOF6k23bUHq90SMvCSSCI
b4pXcC7kntn35ja23TIbhAe0yzAcy35uRQmZXO2KuFFmW6DY3Amw99smwKOe
EiOJZgjsdhe9HWd311Xkcng/b9r4Nv783lO6Djmvipps1rObCp87fUnsXzPL
AINQmpOOy45QJFsOqaicB8O1NgVdzaY6ZZaXDnQM5MtWnEmTSOmpSpPX3SuL
m0nV25DR3Qxpo8uaJdf5tzz9WHWhOrh3TdJKWr3tsXAiY/20wueWGBNpafHf
tg3zmB7Sgeij/PZiiqoz3pml3r6Z43anqa15k11ZbbvL0CQAAHO8gOhMHKvH
glKScYKX9xvbWsRx6SXQWsijfXYAlhVSsf3RrLXh7q+VWIx5LxH5ZnsAszRE
cT+BmgzbFVE/+pSDRHZKP9tz64aWBi0kwwZKcV3wRNWW8H736krsoFbykSGa
faORfaAXVNc4KknEkaA9Z8C3V69hRONCpKDNr1qfVnveW6yFOq/Qso1qkVK0
qxnqlLWQ0iVOJQsJp5yxuY2qEti9aW+uXaOs4P7IifCwdsukfip3MHdLI+8R
cwSic3t9po6psEoxjOljbSKKohISSaIVK5LKi3oSm1mXKoOZIcGHke9VaUs/
yZmkbgw9kLPMCtMouG93ajqDcGQw8VKcUaa12//8K+s5iHL5irulkG4zyZSZ
gF64WB5jJXoGd3LB+oNNE6IJD6IB/XMKzf16TIUcijgK7QpjaH8iox5n0+82
RbajyWq1IW8YR5mk8/zLEWPgjeBVrx8KrFD0VYKnadlmZVKUYy9ugH39hHaZ
hO3+hjjXRBWtGVNR+3xLeTHsq7exi1PSmnLktWdpKgSDlqk+hoCYfhNefzkq
iOqc8R3fWqieqMl+DwBgKa91JySrxu8z3CV6tAwsHD6RvH1OZ7pzQDfOpzHr
a1zbWEFj86baBEmeeiOWE5P6KKJz0tONsUrLrL4PZaNfGJSmLoiiIycB/L0i
HVkThVzp3bzatyv9sKGR7jec78/hkTewba30q4WKrqcfLKdCYYmlHEp+Oqz2
nKceLsjhPJe+OTXvEdw06JzfdQgb9HigWydL7HsKqfKM2XSiWzdCFDS/a4GH
5uzMtNGg79ui1q3AA/3AHRX4WvPtzotyOm9eQqNIykBGq2dWOp6+3P4/KSNu
2JiV8BBjZUc+RlRp5Ry2JLDJDZKWEltNypRKbNF8uQ5YcaLEoR4BaoSJcxKe
9v6gK1fndz6IgDf38/JS5Fe66szgWtK8kk5wNOWD5WCp+hQPMfZBej05gpdK
H681PKs7Iz7EoPeTPairU1d/UIPRT2zYsWNTkF/MxzMSB53TNbgB3fkOiygh
mqvJmpfgJigNkZZqmMyEUz3bJ/FjeLZxx5Mn0m56eqKLLg8Q/CmK24lh1DYA
NFdE8uYPFGGqw25DEgWxvo6NMZLNeuqObijPKD8A7bjtICwfxzVwJI39cXz/
IISHfjR81bansDBt+0fmVJEHu9ODo5WQApQCJgFJWFo41lfc6wEqy7OHW0KM
NvlqB4RBS+ge5JOXb1kWcatt18U6mQMoNb+tMWsVPlutdoTkHq/DOy84bWlg
J1oVcY0PN6I1wiUfmJHHSzHPrVIlLjCu1wIqHyQH9yUnEcsgbCA0Cmz6UI1E
RlWRMjOzvqrNEMbmOyAmBtHcVj/IIQN7XKbZNAdDclNAymOV9ZI/SvAMvWZx
gQPZfhK6ZSzvX3lkMscHa5iVijPnhoRQjw9e1rWs75vsW8CEbnyIzcwBku3P
TzKSxk5rOGFSzqeOiSQbUlO4uC+2b3KKPVVf6hpXv0gwmeFVb7eRiZyW18nO
ZJw/J3uIMVDM/eWGRCdHvVT7CZ80VufPseF1KMyJaGxcpGMpa/N8ZxUxm+oX
vGrHu88R1NEJZszA8DF4Ng+G5Yjt0dYCWE3H6LhGcHGTDwTfU6PAsWiB+qcJ
nmA8cdztjjHJpsZcREi03gr34UELIABzpIbWh/vtrFQypHjHpb2/WPr6+zdy
f5QCR81JOtiUGUlrSfLSqtkD1BhQW8fPwbQa1YK2RqI7qoVV80oA0Vd8QYZt
D4yjMPa/htMp130jGvPOff0+aWWHvnfH2/ZLoj8M9LSfNLpsfK+2JyhyMr3d
OlCiC/pcoecSFFRJI+/5brSyP/Vl2h0H4wYRahb39XPyd8MLERhHfON/xiPb
NPY73p24/cFw1qfcbOMB8qQ8KTjWu/IbjEBJaOmEyELq9SGbY+AoWNl4LXJn
Wpmyea1yzpoFlDwJDUmVt48/MdN4Tn1Ny7L7kmOttuXLFWHGnpCoUtFQFWjH
qKl7KGN050jGycXT/dFvRqmho0oqeOpUZH7MjKxt35xtECDtbROTpMe/70VH
fTXU9g4i3adoJPTOTSpEFEmui++i4bwEHTlptFWsnhQOnn9S36NjFpJEGAs4
E1x/8BWcsRLYOoa5eIF4a124CC2JGpHQDbvQrelIVDIFr23o7RBxfiO3SjW5
oaXKku7Jai9zrrsZizfv8q5V39AxdriBevhrDRZ4fNlJg0FSlCbXTZ/qIE1e
Utr9dhqoAUGufuhoYi/xroo8LupDE9eRYHgRulGWFWAiZdwhgCs8+Haxemwz
slED0lriPPN9+uDKO2mKcoQok91z7GyvpBozLI/FlydxbTeGknzr5CmjGYrX
4KbW3jXpVjJZys88R3P8D5mqewXdXBaQR8eG+Yg+mvnSwa1EDHtiF0yfT8e/
2OXxShnOIOQ4gkGKQNmYtR2Cu2zAD4ris5JUFlv8gHOSmLHfPBmkrRtvzEr/
v4LfhZLvsM+PjkzRA1x8FD0j1Wl+MXroyjZ0ochmxhLPM53AY+iAtkT2DJ/h
o9G9omFFrMf9KwK5CigubyUoyuAXV3/a4vfMbawlH+VD+dCFbCA8XKvAl9X2
Ky0dgm/JGMVXqzul4oP6sidHBUyBv8LVb/H6HF+qE3OpYsE3rz4xqcRUzMdw
s59MlI/nPR37351N7y6o7wPbeF4tqs9y2UbL9Df6FY7tImA9u9gQEpnGwyFV
UFxOQAKm3PcrTdoPES3Pb7yed/n6uxWsPHjl6rQdWoPvSWoIKCCRfViiOiqp
3C1SUiSQWipIszBfataOHt4eYJt0prPbGBFHwp68vnYLsXs0//2TOxHMU5WL
Tctj3K9RpEyJ/ehY+Jhk4RZ+/jI7046OeaARHwCnlkwSyHCZhgOGhC1GtgEq
yspngjrcBYeuWAQxvlhzyg4OU+FCsAk2Zr4S+scS5kHeUQO9BQxysD7bMFHD
2gbNZ4bfIAh2OTXzhavMXM9aEzP56EY1wu6H0N0Xwp2zSIj9wN4kOxp8B65F
hRp/FXN400ZcSEmNjIvv7REZdrmH1pwLx2xTDAfcMux+gYx6DARh23w3ALfW
6x4Q6aqHYBh7WATJ8lRYsjt7S7PPXvdaNY/R50EQ9th3O7QPUUgsCFXaai03
gZ625UNDzy90wTCJX6BpoF9K069AuPBwAW/gXOviW1xB8u8snU2enGm8hH+d
vUvLjpDUj432PjObOMYIGgJXe5+LWFANR2Rgc+yH3euh/hZkPy+FiFYrxKsY
itjpyAvKyFCdIDXy0Vz/KsLfTp8rVUSNotT+/QEc0RH+lwi+mvbs+FOf0a/D
u1hnOaXUlmSi7xq5Ic3Qt1BHzn8PiOPmpR6+6kTjizEQDibRFH2q22Wkf5hc
xQHOnlKhD7BfJ7DoUNSGqlIZY3IxY6ZtPMJ+J/4WemMQqtNH8JPS3nb87yNa
PGShmujIMvgEk2BS/DNI66Cvgj9Q6aEVFPh4AIKdKkZjTiN3d43MGloLjvgX
IVaYIkH2WPZh84EXVTHLpvqbXXqA1oeB3a22pAASou2dyZgDrgrMXIUn2nMQ
KVGgFvC/HV+PdNj3/m2Gv6H0IQFF5PlFBlNxHJ35C/P5oquAdcxsLx5nIm20
N+ZAkbKysZtIPs2TIgSOI8+Y1vg4/vx2atCp2qgNgD8b9wHav8TZPuSlRODo
FGq+ui4qrxEvukch2g3lwBLD3hT8d0AQ7qbT2MaAREOZbVTUCcAZY8v0pBzO
2aMuyKq8AG1qotVHTjubd4mVeHSTwrttGCWJVYxU2PsweaK+/FV0C0DsJEm8
jGkoQzIuLv+0s8GdT2zB312t3O14CAYT/iYS32sPzfz7OJ3m8gh7tOyFPenw
/KRMLfP7ao7lasiVx2eLLBeJB4Y0LwrlmjcOAw3/30r0Tqw86xop5Dt1BK5O
TgTiJRFigpDdmDQLmzv2npl5O1+5LJgkcAsQ5BcbKWQq3sqXclzlvDxGkNkd
NXlnlJyFcpWb3jBkQ2cCGKH/vBQuY+/DRo6EWiEOntMdJHehy1qtDdOq7HMq
j9k/nN68MCvDURDyJOOegm+MD3IlzqGjLo58P+Rkche0nX/e+Fg7KrOwITcd
GvKV/qWxOU6QoVjXHQOMJ75wdHRieTiP1vbnXOe3nyDLIvMlXdQKKcQ0/VvY
VKjUPHuuv+qtez0vteNMzQQ+vKHiEZnit2Cwf07zBVvIiS9FDjnVgTTVoa44
BCtnAJjwfR0UQgREWio+49GWbnHPI/TQQGh3JWop7jQJJ3/Pky3raXw3gA3X
EkybqmntnyVyiRbfhO4D3PeubYrSh9YClkEbkV+nb4CHI65/h9VKvp47M06t
5tZZYKBgdafe+hfbeZXPZ2l0DrhXYXiSAwh/7Ladgrqc1sdDvOfa7xZc6DuG
UIGKAyimgj11RiR2X3E/rQciGvdcsbtn2hT/65zgMFTvtGChLlDlXliTqY2v
E8JIYrwyUlv7888Rs+AyB3EvqTz+qA+EWMGdcy0xz+A2qk5M+Fhnv/HEMFCQ
ov5JNBKylnIv4AqqhHa29LkDvtSw86P8X/FVqVRuIK4Eu2ZvXtVOGbETn1G6
2OcFBGd8VW18pfqCQl8fQro0FNN111SQjNS2xSjED0FJ3B0vvfTnWMyqPQgC
DMMVW+IDBUNCn5kgqkiuHkLKd+Gk3fMBvH8MfmuCp4KPtxFYeHWXnvqc3+oM
LTcpk1GQ0IMyYKMqfuoYesB3JP9F1HcwbWx4C+ITMhcR8HcWMSnqm0ksscQK
LeXMShV7scmKSDn+i5JAjQXFXpPdlrWBlJkF5gZf6E20uy1cjcmJDtB8r/9S
3TtKf2KPi5OjtcWfKzOGFsdlk0uMfl098mn3ssVfV+gwKxGTQRc09ihaNWhy
NaJ+0EqEtPpml8gWJ65/qM/DfmsSkaJCMXvDK2tlz6TCYwIsqmMP/beDJZ6+
0HDL5mz89o678R42rnfPF5yeyly0H5j5GO/KfSyAVwgwijctb5eqH1vASZRB
/AsJq6MQqlW8zyUl/TD8PFT5+4XFaS7Lax9JGJouUNxbnYkd7D6mrsqSPCXI
O7XIjLut5pmcO6Rzk7qFu6vhPYR+ldTrnnmLKmgf5qeQOgojwCuzQMARyJ15
50lyOBMAfPZxSTjyzryJspoeIEcMQwdktXk4FzDbbyypAg4VgWpctnb6TJMk
aLwkPDCPhrXJRq6YidDnC9is3IKw7bUWfs2Dkv+OXZ+3UIWiLmFYgqzsti07
83EWF5JENE2QR/tIV2Tr4NOb+Hb4+8p07nAdfMv5ofTTuwECo1hLXfvni/pG
EVHFlgpI5T7lLynEP2XxNvNtp/l6SlFLuZQdIiHLZjf+oDywcCIonqSGwX16
qcTINDGZ2+q8+PYeGU4JiuCEE5qk5uO6RXaBfxrxttgNo+maJRR9t+3BB1WD
sMHyp3EeqCIincHjMWnL7SrSSGt1TkLBmJ/621SloWafkp6PQZGoIN5LrsHf
N3F8f3ZP/i6bsE87JUrYR2NyBTEBhZhiUxgIAX29wjD7P1/d4x++hptbUhFo
abW7eoJFfg2N9YytcWxJAM9x2XYxX/h1UlF6S4FXen8IYruKxgriKKsFji5Q
boGV4BLK8xLv7GUr+F0IYTsCPk4j+OMWUscGaRcTRP0V8Oaz4hGdsW9Wr/i6
JRorlh6xT4cW+k6bpHClZmDJkvWkulx9+IBo9Ei2OexqJrfuYd3kvTXOKEiz
0Lnphd7sbmVgZWH1s0HO3M+Z575D5zShbSNfq0CySknMmRgV9FsuFSJ53s8N
Jdv8/zIDdLiDbVYgNL6s3uP/XmlunPwJUkgkv5636R56q+uL10YHXCBr57mM
a8rUts8ZwHbjfGD//45+FQNF6yuArZYzYFXEvsVAZUbNIBsaHNFANRa0Be9+
EY3cXiscSxFMFOlZAvOEmLCzWLIVw+ZGBIkPokRR/u2VzesEJakoPlKs6PBg
9Iji2+CdWDpMJ78zSIDbm+C2xO+Jz7lghG2JFDNqeMS5deJOt3KBuqq9PJEP
LBTKo5KLLQbDjiJP9oSK373ZW3IkJhICje8yEIGKEq0k/Rgaml5c2jA8Arv4
NsWpLYZYhDQnryfQ8B6u5/i+BFbOFNaEpdxFcjMGNR+tssCl+eT29UxuS4Tc
vnYnpkKqZk1hK7Tc3so2DLiVXqun3evmRVktBwJN2jaaYHjcVpTqn2/A0lIa
rhdm67J/L0rPzI947F9zKvIeaWT7t4INgDMEQTgW5daXVjlbo2pqJzPUsGjV
u+T7WnQOcGQn56aJybtgAeLUMAMctSeCYE0rnboRcvr3qFV3cEg0RCQ95Qc7
zfWWU2XqLBPvjVJFju48y8fSMM0syFLyx7Nv1gejI30E1wcO2v7ssPMjr3/6
P6qhIK66PSUDRPS7uLMsNdISRvqBfTrz7q49od5QHOYT2fzpW4KkaXU1ng43
hMQWh3xa7mujGhrjYK+iOkVZB07z2Isj4yHW9MrWaBAE3Cad1XIZmKxeEK6b
hb9ha5TIWwQumV2kH9mHqk5/4cTN212uVm92tRF1sFsCfNHl1j5WUc9STEfl
5yY02kAafKn3PhlpNMEvx4uDlYP7w+MB76k5hxLNZV1otfXrpjbSMUvCkJg9
+hwhq+Njveye+zHrcc6NcmUl2gfWWDfKLYPrLNbTdms+sjFuvWi9uY+oY1CQ
prB8LrqrYYHVHiYPOwKkd+J34ifOD6MAYoTX3MSHJqBEpVJorhbG1s7wd03g
b7+JAcCtM23OW4KkzME21FXEqddPzgAvQ57fQNkzu+29z9/vRr9WMbMRllpl
SUcF37gGvW4Ja2wrZhQcUZGE8n2Oa96k7nP2KK40Scy9L1A7FGuq4JWQrpL/
YOYdYkAiPc0l8qVgdGMgdIJ/OH9Jr0LhJvtNvdlVRtbGqnQZjyTHl26SW9Wd
IhBJWmA/M546ed9ysuUQR3cFQ6OmwHj6PygmlbpY+Aq3M8bO2sDYkkim7tw9
Omt93fCtz3/vHQp03D1xxKyMXHTJ7Jor55Bmh9Nv5BhzX69jrGkQvuSKCk5P
gYzqdMiiwC5dghkRuDbfWjWR7Puk9fl5hDNYcVEfXGqlpZH+X6nYLwOQHjJX
BGQP4igDPMknQ9HBZRv3PEVpTDq/TfBbiltQYbjpSTTZHGYrkt4272NvQZU1
lOwMo8/7SsjmPwbWjky8MQwfENQBVYrGKEwb6hbUl7vGHkJzVliC4853SFoz
kNHFCuvQ+8Eay6x3pBXaPm/mvlxqGzNbV89XJW0qbJHysJWA6CeCdtt9wR8j
S81pNN7S5I94ZAWKXYE0WtJ2K67xkhJ5GHjojBPUhxSgaHdBk5ctlDHTH5cn
3Lv3ezjEbUj8cTCdGUbs5B7FbMqjOTeg2JsDb4XFyJvMe/4TdbplmKtDBDlv
84W3aTILo7NcG9bjluP0SpeWN71OhZtDfD9kH/HXRUC+LprNX55Ec5HvSw/q
+CsswR/mRyh0q/OMCtAD3RFMHtil72ptK0vwmpWxqn/ezq+BaCVfZkQmmzDS
g1PV5wZX+/bRgYYA94vedMu8xPGVHzZsK9s4Y7z89SVcwKwknQssh5+e/Ap2
u5RrpVB8JFdiMB6VYdZHE0BrWlVviX1DTo1bYauy94r1v3sv72Uqt3A4ha+G
IEGnLV4254V/SYxewoqh8SIfzyeoeNJVIEPCe3KgA73kWqBdEtcJWwDpViqj
rwGVv5Ned+dA0+UjMByk44MIkCZUQGFcVEK3b3y7mirtZsLUvFmOm5qgCsdm
gTTZ6tKL8O5acRqE+sNitBeLd0ArbOzpJZqU+wT5+UFzlTxo48iRaoh7NlxH
pMDEeQRRvAvP1Gz41acM83Z3qQpV6yyYUFvcVioNFePIK4+ZhlR/R5v74t9p
Sru0hTWt9WLEfscdrmcs7KJK5KTlFLCx6oYfwzeW0HCRF9TTLAyY3n+riypJ
t1o85q8DIO8ZGtdMtbGhQzEVfmiuu5SLY/Dm+vnqi8oR2GCJufiZTVU8MOyE
ZkMiKPgEsxS1kn4UEzRMsPWlx4LekTUf9wd2lXquWs+t8eBOWX+wMLtiniAL
lF9TthH9kmgbEJUmXzBH7f0pBmQlW3tafU1Fy7QKcNxO2PEAF3BtHkPc9/9K
LkLGmhEzt4BH++mJugDUgjCbMosp4HasyoGMc0YksmC/vtn7Ls60iRSr6xBP
ByObiTYTFHaWZNC/h43kUYxThKVI/CqK4SAyr3epF3LdDivAahbcHrzH4vQq
CgQD7uuXRMSUarMX/o/yHOMJORKOiV85nQ/7bTclVQT1FNtLCWVTyV2dYPuJ
g3Y4ohZI5V5XXEUOM37hlHtZiLY300Z1gr85FcHUFVLVBvHfC+86AXTlTk9Y
w0wl724P+qhNZ8UWNNWFNtJV30BjjRk9aHn/mgWwN8KdVDqn2DR2blHJMo6I
IE6LBAZLNOh74HIseC2KRSspKOLMzIItMuZDXVMeRAb3s4NdaOR0z50CrKuT
vDxXkauwaS3pYYm0ApFzYsGligmeUnq58KCXmxaduBYyn4LzLFsKY0hBB05J
LkzcFiP6AIMRn1A4PoA9ZolPPdy17djJC3sk5WXID0BJTOK6rfHYVq6cX9M2
Nw+pOW9NhliuIBsuzLwiom8V2cVmJy3aox97ZzwJvHFHWg7y5dh23Hk78P+p
OD9Sp4tfTiUSRNn1UhGmexZedP4YLrKVWgg/uz931ba+TEIjZmpr8wSvF7Kx
AL3NOFxHLuYac5Xxzr9Wob24by0Dl6gtYLatrngwkERFn9Fq8q82NFc6tgBI
w8IOTUHWxg0OnqdvpfB47MKJQnFJA702Aiiz4w4eznq7Q5WhzkUPXqR2dWvs
IK2OJykR9kvwfjWgXOFqeArbMiD2CotmRbt9LAXzlqfLnaNtXanVcEu7Ujjc
KHxDCxlIPerhkjNv1VyfeAy17RDZWfOyrzkWouaodSr3Xr0iaVb/LMVX4DYX
HE81Tm8o6vdDx+NrwYGEK87MXhMTM97iyrc5Cx24fb2UkMNVwhmoq1siuS1P
parqjxrkvUkv7OWnndTRDw6yo+FW18bd6rW0Hm6UZiK5WXEP8wQMOPvbs1Ia
VVevvmv+jrHldiKp+pJEat3d5FkWoF7AK+D0IJNn7wWlNcfZdmW+muL31Y6/
ywn/iulJg1gJ4ICy5LjppowEOLTEon+dhtSQKa/cmVYQxlk4F9WYq/Rqs8p4
KFX+tpBe/m1zwY5ICKJZWiQ1d0B/iEwHrDSwiSjuO4Y6YIYW+Ime/fuAt9g/
adUxQKMhVX/wvC1jyaGLnrWHTxkyPIl1PgIqAb02uQ6N+5SKGvTe0S7lExNN
XZt4lOdfHN6nN6mnAqJM8Gg8zFt7PyqBsOynAGQNmqwOo83+ah+wnM4/VJdg
+qOJB1phprDanBvjRVbHOTwpKXo8BydLLxL9h6V3MxOTimE80eWTbVi3ZRwE
9jAPMkdu8noaG7hIrr9MQKoPQcy5/YymzA215WL9yH5lHBJe/Cvo9NRUxv1t
Ze5xH69ukaQbykbPaJcMMIPImpGfuv54nfDo4Iv5nDQMWuSf4pf0LI9jNyST
P1NWqYu7RAqZ7Z1k2LCm9q1l8TgEEGV/Q0dpiXyJxgXclhBZdiO7GUUT/Jsg
fz78A1l0NtNfQXv/giy+mhWY0YkPaCX0szoOVqptBz4RzneLiJJeF0/oaFZH
MFaomB/EFa9D3q5FaMdq3xAXZK/xeLl28YwZuLUgvTwhsI3ygeMswsCbE9eT
ieNg2U8UVVl1+xH/WQ9FimUO9isn5LJxvezE2OxXVd5mkRPsFjlTs7pXfBvo
Yr+MqRjA+rRPtVe5oiAnaZwAHk+kK2ITkorvK4WpzY2T1H4ZyA3XGEQXy/01
gxvdAdHDWwHSm0fiyHY76CtvJ0DKZsri8gPTyoETaTcjQFMK3i2v2d9KSk5H
8XxMEQ15yUp0IkOn1T0rZLYrzgrrWX0cTMbzmlO0Gmug0gwnJii/Uyy0IESw
OrIJXJ2SCAyXWg00fwSkteERGEdUal1NDWrujh19tUcG9fi2UJftO/7mQeuW
LATRfuIQDEp7c9DdX34YCtxkMmIXGa9xM5w7C06E+sUHo8SVvPSXiUbgZiCt
DEzNIbIRIxJTiIH3gocb4+BpFPxbZx8k68uF/O0JazN3PlFTDRlo01VXlZnI
eoXkv1+jhcfjrd+U1szcB4//M0u2cEIyJZBGiZdv9wI3V0FsWdVJ4OsY9V1C
QohEn+01LS6+hcFqm63bdCOhqnYBf6gUgZoJHHEkl5XpFpRj9rIohm3OICDk
hd243kqFP9LHuNJoBmlATlJ41lSiG/kgjcpCJr67lcJ6IXbBmXheuP+lhMhM
ky6aSQpKrGWbACOq3BUstEv32e/T5S31BNQBK9dUIaasJkFMhoXOagXPH6a+
smBkT2CYqJ8X6vCQxWr5QmBCQCiz5zmcsgITWDNpB9ok8564oiO7hYQhHigA
cQlf8lMLnbFFaeRVI/YkVdrPpJNNJCXo2gJd2a/K5V/1pRvjj2kfTyXvNLfO
oZ9eFLU7tPNk2b7e8Z1Rzuob1sj03dCOFnFieeraC3K9UFwbukUVeY8zBW9T
2EXTAjZPH+x2ySXdbcB/zZ5+BnM2ZjGaO38TIt+5oWBP+5cuM0Y8O7JtOyIT
xpWjiiWhSiHiD43znQNA2MCn91+2do5zsT2B8QnpMPN5Ohcwrw2CRlO07iWG
WC+RMzxjIt6WRmAzaPN4C34mS575rnPIzIrq8aaN6l9Xb9gftgmaK/2lgNRY
2ZlVe+SnmbAvUNW9MwlbYBkwe56D+pldpW8z7NTcDDzVX6o3ym/uPS319INN
nwwadbMPkzCtaVW6DdZYavCeYq0AuQ8IAmu7+5Ze+VJl+zmbrl4RqJ9mHYeP
huyZ6unq+khhs2BP0Ys5PbAxuDrpPeKIjF6xah3t4e+tTjElyrdUjRl7ISNc
DCtv7PFiaj2oKjY5pJ9oSngid3KjigKqjkRIvYB2oFntiLw4fOCwicCQ69MQ
QCkqvUF7n56/gQayrRBW+MQN3pS2azugZ/Ti8Wodh/Xx4v8NHFIdLJC76tgn
e2LS/Uqacwhutkol/lxqdvVCQAlxxsjoKsdLxfecIgXKsIVS1ocis0ny+9IE
trvT6FDyy+DF8APmLXxki5I021atUQq7FjLw1IMTvUicPf9wQAfGeHc83uMd
sVdXd2ZCraxnWZSnILuzjgNj/fWI9JySZA2O0GBiSb2a5g2FJn4KN0EE3evz
sEJbYt5TAvf/rJCq4cuAJfdX+sPANsQprDioEL/2IbyNybpS4Q9AbSUvq+7m
i5b9j0pYp0+NrT8gUzavoSUwFUjl9JpNwfZvgq5ZRxPn1XnnCw3mxfWf54qI
jbUNotEfAzW83SrHv8WNKEwDmAP1HicWDAPXsx9wJJYraHk6+Ggc0CtRyHEw
HJdwH3BrPERnkk6gXyFrW4NZV3P+WMcQla11Jcwx8/J2/EDKHtWjICJNfm41
hvvdeVnrrAakfnmE53hJI7Tt0XNmtmfF4NYFNS7fI+0Hxdpfb3TWpTF7DTq3
ZRmTqiNCuUQunLhBSn2ACvDK5ehLBYQFoCml4o2eaKhSfTBp7bGoPAVmDXZQ
fe78KQ0kQ4V+kA61DeSbjAVm7gM7CjI6+EAHt81eOOyrPtFcgMcycCCGbI42
f1+M72LqdSqcQf+nC1tPQnYc2PjY7PK6j2TJO+cShLdTH4vQ1rmxxovvQGaF
Dg5IcOiWfNHuQ7RCalah/M9q8e/cmkYywNuCm5D/EKIfB2G2yhFAuyw7b67s
uNfczzT59DpsteGe/WaVxbxqGLmjI2U1MoNwIOD9/pmCFLPewz3ffjHqEU3U
DGRw5k8bzwnu9nk8UtWoU7yInvG0n+rl4unCDUmpjBeJOHMjkexAG7gump/0
ytYgsgvqjY7jlkdmDZQWEA+7TBQKblHC0yN3ZN7YKLTvK6hWB+8o6mzPDPbo
mcfQyUDdJZ+LqLZUynVA/NQNzSHF8FdRlc+qJ07ykpj5QvygewjhPMeXZPuA
pclWS2Gnc8btcz0SNGmYju1PtTw7bfhrgQpT+oz/JcxbEWo4w49sGGHXlu31
5G4Vpak9OHYBTYMObU9boCTSWltaPYTzBUj+6txOmzxNnCJtozJLfsTi40wZ
dZ3zSIUOL+sJCvc74ZOT+9G2WyRc6B2hWEbXanNXyCBXI8TsfU0iAKowKVsv
YR7PkuaX2kl+7h7Ibth+3JaY7w+YHoZAkL10Aa3e9khdx7ADeOOZXfZhN5IZ
7VvC1f0TTwvutzHDAvOESVgNgYeBohecBY86BpyDq4T189WimhdUFl3MAMLk
KdXTVOVKmIHfA/A3sSZltMAFaEseDrjAVlD2RkAwUVFIv2h61qjTlcc97E+F
ezjhxFzXrXAHMQqrtYcK5jgDoNoUAuUbryhBwSSakyJ4XLaKU3QX7ruc9jYw
VHvTIInNbj5+KF+KY55gLVMh3gB3SIxsQAigemCFUfw6FGouj4RFmleSCwnX
AlFfug9LC7WurOirIDnV6pXXYhLqSlZ7auqjV+d3JJrwFSDl+ctJtAklS5gZ
CuKct88XVkthR3YgrsW6hY1hQcNVkz4DX+7nIJuICguV5dKrFKxXCI7CP+kJ
FIi7d+oXI9yV4SeDZo8C+QqkGn6rOJdfuQYHcWd4EC5snf8wJvedjDI0rGjT
yP7lUw3N/Y4au9SaFMPQwRmUVujBwnctiC+gbVxd0a3Hf1fxeUun/501MIYq
l/kvZjcQk+bmBtwtioRH87hBrslnQXtF6FVOiEy4bSLu9ohigvSmpb3C+MpP
x2D/NsAj+cXMKzYbDZEABsTmBXSJ4xnJcOlkd8Iun0+U9pzm1kPTYznr/zRP
gCxeBmkpSe9deLeWnj5LYdAaN8mErFTSEYVkOXMP+h03DUXL35BB/nu2705U
HYY4+vIHExLeePBcU/TTtviGN6t99fp1wTNeitLgn/sAn+bAV2gn8npCzW0Q
K/ClQEcP5iBjbNMN+cpxtrEYwVOMj+ESQBVnDjHF1loAwpl9BwETkWWXGQik
b0EoVPUld2YyPjsS7/3aO5d0UimeV7kwhNbx3R1IMuhexUqkXUuYnPwq4HKb
n+Vm6EzPpagPouYRpj8YRIx4XrX/0/+GebKzGMMD/yB+TTVALwK+V5E+qYUz
ZeaIztuQ8Yx++GQHyK6kZB1pHXnBifri8JDeIDHN52sLPHF5UvDEt9jdTmNl
NRn8j7SeUXFwiYTeH7VgGTF0/LasSx9fZ0Lb5h0MYMidMwCRKq4icAVYTzrw
mUKS859iHhMZnGvC22mRYLcoREfQ53zJJTNWIaXTPhcujSoJYJCH+VA9fiBk
YXGAkcS4Bod1DTX5u7Sdd8NKanOMl+UrRPjVgHMcm6ekK3bf9/JHA/3whpLu
tD9Ba9sC0Bw6SO9DHnCLU+Rw/zhPlhxtNop6VjmD/Xluk/dGbgatpbsRQQin
9+b1sJtRWOq0JHcDSnWDYKT3FpBaVlG7757KMtSiFEI0mH6UFBSzp3srtCU3
Q+0ZcXKVGXI7/Cm8uUQZV5ePFecp2RJ25HYIv8ZNfqo/vvmnYkauTU906utV
vrLUyXjNLGRt0oYbntOBn+nNDLqaZmvl+//NdEs/tvmQ7YKCrshXjT7dwKtx
ec1DYeLVjUzUE/AGo/kb75AXIa/ctkWdSqfZn+mR/4NVustXM+va2FTl4IC0
Er+28qHqxt9UIVYF4QX3kZ9/gtrnS2Zeh6T8DTaxNzdFYiqwjmFR5+YhcAwa
b4MqfiboR3ChkudXQil15Hp1vBAFahzjbooUKck3Ge68htv+Pz7uEIhZsSKj
qLl/QnrnRlyTS7McufMVJPAHN3DXnII3euORHkMj+U1gPKbr9ZtBxggO7KNX
rO6OMz0yQHsB3wQFc0+sM5LrLJhs5N3Wbrpr5lCjGjpiMLVapg9/rcPbwN0d
XsOKlCgNNkQ4FNl7WQc5hH6FiQtXOhXSyxuIONqENUXbK2k52piTyEEzN6ZJ
XVm0LWQN0U47ukOUtA46ba9j+cFDQkbh5n//QZ5STh1REdf2gmDreO8icsdC
QrUTf5Rs9OZtP0fFFq9ANb1ALjtIH21ZR8X6UsWiBvMou4SrWvKAFEwDjXIN
5Df2diJnXEPZYilVS65D7JNrClnBbTg65gm4fCXjGcPub+krBf5iS9d1FSNE
C4bpNs2T7LHtDlNFgAyzpX8gtp9nLg+x1aFuJl/1m6CyccVNmoLbhS20owr3
W+mLKSZyUoRz6lG3Pif7YpV/0Qz1ih1KckDpJWPFjA8gijVAYHj4b4mBd5mt
ja/0kgBB6i609aaIniV9oSNwznNy2MxPWLrKsU06zvQzlyZiggzpHkrlmHry
ZQL7djacN8pXr3ktwVh2Naf1c0t7WWQr5FGK/pY90Ih/bhra+rA/ko+iesIb
uroc0k5OOMXGPv2VtbcVZOzyjKxL5GsmD3HUJnALbp5GzHAcpV2u6XapX7a+
Mmr1UU62o98LVB54HUp1Zubc+7r7fjfSRXa2H3A6Q9NRggJehqMY+3ymf873
bKTkumwi/gMUNXKLtQnB/wVVhhxOjVuDjSfSy0XTHFiLrqdKeAHt9NRq6FxZ
djZBNj7uZJc2iJ85AuIKRNik3br/t6RY5FQ6YfutzZZ/vHHWo5PK/sPxI59O
oUU/GFDhw44pALEIwIHtzt1swDjTrhWKsF70kcZOhYYyahqb4w8QrhEeUC8j
blsfTI5a3SPBQqdViV89hyNyz6WgJXi0FBCAhhogyGzlP6BAHpvn85ZwIHlM
WQXDX9sTFFU37IxSrT3Ymi5VPDyQzXcd6EOWlo8HeSmRZEzmBE7J/4skj+Wb
z+jf1g83oCDRqIZLNGswDXBHuCZnR+ozcBbSXSpsBo3C9l0bUI/fxQglJutl
LCM9m5K7XsQ1ew2qy2Kz/eJNr4jbs1BrZa84/kofAlFTHNAnBPvBan1adS/b
+UO+ArRywjLMHd7JOlgenpgi/KX0SoC95HvedqRYXSn8HQXmc9dOmkYpa73c
qhDNBp2tsIBEkunA00kQpYdhOswlKW3F0g/DohczeHzRN3r9bXzE573tPJGT
68y408J42bUcTL9oLyUrL/bZphDCM9zX1upmocEa14WBsrPDJ70i3jb3YuQ1
ZLvgERCX5lec1x8pBtBJ5tttuPHVJmloTIZcGRmwDcbbDBqpkttKshkmCfjK
6XsWjKlg6/8N4fVnT5XQIrsL8q/p86QoyypNll0akOUNmz8gjadxY/HdtoQK
HU+TK7l317J3mfov/UsXKWE/jA0e1XaXxPLCQ5V2kn7yYHyoAybh5Zm7cocH
2xIxxrjF+fo6mqDR0NiIxHBN+B/9EXz35kiWPGRpLvyck+NDEAyd94Lbphqq
y410O+HneIKdvRopWcmty0Prko5jAbQBpODpxwWAYy/mR69ZqzqMXNQY552f
JXcxl/f2weu/4NQTQRJHFpEkOb2UN+FgVwIReSjWAJKBJEb4yNzGaXrGD6F6
jCZDdxu3elTcS0sSYdthRkBV7/eTelx22qohvXwXE58rEjPBvvlfKBM45s7a
q7duwv8rvZhSvCn8SZlh958fnVG/V7pOyijuDle3at2W0zbCkzMhfRL9MfRj
0s1mRnmmmnwacIPx8bM1UtrXB3y9QEja7eC9CeWhQGt92oGmbzkm+gntshs1
ICdbFlih+m3xhGX/85FMmFLbvDlWbq/YNQ4qarIeKWCr/E5NZNwGOk7gKdA2
IuMzjfHtFN+tavU8TQ83BUIeB/3Xu04Pweudcumf+fjLgtURahlA3STIMx93
BZE4gB19yf4RvQWaKdVhKERUlaVas2vBg6vseZex8HUP6JqtF8/5sfkqkqEy
iJLpeHjoiFr+VdCYuap0FLe4elMiHnAelQNqvY3iuEUBgBTqwH++0iQng2Fw
t/RKF3/+pHYh3d5sE5bF1tYT4bcpt5wJckugfVkpSRzMxRzEuVcwuRGXitzC
Rzxk+BeqPciOtewiWFKTuvZsBna9nxKp1DHakoCjVd2KzJdO8nomv1Bbu5Nh
WMWP3+XWzX71OvOW/W54g4VEJdThNcg02SOXFhZB5ksebdQyqXv1kfrZWfwL
MkmNDrBRyghZubRmvb9w1vEl23liNVfJfjO8KdC6oBzms4zsdyqHZ2PLRm/6
DKB2daQZv8z+wJinMP1mmLWpmxLT/GG24Q58LwAMO9ZSySdkEqzCZeOWEnBx
RQ4XV5vDQYUu2JtJVhsyrwq4B7R3qT1DfEGnohCvTa8cF1abuRUUpYZ+Fn+Q
zX4gptWvugjXB3KL37h1L6pZwjony4PKOB37Fpz4q7ySwMPhngQPr6QKlJy4
SIjVCIB9RZJY/AilOluANQgtq41GUjIztMPh0m+B+BTnl6Iyv0SJXUzhWz+n
HzDDVs6e3XwK8jZ3dKgSg5oasbKsIu44uCdrtg9OvJG3QqUSgEH2d4G0KAzX
J3UXhULMp/7XbGI5M3YI0MVhojP9NEpeen8dT0gqW0S+zPvFdpHRUxRZE5l3
WWIdDqqstxYsJGUt5trvOKQXzr7CnA6Yk1FzQf6ONXKuGj1zQ9m40Y8rncam
/K5Muyj4jCj62DTJ86CIKQdNVEp/fbOo8pMYVmOdzLoN7bI+OTr7WNetMTF6
OcA5VSRh6FEMEqxhcpeT5e6VLWJ+p922JV5QcKg0Sp9Vvajdmx4H0bGeFI8N
SZevR/xtIpfSKcVVLxq/S5vE/o6wY4s02NHl45imSZF3tkEi/Eyi0R/SvtYX
D+nnm+eMz11atEmzbfOIKBtOIOxZ42GzqCt6slm9+HbceukYpttJ5cP6FJ7u
gH5TvdyKwjwtP5RzuOtBT7opDXNKeppOo+xeWczE0vRTbuXvvOGICwEIIXmE
0ubRfDSzb4Xa41z7ThTqmnmy5LCfiKom0CJoSMG7Hz+6wjaFEzJ1UrCH+Sj9
dHuVfnj9kkrfCSOZw8VX6W5FNiKa3CBhnNF6qzOE99hnWH1YvPnZJyt9sAnP
/DNJCRwXGhWlYQo7vmT/XO/GxMrCMl4NZRzSeOu2yy1O/yUEckFPw/rf33Xe
npxk2nA2pChlwfLGDwcV93j4E5CRzPR1vjpEjiFwD2IixPfXgGs8ojVx4hG3
Z4ptXnm6e0rh2kXhRr/PrWP9AWiFFoAxl6U/cyq1mEzJsIkEVx8Bs5LuVrAh
uQvCmFtp0bPA3zUHO1hB8p0SYjcbgEmZJpALt8b1lICTpEKCGJ3gCIl7fQaT
Ev1IGsU2idj11/0J3pMyGe5fbr6EVJ6Gj3P7xoHsFaJhM1PqwtUccOPWygP2
sKypMvbHZCT088Dipu1yCGoVmWRT0MCnh9mBKZR6rCLiR+nkRvd5P15WghUH
LRLagnlZXFkjArXIZLPnAKfrwedFXYfOa//JlaTckt9xk1z+orRT4izX8soj
qufZ3Wkduddd3eOHdN3Nt0tlVlf3lsL1tLOqyhGMX5vGRYpl/0Vb3Dk2Fr9l
DdGz9eqlQY082a7DhcA/aaXmOruoD+fFeLgesvK5zcHxjOepKDvFLTK/fMCY
71RakYfbVYWRgBjLunYOiyqnLjhx3a5lVMRMkqKAC8RlNIYfP5wtUOEtE7nh
rGfz+Jify3+K2jewP89+l8I/1IZhziFH3Y56sGHVurVy4dtjp3a2gKsiTHNJ
3TsC5+0tWny2xsSOw/nYjl2HQIyixX0ONbWoMMw4E9ZF1cy1+ISh89xgS/mG
QRf42jHMSmCGA/rcBK0LB2bzkNhifsFYg6vby6wyz6XX4xI++3NfgmpiNR/Y
4n196K5KcBQW8UUDEUCFWW6sh0t58rN7iN5yyABGpn7jllvs2BSuWwoO0Amy
fS/OSGtRAzwc1k2PFKMgSQGvmMCtn4lh5D1lu6z/QaqGiS33r+Z/A7WrlZiN
aRmCS38O9N98CEqSidx3ucNVpQf7CIN2wxdlmfWWwUXpjF6mFoJnTmPtzBwv
gzU+92nXWMJTjMMCHcDv5cv3DyxCdbr2MgaiAXjnQT9icR75GUJ/PKmiZtZi
rIK5uqSrlKiVB59jlzl1Edkh+vvX0khS5/tLZq8F23xUeFO+7XfaYtHfEA4C
whxN08wjKk0FRUzcy7oKY7VSJJhs7dMFdQrBWQke4Mxh7Ps6v83wSmApTMKz
3NNinnhjZEdvy5RSVLIsvc7xaLKMr+1kAgqKKUQpb3377SROuK7CQmtLhJP7
gAc5o/UK0036o5rtgiqIEyGyVOpkXVwbooFnkLFilPElrLghyuVl2lmKWWx7
17kai1xKqyAZVAA47vgnkG/t25y84YMddgz1FsW2PVpbTiiTgpdHbqN3Lkwq
hKoM+f602vfdDPEcBR8KRkUU2p8E+Yx3CFyffQRcDCC8I/JHxt2BHUMZLlAr
Y38mj+nKy/T7DkcLj6cvdfqhmyyV1L9DGH41JBVR10AUzr8gKh5xqTV0t3zm
czrlzmUKFnQ+Rs8QuBLv7Zvo+EY44wWR7e350NovEpdmadYrQ2JKYEG3lSYe
iPQWw2C9CddX9fgxRc3InFFMs7u9SARWeBAr+4AdUK3bepDIRoBjXJJjD6XN
QPtOKuge73797PaDkmvPiTtwgIBnH91UwN7Awkg5doukaS8qeIGM73zUrVXM
KcxWloI3rezgZRCPoqlPAh4VU2U2Rn4T6dZUEqIQ8sl1bta/bcnbOBJliIof
wIOfHIou4NyJOplPDa+77KnuhGQDkPIk73hQ5EVbTLp3ZkhbRq2eJkjgMoPo
EBgS78tkLPePT3+0M3v2sacitEcj2XDuFqvxKdGRu5YjSA+1vp64teNWau6/
twVLJdMEOJIUTxei1Neol/b0m2RqKwCsq33zga86FIN2cpTqc00cDpuqplKD
UXY/0rvmbDWmHKx2LbhrFk/aIPATNlu5c3LcePi2dWGOuDexsBf6r1PijDYs
HWJAqMCws46YNyIu2GPKqQq+yYyrWmQCbQuG1MCMiVBH5KSn8rO/v/BRBMNw
1z6QzGq2WG6hW04mGW4ppFv4KsrinaFedWUArSmu11UQrEoVu7GWAXhLUULT
6DrIbbqOqLNDlSydR1iSaeL1JGPPrlwAKdcOVw/gHAd7bLoetWc97cYwwFpe
MsCYi8FX/Vq54l9unODXTnsqHIC24KvuHAW0tpbr+cHpI8KM/KP2REf1YsnF
J8aaQ5avzqQ36ewILZwbit95P30+oe/6O4ZmaJWTsS+Tr5BNp6RclazoWceo
CUBmCdS9EfS4X1+GTUljdvnQBBuygjLmVXKBdei7v4nx41SPJIbinjq1rTH+
Q3u/T+9QBOJWfdgjgOb2k7it6297t/my+QqtgEHmWsRhoWdAno6BRPgZ2MaK
zY2lSRjXeNCrdp9J/8OMfBMVhy5DMpZ42XYtlH3N8/FqS2Vs0rrixV7Ms8sO
FBCOP4TujJamIyVa1hyzvWPTyWplvjUWONmeakKyld3+VryOBwUWwmK+GZVU
Ac55+cqHQTsd8FnhK1ZuqeJDH5pyFQKif/H6donB9zoSwtwcBBTILT37l/iG
VqUJ9aKLzdn2eBTB/uvCTqdbOQJjJb8Dmcn0VUHjWEe8of4RoK+0PfpLfose
pGisCnqhWi8v0/Oz7XKxXpOJ81/2M9ii6DFMnpleZoUxMVu7oR688WnpGc/6
d8+MC90cr+jwjBfHFlLjWI7hwYO+aMHqeVzRFqUVe1mnjlzjqiZu5mTsGeJc
MaIOpmVUPifVy5dm9Sj7eZ8l4vRDU2vl88s4Z9ASZlDMW0c0z/HlYjyJ7slO
LNagpgjqXBiYLNZZb/AdTckkyamZZYnXbSrfJKlSrnxwZjd6R6z5+I9rwmWe
2LbUoWWQf9ByYOoHnfGE5t2ZGbX4qFhbEi87h1YnpycyoTNs8cVuLIdmcYNU
+9+HUKjXnOTPvM3NKZUSZZjUhB+j0KdrzpUe0k4CHYkFQQqMhJq+T9aqdOww
dvZ/YT6HB4CQD3QChqkaXKFF316vMrXAzJFKhlXVpe0ocMyrTXXTIEVBtEmK
ich2yNP1tq8Tb1iIFFdtfsV22IG5eTYbezJHicPgGBj9XGRrQonxVrAoqGq4
fxr62mlGqslxufMGtHsi7YuDsJSJrR9F/EAIFdjF0vBbkA1fTfoYjgK0hkAN
9oMIyhHFFOlLjlgD1r6IlGxDovBf7MliPCweeJ4GRVKn1W0IgGuyC6zKz1d0
bsDeqciE7gWajNtU9RuSB5dqhFFb+EyzheK/iihlwAlyi+mNGrR4ntRg7654
5MvGSG3ANLHLPtkOPdrx073RgfpOZQzeKfHkNzBQvyXSOVjfVtV7mZPIJmk5
P/RdObP/V5806zY2cIkCfhSVcHmjJ5hZh3zzThA4nONKITmYKT+wDUyupsC2
pxOAoZEaW2mdlsaJwy8wzizREQEcMaFEAkKkildhNjnB/E60yF2i4KYr2PP/
CfQvtArco9dUFJ0YFQTMLl2xJWjXMVf4JX4jRmjAmPel1K69gKG/zAoZvIEl
JiQr78jMjHT7sMt6TdJQ7yWYQCXAtLNX3fmVcRyd3PlQswsOONK/AEReguPN
kj2vD2weUBOtraU4Et5b4VL3Uv2DOozgr2450C928uZODbhkmfimsfHfpgr0
2CkliwCFT3Gx78cEOc8daZwJSKSn7bsbVk1QwuMX7onjcM6CKiQxUJEsdUq8
eXJ2XbBooEShY8vuIP/JwJHVZqkRiVe0zmSzOzYybaoXCGcQ40p8FQcSO5n+
o9dJs+8u/sh+u9FjNzqkM2NBhJN7BKpxbKfI4vQhqaZOlyi8FqMXAX0xd49G
YIWr+u9hgMdX1gea0X7SrLT18mYL5JxIKHV4jcgy1Ry+paHsdJd2oL+zlly1
D9XDd5sOX1Fd61Qpjf84QDApI5J/g5lwfeqorDiiTMw82JdVfTTJN4OhRFYk
i4fg6g7YTXQYv0Mdv23JghXmpeacTwRLFkr2JFY5CBN12smHXHc11WDw65+3
nL2oShG9yjSVyNuBQ1Lg0Bkmw8FrOwwdLfZmQok9gqdZdc8/cAEpJDZ4QMIk
LPXzAGvLIjagNbty18KBtoKNts+yKvpM3Sy+bnkM5VM96aFQBqjAsexhtmEH
ueNwPZpWdxXlyRzqmSObZXJTXa5yS0tGbuiIVeguqczONIFys9/y0QPbSEI5
+QvpN5z9Xf0h+MVktIWXFiAhTGzjgmYwb8o8uDX/eyw0eFHp04kawaDJbdXg
AJwkPVZBPGIZccbxRbPPUxCk3xb9uZqHFbuPMpj4Ww0G3QYH0Hm3LvBy6jIb
v+Zrz7VycFnzGp2Nk2A6Dl5Tk8bGW/PkCZyW5j1gWOgthxRB2utIi1ZwfLUN
ryQl0WByXkzHQ4IzElmUd3f9OeQLa63uKbCCqR5NWHt5fPNk4hBPS6Apt1ao
ju00fZN34WIAMavPYPmASOLnSGEOmzguj0IyoHAD6VPF0txC3OpUnNyD0FB4
o6gzPaxEAk9t8a/kE47TtwjgIKGkv252pu2RguPCkfXlPgUG949L0KwV96X5
4Tdc6jX0IV+tI8qP/ckjJ4QtbOQdsGW2F3vlGbAbemW78WURCVlg+inRgTGE
j+2hIBCa5hfF2RzBTT5ePGb/SM4PFIlzuAraLL2zq8eZQbaEZVJZbCauhxmb
0zopp7QvXuiWh8z4TQpmW5fceOxdFuQ2VVpg8C7EgOnY76Z7i5eDK1Be8rW6
8ND7JcPRvU5SysW7+RL+c7mnsPsXG9JO170DqvBeW4ZK5CcJB/v2iJwaCSvn
1iCJF2hgJ1JQGRAU46u3AQaZuEGBzw4d/cONTfhWRZLhyziLsbPq92Q+vmyQ
KyuVlZSIN3l5DiuIS8QxY9J3M4Xawdr537MIvHTHB8S9h+a45rBr5Kb2T0nE
nQBpLyjyIY78thzC7qkRmVbRe6hT6hZ12ZUJjbGC4xmTBxsL0TxCwzBjf3eU
vBgfVMKlwIDR5UVuBqHJTGc1EwMKwcEybowgkgRygB5JEji2cp40wFZpCI6n
dOOvcE6q476yL+EbSd4rIrco5srZwXHF+J5el0ZiUGvhMVbzToEf4gZr0sAP
Szr1P/f2Dx2R65b6u9dsZYyA3m1LDK328wsIeNdDb/WX/aYxvodxPpUVNQvQ
mbRW6qwAY/MhKR6PFBfpKibX+XMmnEszDnWwQWbayC7AuEYtb+7Ub3yWtvz7
uJX6S9u0zn+ymWBTMOPosR2RzxFNXj292UN0gXpk+L1kPps7H+CupMLjxE2Q
64dKN7QURsartcWeMVuO9sLG6Xry1U+9LjrWTB7Djwdy03Or/BuSBoTUZlg7
i9hVSw4mvVcInkM5UZmVrbw15RAgYcF+JT5awqp3VITjCQqsjO+foiJE+Xw2
sfCjLpwpLEBr+a1T9n0zXMYjlTDNkxOovBmQ8/YeAE8GwTUkx6U6CiJwIE2B
TltMw3EGbjoguJwkAbpqsSy21/3C9dnUmjY6tucASCBlLP5X2hnyBbUvwJyc
pGclGur2f7iZI8l5zLGKs8oUJGFYb990GC+MREpj8zw4U+owrHVw4EkNO8KF
datwr3QDRJ3WuNttQnPq7kkd6K1d+L4gFXzQT9motyM1/NJdkhambD2KP7iG
098luoXOPXadbcZlFgxdwtWAC+24SquXyfwJHkN4urUQjKG8k86TDfIk+AX4
d7R7IHqn3SKulJI4NBFcbzMRojY1To4Abwr3Q9/TCM1WMno8ctMIWZvB83nx
O37l5uO8hSPD5hXWJa7KGWPr7fJTKd/42qwM3mS80cOT4CN8usUDAhFw0gs5
UpMvXFbEytZ4+mJO0NHHp24agshlcRqpuiAx3/2AKublFAZqedh02hEeBybx
dFX7KJtWfGmaFcBMNnrjZJLnPGVedbGoPYLgcWdDS21XUa6rIwYyLPMKw4mk
yXNySW3Cc88iQmla2tmZPwETU+oOKCfVBfoVSYc0zI73D6rx3jv/vTXqa5QF
vVdsYLoSTq2w/czhO48xXOBaFRqTVVVWi7QdYqP2t2MuMW2a9LlzM0DDPbin
tGk7lZTNuP6ugpkJjZSSW3MTAgq6otVbC6i+Q3QOeGenkL61bzVtFQtUNhX4
JgO//C4OtZpHlPDh9xpubuN1Dmv+p4x6j7ChPztqo5Gw5OzMWLHEdAHT54vx
AvZS6q1g9UGPVYEWdf/qdwkh4Zycv7nhhlbFtED+yyhn8TrAqkrr+BFpvmY6
qOZXPPj4FptqxJocqjhdlLvJDIum0iHb1MLgav1CXbZkk2RDkTfzaXrogshV
coG9fbdJOPV+VxSz4vqr4JxJjNWh+YsR7qk/R0qys/0c7/cd9Pb+0I5SPA7f
cQ+hu964qRQCvE5/1Y91lq537WKGO1CCfOUEiJREKv6llmzz0r9ix3vwnDdx
+gWTyS8k86eVYGsUWH7VcZPHduhLqZDHvYi4KOJ9ggNqx5eLJAIYgArgMiKa
cj2ACLdIe+QAEjOnOMJ1oVOoqRpRNpJ8F0f8yTPp0i4I3tTvBWUzV7O/LuZb
QzCqbE1DiUcXzLvPflPdfMgjLmzRZfWVGLmycJrRAkqdVF6RRPpzd+HIghX5
Ot1GqL7uIVecQzS29eLrfvb2cGZUZgDwse4eqNZ880BZewmB5JHKcWm2YECD
fck2BIQujnz6zGYx1rBAWt4K1PBFVULY7NGsJI7mnPPNB0jo9NJQ8Kr/DjK9
WBj9yaR2O5BNbvcHu8LZwLcgOKdlMq7dOAKaTfpkCTu/PkVr+hImosIC28ZF
OZ2Zd8lwylluNyh4s5aOUV6eu0JeuT6DnyaEPJjxQGNwI0nQjnWN6kelldGb
hAxyA3nao8/92dnHWP3YYt54ZeziWxsf9nHiGGlIjJim+KtaM9srgSm8AnIR
RFiQmIi/xIV70OZyYZoe/YRBDv8qUXq6YLseNypHfFKEF1mu7V64uy2Uydy5
DaJdUOVOB8ToPXBSnHFwTOcdLOqB9xNiC4XES1fHmBWHwEAiozHuNcW5cQLj
MFepX1pyVEHnJ3Kir9NObi45TrqOCH0tO8c+IQERxt/PGIjtymnp8ylDUYGK
2L6zR5Tch0y4osGgVxzcZJsEXhn0vEdLS5ECeeBdVzJa88FdmegepLJl4x67
ldELFB0COM8yhhAuFpHL7b4rKRu1ArK9KuIx5M8DdY7qmO3YAeNkAIsHXv9C
b9ys90maGQC+WDCTxygc55AdH9kMMPwIokcjFqO9CVGusF86p5O9RW5x1SL1
zS9++++mSdIwRfDzuBtl3mtE7aMPkoZZMW8O7+rRFh/KwZDUgrvDwPg/KeUr
hsZOLsJ9z/N2+lWxxWm28Wfw2NeWq9MhtGmU322Gkn9tqlPaRqihEiou7EM6
e1BlHGrCTZP72Di6Qy0mFeNvjqdhKCFDDuUcCpfqtHrWH2LDL1reBhJ1FNvv
Qu7rDtGVZbeYVhO3KQrJ4FywZ/DIoPVnjapREI2tGxZTiZpdKgqf3Q0u9xLQ
VAXAkTzyuOLg3LCoiEQTvWqTAwaoAX+sUBTOcbdPnAooEUT+eZuwRru3g4lj
6+7kMgB6aVMp1oEaLOLIDzgeYLXr2E5Q8IqdeByakwlT9MTMfDbSo6VMzGBa
weNeCfEWNABGTsY0OTV4EAqaiv88svzx37uz+3ikNF68ay+goFbSio7iQaOy
Min6iIZ8tXp6XUboDY8aVHOmZtQbJpEbljbJ58fZGbdspzBTnSDcW79E4MpH
WZE4G/zrP8Am1rMSr83PMjqhdwPSPuwVxKAUPHgM5ifOM3v4gKP9Jbab4Z/w
UaOllVZKAcJBW4eY04A63Ao9D2zQytyuHG9MszZ/Idu3tInKLij4CLecsMsX
no86k8eUw46E/gaEzdLd++NexDBFZnsbn493zg+OZWu7IEp83g97THPjj5Fn
Ju1as8t0xrCHgYdU25SyfPnKu77+f7Z2vj/Iro2x8ys3o9S67eVK8lmv3M+i
1nmdbsVNBFiMaEbtO5eCbwhkS6BEnEp6TX2SvzPOgU9FI4vuRR6BP52TO6v9
QYkU9jM6aKxHf6fgOkFowTvcyK8kwlumWyBia2ezb529huPVl666HerJs5it
kPdzTpYwHtGtJ23ail6mNJbOV+6Xrn0wODQEz9pfzWR8J1Y5ft4xA0vzseK1
qRXBlOY5wYpy7pFklZlAy8rk2fVxankI1P0y/opnLKK2+o8lxXIxdoOivoVK
iHmlmJsLSve1DbdUth2ENK2RAqozJKXLYqZ4gttdy9VtI+yNdOsnhj1aJMbS
CEKGDjFUw0pxXEBRxgFu7SsURLLzKyqhzkB5xZIxHFFWmY+2iy0sR1L4YYdi
lbk0i+Bt8nYa8GutyVCJYDLACn2pV81n1/L1vqHZn+gl1Gf8PyV0aKFGtZ5p
GLu7Kb7v9tWfKWNWbO4SlV1SMJzfvVQUB/iSGUh0Ju7eaLtB1cRZNfHpXo85
LGXnFUXll8RAn0ZBnqOiFHjMhbhpT1XXeKYlTVzUXOnTXqlaxQu7HGkMy97n
fuyr7ucAfhKlpeqVJOnccOAJcFhXzTYmoMDB225xf7WLOPRqobrBadPIeCYi
9tiVtMaPYqoCnzN+zH0FcEl1lP/eIIpGJ5K6zXhuTXjxle6JqAIOoi2RN042
Gs7rI/VBpEyzOl8QmBGgF8LWyiNedgMSTz3PZlHYPRr87kNxIQGmW7xoFNI5
Uh2Ggto1rBdvBGfNVkg45yifV8wuH1hQX6THNwhTR9Q03L3/GPsoa4YLLaS2
hQQ3l3kaBZ4h2HIPBV3qQBnvQ4J6BmkQ8hFFIVA10RKp+EmijsWtyjP0mNJe
GeedjaWrZMl4WpWMba5rh0d+YEsqIhbajVdWNHetWsFZfhXCAG+bZag7yLA4
OUb28pm2EOikH5hjoURuAtYDnfSyhHZhhNVGveY5HNvB/+LaBK94PToKUXV9
2DYQA0Zf00j2iiAEjs7dklUFpE86R5SeEX7gPth+iYMFP4HxXAHjaD5dReqt
6Qg/7+xVJHybO51sbDFktKarhboHVWeqTzbtynvR9kOuzv4X3n2xF09lumer
lJqUwLW9Rfv13YJGCyUaQnfoTBOZKAJwquykrSFgF1hmoiBsgKnakCPKUgwg
M1KmPE10CZMLGaMaRQIARb5phmBgbud2Ss0QsMVf9Fd9A1I+F9+Kwybs1/vQ
OXSPeiyX6uoOh8sIARBTjIN8QZCoIKJnICyYT3KMiXaCV83951xMQ8cTaK7C
+87AQ3rberev7IB91e2hO6bEXjmVCp7dQdrBWAlcKof0Ns4H7kBcVrTZXOnc
xVZOi3k6jy+1ApdsRJ1HVDOcebq8+EQOeLk1r0dHU2B/0ImJ5YFWtgzhVnhW
cWH7LF/YaVKOfkYmOs4Vpz1TmZD59mIU84TMFzNIFign+CpebuITqO6yJsii
1zJ1osmXFmRDtTFm28Ps/gWDnU1/jJCC69P5ecPIjBs3JLrLtIEdo93/DCSj
jPgnc18R1XN3biFwt07f3ghselgYfVIgH/uycBooyQz8IPtQ705gaVRZ+uS1
HCOCyUgidIHn8ESAA8sDNIkvPm3U1+3TFZkFW6MM+G0kCDj5VJG8WBCa5m9P
+N4k21y1M/RtesDilJuwBfhjDKTcQyoiUx7GtnTh7SzoEMJV/lx+0qVwo056
ncTimy+72MRxy/oLVhww2yxRZuBpswPmlqtylx+M5t5UVHvT/4Km9Rm8R7qR
xrwrJM9FxEnFGxLhbx52LAPFsruktaGCSKdNgEp8IBK6aHXD9EXqcFRLMiFY
lkkMwzZj0ke7urbB3s/oYU9eMNu3d2OjqRQxZ0sgNNEKDBwEljQeM6yc0b3M
dE7tiZ1KlJw6cczaRRPZp5IWpDR7meKpXJdvEEd1Sf7bsdf109eDMvkL3xaP
tHCp0WVR5P8Hq7NIa6ocROTY3oSVg1J0nHn/IXEP1EpfWJKUamf5VeZIRGGk
B4M0+zj4eBwhBmYk6Pluyq0VcZgHj1h44od0fhK/WbHX5sDgeuttyfTtXZky
x/W85lHGYAzRnTn1BaV0s2I6fMeCOvwnpx0BaG3pnQLlD8ZtSc6BnZPsWeOq
MH6bYH/WA/T5RRK6Hkgo4SGleEaozMxH2AZfSeej0umffLVHQTSUkRnCsnAy
eyV+I+4tXMKnDalTP8z0cR8ete8324b6VR3Kn/PIlv5/xzEUiGdZ4+ZUxxQA
xYRFOFqH6K4tkRQYcaatYL7xAjCUzZrnkqQv6CbmBOVN8Frtk9Ydpy0WMVfi
U9Bo2gWjOdn90uMCTDXLKTTTbkY9oc4nhKZlro7Wx6t00z2X0w+UV1ipostV
TIuWW9PX//xxBF8CjcsZqPbomF9IYuVqaX9tMuHSwNwJqUwt0GP+kjSrrOv0
B6U5O5ZY+w+1a5MZZM3xQJv0hJTCNT+wTKHoDb2v1cYa3gqXSwaH9DwsIc52
Tf+CT5vEhL6US8kl9gobKnR2iGTbM6/rxRQFpybMPQi28vkKmYPWiJVtKdf/
RZZf84XuYC9vdeaNy2wreGFR2lY1RfhOugbN8KabekXRo/BU06GRzy87w1zq
scW+oKpXe2imN05esRjhdnS8/znq3qGP069wZACHMVJRS+hre/697C+X+M/C
e+YY4dEpl0cjsnD0R/qeof9mGZZFGSqZX4czXrNbvOWEGgzZO6k4aKKPF5Yw
+Kg0HznajdzjV5aNnmeMwHXUjk4uN293OmE3WLK/RPRzefITdAG4RwM27UBx
8fMtShPbiuut8noOCdwDSQ0evLgA4MZnzQz9BrIQ/Y3XIWtFi4JdH93oOZPg
du2G5gA7YM5XA4EQ0NU/uxBx1q+/tXv/3Dg5aF2CroAsfwfHgp4aMvWx19Lu
LHzpFYHqZnmKBRdbmlbUdmDnQZ9JS8/vi/5AF9stce6pdt9dorVeUPbD3cOq
fi0jiqvtpUB8m06ok0ZTRmNyJAM1xQGi3eKtNae2nrtE0Fa/i49PDUgO6ist
VLwcq8iJv8X+3C5mU/aPbKCg+Gy3G64FDUHnHwb2uGRGoRT28qoO/lak9Sfj
RtpYsQ9Jr9YWJNjzGq11zu85YuwBPs5D0dS73kfc66U2p16kM+QRUsD6L1FD
cM8J+KSTQQA5ECG+wv2RLoQsUMPVeBLz8YQeCLL0AynQmVG0Na80+bRVq59l
Y0GUFRHF3B/GTotm6mT4B/Ig3LN80wO9QrxT4KTPZ+uGHiR2tIZ8ql9wO7Cp
L0m0jbWwBkpNzJTIJ/FcIoYzW/5Aoi3HDyraCS5qhODFlrlz2TqOICBi80rn
kkEeyr7oZhfsdEKj9yaekar0fjTSppUa1+O/vI4sD2t0dngMtuMWsQIu7/go
Ly7QMBwcUdbJpSlxZ6/vKhJoO7YbJt3sx6IoX7t0/Mnperf8wxiokKO7eTGe
sqRneSrez/7YJN24eRgMzy81aIta3tZ2z35JzF2A6L94JWgb54eSjQzQEBbP
cV3QOYMtoCLLx7VpGVMHhFzPuY0r3vV8sAti59do2OiuMAUzKF+1QB8fkpIL
441B/LFTx88/HDCrh6ABdndZ9r07GOCGOKZIVhd9CotPJTYHdUwLLjGgDQ+C
dIlv8frpQJzXPibpLZN8NyCUqT+5jj1t0k+YOwaeIJUL8tzhCopC6ToJ67Q6
OU9O412qS9GBbJoCvmT6GOp7rQj1E3DzYG6EXbUyZRNCBMhm9vAJWa3B6dRF
oz0DHKpl3mpgFdpw2AZaXQR+kE4jc6et9+0xtVQq1CnO3WRy9+iQpeGqq1P+
XzPmWsaD78pTA9dSAdKXYY+IEipaS0QGF/mTAUxQRSM9Wt1vCWtn+MA8bGe1
wEImY93/eO2r7Ay+OFDoFz4KIAetT7aSS7EIG8DKIv2N4uDTbywNJYlnpzKe
A0KtRfPZmqkbyKmgryX+MTHD65NFwEZwnH6jZDYz5es+cbP9KzESo1/xObLu
Y6koku8PBk62bJ2vEuCkOpGTHfnXlPSYKXgfjjbc3hLUieXEiRHOiSLyNzgK
/QW9+Yg3ATunk3ezsrlWLxe7398UeqMsPPEthyEYB0UrHNdN1gVJ4BW1Du94
GybCiC4utUxqc6Aysydg5cBltkQySW9DxILkYh8d5mZVmCsamXrcFpeh+1WE
+ZyhDYSfGp3m7Q/MiH2gMLhKe39fF84FTxjXcZ0YJHZGBMMucHbhi7eFeuzx
yJB9MYAWy56gE+PB65l4Oc9BE14kOe5c+iX8mAy2Im78zzMYU5S2x9mVqbjI
z4KVAnz4l7471qMWIWD9o0DO8kYs65oXytbNsTOlk5aKyijpPcq5XZoGVbSg
HdgPvwiipmg0h0z5V+81lDMaJhpwPN8Atjfoujzg92pn9vJ3hnDo22TDQANl
V/2qRmWefAMXIU/CdDbwYPpuFwa73YlqoordunxVngLIuLoBEK74sB/pGr3d
BhEFmprvGwojpkgOsXn6n8+rix7qFJq6dLm9IGO6aiHQgh8WDfYlmPotR+BK
D0ynbyoFKp+T5iGuIhq39L/fzVyQ7o2bNEHURpGa4vogukpVlymW24KGQ/wG
aGdGU0oYwz+UaVI+6FFql9wcthswcNyNk26yyJpfXwlotFLePpUS8MeiOaSm
dK4k0vQb0Gpdu0c9oT7tVnd0qP3tR86wwNetnz166hgHZCxUat78KA5hQ794
LX7pr2Axj3em0RN2qbmjCY2G9pu/uZrpb5yVFUskXtQCpGxNlk68Ql6Y0tC8
m2KT2twsS+x4Hsdqws/YEIqdPPHxN9Dt1DhhN9p2t3FySv/11uR094pAlS42
dpfJfRIJ6bR9CmV6/82pT6Z7AVyWX6ZgwnRZKKMGWeBCpHN+R3MzSQ9TxeXE
SOAKAq69cZ3/I1J5QTbMDDl3/DvlVfJBxxRyaA35RvtquOztf523UCq/Kem6
3vNmKYjkpFSvSoDrh5aYoWf6FvIxTRoQRYy2KdNOZv7eHU4/DYULMkZS3GvC
cKwJvROKdm6MQ56KGeTQ736nw1yuV5UOuWHyJCQNKdLkknUkB77enxBYNtwj
+s9AMozsUH5baGmXTy3N/oocQNrbgsEIwFBnCcd5MgtHkmGPyU2gDrdiq84W
zRskMS7taHd42P8P1FuEZAUj9X6eouDtrpb1pHOf0Dcb/isyOwRIBcyA4ioH
3ZvVwo0BpdJEazVAukNmxItJUdh747iCcul2h2xpuu/4owjNGVvaz1FsTSbq
FKoXAXMSp3lsTWISD3MpVjE+RJwHErcktFCo2eGsn6ntRZZXcaDr9ypDlMIV
oqB+VAHgOuedmwcp/5nM7+MA2KwQIPI6ZRI6SFOzxO/Q6qwyAIsy+w93kLar
J92K29r5fXKhVggP47Zg7U6nr2kUD9QmzVIKbBaoCGOWLxP/EdkE+iwswmXA
/x1bF9zS9XNWFyZ+qwIzXYURGWIDHr0CWc+5ePwVHWVe3L4RbZuxw3vrwbRM
SEBlXq3QhrFLfOsHrKobBO9G9D6Rmg6isGTN2nNAo60DUpGNwhqV1baSQ+lM
HnURYgIk5ull3gGGFDJirZZrmkXu7QnauafKJ0z8vXEXlbeMkxdMW8iQMDNl
P4OiXv4YVMCcEDB7ITYv0bVtmkjzLQR6iw+g4pMSgwiIAFETYsjP5qwr5gWQ
UYcgLQ+t3CEJ9EzYRHCLuaCphxeuP7wY/w6628DJpBZWZxBdaJMEPen7/dx8
nGFy7JqeR9sYVs9S9g3wRwy06tbFQpXGhsbxRirHzEKFj3c6RC8o5QQJ5Zt7
pXxXl21pgUSWh5JNSYkgddrxobb4g3Kl/nCU/25M9pzKlM+SbWCp73GxKd5w
WPnOg3Q5aV4hiow4rgEOZmNws0Wk6ksphW45XeIendlEOWaanYynNvWCLu/4
La+rM2FTRyaum70Vj4ZXnoFj1BAkqRf83Nhmc8WezcedFaaSPNMSTubk6Pmh
QYXzaN3gUL0btNElLW9uC1nt7+cxsxAnpHzavtAV6pq3/Hn3JOybDMMwypRo
Zt7dHM+XlxGqAiEH8G4VWdqzcVW8iTtc2RgS27cpgkmP83wvOviv7ZfnLU5O
6M4p4jRheP9jR/rL2nY36VmkGLHYm7NLZy8bGFPoIAFLZmvhz1GbTM+Ad1Om
+jaHYFEsoe99TYCH39RiIJzuRTt58jfi30rZXzgvjNPBVteIHeR2ocsNaDn8
7yvC2gFj1Q+8eVZ8BRCtHc4AZsw7sPsdZyTW0fkDw2VM8LglGX0WLi13NC8v
ebvmZu9bNTJSsQrurFcZ9lDyLID19b7U8+rIdI4uZ0GdgWnISuOeElj1PR3I
rT3tSb+1/7coYsNxSIgqH2sDkVrW5W1hbvGA4BK32UTR0dtJ1BTR+Rsrxqgv
SM0bNNu/PVJhrTnAmzF1VvY2H97Fphh6hw1+N8fEwvGlw0lNZka4m3FuaOve
yb23eJeK8QboBDXj0BVbCfJh2pgfh8JN4InNNm0tsNHUFov50/Yqr7ZzqvbV
mMk5BfZwDqkKEJ7o1OQ+Z3pNptpwAcvIRtpzalIBYth7mbFOQETqzRT2SzXJ
MIb3AnsVIyhh89nAFiZ20WBRGSYS/lhEf1Y/izfH+nYQSC/65JChossijh48
tXdLXNJBOWpoOR62vdq7Dkrrnetv92gB2nKwErCUm8XHG7Oum0yhjFUeHNRV
oR76QB8KMOIWU8+DYy69WUJVXGjvcc8eb0qza6W0huHZ+mgDbBRI0b//YlWB
AssQ2tNXMHstiTf4OSJHLNDD77usWBMeLtk6kgeBeZpGaWfjPtP4+xD5ceNo
+VwbGClP6vPL1ZuxWkXgIzwIpV6RhQY1BcOMqkLoC4MyJ2YD1bwbM5e1xzc+
PT5ffPni04V1HWz8Xq11TFJ5QghvqJKGYZNq7AN+yDW06Ml+vemC2JsRuV9W
Af1aA8bQlVzOoBNUPe4bvuf9CVOgmKxenl0PSYd57wN+HxbLUP9V+caqd4z4
lwmEuZa1iroiQFSrhPmQLlbCozCYkuZYFVcnszl9pTBYOSp34ERSeH3w+nNK
fQIu44oHHZtU8ZjWWV/mYMrMszPQ9AEl9guIpALbI4P6aRPJqqY7M+NeNLbk
9uhVZWNoFpgcsJ1JxPzJFdrQSi5lsmD4pTcsdYS3cA9terF1nWXeNVoVkqRB
4KpkVEtrcYgyY6F/d9O57oF2s2+ay9/hfrDKGaJjHTDype8KKqHMX/5Ba3ix
Lb3R7Zf9WigHNUTskTJ9qGNoAykZbtQvXm7gOJuBfLF25h/H9enitey5F2nx
zun6u3OeY4ziTTfpq4wzA2lVLOqsC1xN572QhEu5krKt1ibMGPVT6G/RUZSM
gJkZ6w2U0JDv+LnRM87RmrYNVJIi+ZgpXlMUIkjXXmE6RrlSizkBGsWQCl7s
r3/83oRyE+o6rh4JhoHFi8/a8we3c3hhsZhv0hy90Gm+MX7UJFmhYYbw6L8e
BlxShU8S9fgvh8wQtGHzUHVj73q0ON06ZIDxdz2vkfj8fqRU0axKBHXqEgcj
IR65DXfJRCppEqBZl55NoEsc6IstEovneVrq5yGmLcOLcsB3oxf96D5Ip4tN
A0+G0cICPyg03H0bekf+gEc0hqZh75CpdByn5tMb32/lEAChqEdH84BDAssB
xfK4u/lYuRPTlr/kxdzOmPe/3+ttbq3GZteDXed7Z9Kwt5lxF8/tByUQrx4z
Kf2Uo3FhDUbcqEGbbTy52JXAYkQUGOwsK/Xr61jZqNv9c+sE1KdD5AWtoDYe
Oru4YGFsY/bVAyyVdhmlDrUdK7jnUTTM6GxkeZbKeFUc4QEdYVg1bRyrdX6B
5mUiNXET3zANeuOBGzPnBfHOX7uuNh30hRbYxSSYruPGIxwJ1G5W37hsyGsF
QifyhRj+DMYuyi/pcYo1F6gcx9uYKW1rb1B5mjdx6M4uo3d4go1lxEjQT1Kn
TQ8wFzuV/cCXANIht30gdHL4Ul532AfZ9PAyda/19/ukB0raX70+cUnRSFZz
WzXRUJyu6Ell1sUolu+C2MyOq9l/f/XtHSXiXyYL422KR2ejOAzdTuflSh+t
xEqW9eVeqPziirP8cvrbdyJKInJkLb+hntxkCsPl1/BjN+FXInIBmHSP8yCT
EL3KdVUFm3GG6B4oT641iQz6jWqGxBh83HSihKp1okux6+K88ut03Dw2OU3K
Gwy8ZnX8JIR6pO2OchkSJPwp+rBzyWIFkByussAI3VV5Clq0eNWQ0f/K+uYR
fdVViGbb/qb8vN3aF5EzCLanl/iksQ/v/LVMLLqX4vHjDnG1hebMGIcbU076
cOuea5dKp3JMpbXJnqMQYjhehXK12981P63SJ4JClndOFSiq9LcNISgdBUlY
YBEegce09DWtpxSAuT3tTYa3W7GtXMkoPyUs+h5n+j24giQH62rBV40Urq/L
ipsE2qa8uCyksRZ1ZA7/N89KizUiXCNWDnVm1kERDyuQhKU6TCm20nIJPUys
OSkB0Hrl3wfvEnYD1oAyclrhDYNBP70bsaGES8UlB50EX/btoNxvaQoKloGa
KkxtOjBGco0EZHXBYKZqo99RDs9fr+KAnY3BGLECNSCa2zoSreahNPxVQIs/
XG5Z9nu/eUbaoMc+NGyEmNeAzMvPvLS/UudoHr79qWGJI9i5Ubm9jJT9o+eL
/7KTqroXB/kuoppXZfn6k9XbUli7rnCrIkDiw2cNZANwyOj9o791mgZj3u3d
aJHaCHqwYMnH3pf0A4ND/B+mqGPMbCLG8tdlKJqFmuGj+/i+1euLNp/1+qWp
mEoqf1P63YVKAAso8MYDr3uXMli9q0ugueWZ0wVO4Ulhk9Kt0pnXMEr8RleP
lMlMHCzApFbSJGK14W0in3QsYLjRzCnf8UCn7A4ldV+l9t2WAnBvgtYeYL4K
/aj0ToNlfG827CXpM0/FqWJvyk2NExFYKO35c5yh26MzvaeIK3KyPp+5fL1n
xk2mM+AYMdzPGv35BDyqVXA0FRG0m5N+qj+3dnGCdxIcYlpGIOiPQ2UBUUti
cWn4DGopLzbo0LowIenA+RULC1jtzVDQ60aMg1igXzyK1f1rfqBkGEl8WcSG
NCmfg1AQjqrmavFCBk67NvsrGltbBrqEAj5BYb4An1IackMey0wwacicezoo
gJhNzVxU0LUloEQwnxcdmjd8LKBrC56NzHhZqHq6zWXQ9ePNPwQdQgRYoOHm
suQwuK4uTvumJ5l/qq3pYIwMb1No8xRWz1ohYmJ/cgcu1pfjkQcV3Aj04COa
JtEYRxK39LeD9fG68GZF7qxpam7pR4Jas0NkkN6LL5O/KnjV+NqUea4+N2OH
RmZ6uGV4ObFCTWF6cMPMqTlzAjH7wpgNpzTvwaREOcBH/rZBvKVoe2wLxfDm
9YhxCrr5TTLNECVvaJBFdtykB8RKZTZAhiCc4siyAkoe5YBVcZeg62H3dliC
UGFp/Ujk17bCWL3UTjnjxEGN8d9tr84OqElrqUS9OICbqBudAGN549+D5VYX
avB98Ndfz+lHksNR6rus4NMwouqDogArmAI+sSFZNQRMDa3pxrqVvS1vLaDW
ZmtdUsN+fWKhtesuzN+bWTTtvUlOslFC4KOCO0Jx4ueYRBfUtUegt/ZhVAGR
o6gnCW97FS3RnGCTmzc2cwPxOw0AbX5rzBcDe1QEfykdKqJTZ9hcOzz2yehG
cKCHfnpGsp1zi0gnLiB9lUp+zycnJvqA0AHlTduhUS87laRlBGqlHkM9qUrb
RzLknnPT4gz92tkYx0WO9UagPwFEzjPqNP2AKxAPkNboDpmwsZAETWlcWBg+
4MA+iFF0itCluTD7qrTcAi/1OPFDCT2H4Xj0Bw4EvC/6VrOreB8+IRGuwrg9
OHw0bh2DApfVRUfPg225awM5XmdXyUWkJ8rT6nxAGjtutolChC8GogNv1l4I
A85tz9lbtpZuej5YE76bk8x7U/sgyoGUTH6Hkj70GcpRJLtavLnDWzqFFHqQ
QNhXMHd6eIBzfTVkPonNYywtz0kDNkQghiPDatmVI1xq5CREfMceUwJo+TU+
MFcP9DRLN5kEQ8q5JoZXg5i4Km0Re38pA8kx3rOTy5UPQ11/e5W63E/H8KNC
/LBdY9aAhkGhkNVt97qs4LNUS0rAg3YEmYMT/hFSFsJuNAwFj0t6RwSv1vtw
jIrICDEmRdwflSxQpw8bvCPNa6iWXGtdF9+RteKWqqqpBa5qC3ZWXtISV0SB
3GdjR4PRcGuTg/Y54yFz8ljvla4dHJa0dycEY/J8pI6yBj5CSiiE2mYCZE4S
htjDdt7uPgtdoH5sv5SXteGjwMK7UT+8T0fQKrllWqqjC/85AHqmEpKu85xW
BuUZVvi6Rkkupiy66ITNMNFIyeB5/1FIdRbm6S34JvOLZm/i4rSCONo7Ouvn
6hnB9L1E9L7m8vmCh8cwV7EARxhJIr420ynd6hjPVqRA41cCcpvNZ8n0Y+kr
mZ4hiEIDybqLWJONiJ8CjPpZowsf0RBoPom9ymEAHZZR+LLLskcsfTFglDia
hfx7/yBsdCNxcceyaHFtMxKnZ7bu8aVRiNRnO7PXyTP2PclG6Ewi8crOZggd
mQdDQs/W4G2Kd8j6DUiNuputZZ0BybCeChuP+EZN2nz2onDeArJ3yH9/XwKW
eClF7xOgjS4HR/tiLlwjxVWAmhMuPatbgQ2zEdjmTSUTqBJV7yA3xfJkEoJC
eKobJrNMqJ75ReDv0uVxsCAQsjhDWiaciC9jfY9oyAfyngs2QTf/GaRbd+GH
i1IkcYh+ntKiqoYDWCF9lTs4uJCtXb51xKHq8qYXz5OZSokUstOfJLo+KLS7
pbwhlDoxuLt2UR5NQcbdgn0g4ocz/8GxMTkhs+srENdJZ1XDukJQ63bI3NUO
unifiNqEMESgehkdYfhr3QrFtV36oBaBSG8NXCv9HXNmLnAQ1XErMDlXY74H
2iS61PwT3MOccWhsABFDv31Z8yEIi44IoKazr69PLBk9jXkQtA9pT2k+0jsF
cBQotMvmMwKEYPJJf+m0ulgYaAbwEtnH7sfolxlF6B216zmovMiYo8mYFfsV
lqp3GkIrRJ3cAvAVfbhGg+DUBNMclJeRNHAW4nePn/0uRZZRkLvw4L6D3WPL
abAOjal/j+QjldPdOvPMgkd+BnHC+4vvLGlu7ZhWxfxNiES2ndBFH9vlYHU0
uIufKHE7X6VT1lMTMFtj0Q5Kr6VXTuGLN/TxdhUQTLUcSfUO7OqbR6yd4xCv
Y90xLoma38Z+nzX2rEXTWbSFO3lCg7kCceWG35V087KLxPv6JZx18V6dLq/X
lOv2aNKQhXpx71V9Thw+ULCnd5YQyuDZbilLpIWZ0kixVrg8kH39AeqSh+7f
jXr8BpSKG2mZxrG25jjiucjoTEja9swGtTEybvLC1X1tt9sl2pxuueq+NQ0J
wl3g0+aWpZ1xRk5PylzBfVe2juzhfjgoT1DWq9+mQJLROsZecANzFmobkGtf
JpKhx+885UWg710U7675xLj0HFY19OUjL9ugNZoRkd4hHhOIiWFrKyXXBEDc
TP/A4mr101BERzA1lE9gJ0DOwVj3ZZMJF1dQAqFo1ABe/P+j1BW6P1POfzNJ
pQ8oRJ3qZCGXILq0hEQj7pD4DsQPCSGkE00o8kA0oS+Lycj+TQMs9bjTGARI
/HS7cHNBVPR9V2MICCpzJ5RluBNmii4T3ZlbQL03e4a013WKYZpavRYwtnFd
Jy+9C/vynyGGl1GGUbpaIuqujSQqZf5tMYt6ajZjzkgVHqV5fGHYirYWiPML
vL2m7k7oh+KshTnrySGMFtX6bkYn+fAcLYz+8ykUFZPn10P/Qy6B58resRBD
W3W4y2gNFbY3FTsoIf/Rx6G5YYFjA5abXuUnEYL2bKJGTD2lDZHLxW8s8D+f
ZdNnSJYJs+Y/qq0YiuktlmeiHGX5zfPD7dhVh56rXYuqoXmKHm96DzgGtSZc
IFDQIgeepO7TR1/KEumVYQGPeFVaGdZMQ6QNi47wwWHu0giFNe3rsBtwcDFv
+uMvDLdFk0njcqFsNdQBS+oVMqXhmlyMJ39elO9n9sf7OG7TuLgLzg1GeApD
lGWCfdx0X3SfoGn0KxtCNWc1QE+980dC7X2pPLiUDz54YtbEMKDc45yuOUrq
HNmUpWRwqmQyFuCcEt/yBmZ97SVTwF1LYVZuK+Hq6+QLrVUDtDAcmlJtJc+V
bXrykcqHB6BYrvcxnliW6AibOUYC5DDKG7DeLzMyveFvGC0apdCZb1eo6ESc
SHIyPO11m3TQ6rqCN3777+x4z9wLz9Du+Kygl7kDjmVWfF55ueDg/EFjr7rP
fobz9kbePQK2KROym55mdYoJQCTvDVL781elFMKLqwHuK5wouy3qPRLNvRB0
4hggQ/jFlddzpCk+QC3RYkQGTVw2b1KV32Hmi/pgU5iw3Apv2JQw83zVhxAD
rvO89yUYmj3PuimhQBJ7kuxknOTs2XASBbrljmIF28TY+5zbwIKDk5l1KTGD
Kn2hpyWyeIlgWFeJgfDCaiDL5sMGn0XUVpEGqymOrSJPzUTJ/BPhIcB/eQtP
XHgBZHtG6hPF4jrsCWtbDwvB6MIYwMLJlzLMcePEbi/OSBu2L41nF/HvVfym
alaSBKyCHuY0KbqBrTNjniL8cUeKF7QnteJj0+K4znW79eOhHompd8w6oHZh
lzWd9VpfrUO+vaBglKzCvT3duIhCvnC24eRXDbyXQd6JzdTMi22Exy/Sfdnv
U06FjSj3HXXDjOV4TouFBRvpsDIoMobPdZvjSpYlGnSqZMwdrFZJmibeg/Vn
XWdRUr8amNFJFbC4aoOys1dzHmhZAC6YlCYa4rzQ3/IuBWqvyfCtfCC4qpZh
HaDvS4LXu3YJkYlLfLFfkiDuChxBLg+JTMu+TTer/I1BbwELUlYkvo/OrkTc
lAm8nhnA3EBGhfFjv2xyWJfdaph6i5Xq+ndKeXvV1Un6iWJ/663NtNHkEIyz
yeWTgzh9i10FBTtkwIrQeRFEVy9nloUBMJP5eMLd2PucPxirY45uHns4i7Fk
9bzeya12RrQjfVB/mpHapeKxhEYKTKBewnm5RA1PAdsIm7xX21s9xcrLhBcI
VjFCg4/yf9iDl4KXQPDnufWSH6kR4uUqsh8tU7pgT33z724WQcm5KCTG0NGL
iF16CacoX4rrqHLf4/4VmwHibBtm5INGjWoKcsPIkWr4LJy6YkfqTgJXejPH
8i41T0chQEdIefc6/VZoBQPg4yrHeHyo7rgJ92iyuIPpYgWikdNfCwNwvyNe
i9kMBJW1miIhYixM6+wFuYMCmfPPOPpaVDlo9FaUfvH2O7XC0w92mAn6j6Yc
jaazgu0J5eSrzCRTLY9i6yCPQrsJ16Tm9oZDXexa7QCDtGknsFpSlX9nLDj1
qiIdjEmW1OnGK2OAHga0ep//lcFDDaPo8hrNe2quBs2Oa+Rf7HB+NLwEOuD2
GVK9qmedsbcphvoPT9gGxj0doPdfIjhNZhqP6Lo6rQFUeLZDDa2NOZ53Jyi3
NIz+lzO0lslzWg3vqtNnYYv1Mohy9xRDdpMtWVZukqLf7vq/Q/P0o9khudjP
PzXQcx9ecvuvOdy1RXYLxTLcQiLd9pE+32VS3vTnfLnjBdCpITCToAcl1d3m
bkQjCrVM/ILzNzTo7K0adEwnIECQMUJs+Efp2wDUEGxtPeR/mm7fqHuqnhlH
KfL8gfN6ylH2GhycGUOzDfvkHK8Zti5MpIOfiJ7LwnxUGD9/0DfWSUMDDyS7
3T4TcVoJF6QgVQSfURKyXFWNrNBegUNANlMKGdAoSzAiynfjgDBC3j57HbB7
UUuJQmmxTjyRyQhBx+6V4qRaGz2RurdMYY2MFvbRjBDaa9Ngl9spTZD1O5OB
S89IzdrHnIz0eclLNmhG22UMb2TUkzXTS6tnG2UTp9ZkuNCatY0YN+vgNjtf
1K9Zwt+sZfEAUg9UScjia71b+/N175qBRUNgn8zCp9KADbpcn3HdiF8WIA05
dtwbl6Lw7qF3d91rD2Y3lOudbgCiFDXW0oTeAv/HEYoOfVxurrAqy2Ipwy1i
Sun4VFUapCR/PcX/nkdJl7CZyNQybi/l8IYvWWuEGkXHe8/zex4gRrQNaiRT
VW1PLwS9rQQFLuShn6dX7csqDDCR3IIUis7DcOTBnfRbaeiUCi9lFYSX759b
70b8ButMKenZ+yy4nDTcD6bsJ+tpOwxz2qbNELgDABbRnZWFRDdPxTE/wre8
y5rK+ocW5Z0vZtiO1SaIEtL+dxk2i5paYD9wl/t1LAnkLOUxkQU4rjwmaQk6
m8jHTs4Z/p27fyeQNrpNFx9/TckQsww87BZymdu5VzERQWAaaS5sq8aSLtS8
SDfaFuMXKCsmBe5Pm2Vi9EjMYuvxKKBUKxyJp7qD2Z7gGvVAyiDACdwNoR1o
7L22P24M8lwVmMFBKMQsBbVH0aQYnBFs7M01M5VugfktJhUZURdU0okPFcCh
s76Ef+3C4m6ihQ7FMlHh5dAqpb3n2aKRXMTeRRghUvhMMMqxbG0a5w62R3yS
PS8xeZpJly+UEnjpZKnQV7wSKpc2tJi8uR2VFoMFC9+EjubPgICOAxWQH7zD
3gUtiyqeGcdGk5QaK7Y3o9hdOT5ePCZiGHDkE0FwHzSFj2m/QUdX1dMIZo+o
trT4wkNOKL5oaROr9z5RTduQNnm/MR4wSGOHZZm1DoQCdfAr7PASDhnJ/ky2
TMzuXm1LJQCa/y4+w7pWFjECRCwizSE202jGLLAUmpv4Sg+EPU9jycckK2yb
BrfpjP59Mnq3DT0trznzZGNq92/hdo9R2cgBa3YKfhZ/YDmbASFBgVflIzFZ
uwtyGNKawIkA2nphya88sWA6UZ2OsmY1+gYykWvv9XK5hBEvDp2v952J0UpZ
IU8tf99lHqdsmiXZw04JEqtD0VgC8Rg0cWUSVhSnOJ6TSu7gJaBlmNhHR6xr
zffWPzlrM/1GLghXSgKNEQziBrl0geJtu2fKrMeyVHXK/V7DRcsBDoyXY+kQ
y8w5yZQyxLqKuVYpfhEH0e/n9wRZWW7Hu0txCVBu4JCVk2kgnYaR7brPaXUj
tDnkMyKyfW937vad1ur5DzvztCIiNpTrwr7rhkkBSvKq4B6LHnoh77GQx+E9
u0bn3/BYrna3D29bworA1kYeEDF143p4LFHmm6L0/ACWHE2r+C+DHahVr700
ER1n+L35rPRytccaSUmOCS5TVadkp28vLGwZNffZOUI9QAAs6Li66rslTP95
+DPT6SlsxPMTH2+JF1z/aEIzg2PeOBe2K51x1k3uBMP92gxxgoZCd6dOFkNM
zCrGxU/gNrp0Ek77ZlO/ySb3RnmG/+ov6kKmVlLa0dKCX95LHpzm3M2bq2qF
Mg6Y8u4fu207qD2raJTEHJV3B9OKLhHFzuLvOvv2X9QCjwU8yiWb7gge8DFK
JXc9h+7SAXRqfP+uG6MlwVgd2fw7AQlVVJ+3qjZzX9smT2Ac1olalReGeXzf
vGmQReEROS5hWPtKcB4Pwz5/RyjEFzHYjig4sTlUKwtkL3PbVTdLyI9TwkC8
frDA2TIvtBgKim59p+uvQoFbLKIh/XZI9zSdOrMdJ5CKC2WraZ3b14yRHf7Z
p+2vz1h4uB8XvRdMUbmPTBMx2Fu6WLRu6E8DTR97fHSlJYgmphZeHSiU0xSl
rxzVXNyQCKMDhW09LuaXNiF0e51W4y5bCzkaQRV00EAr7ZFOM6ZAhSIH9xeN
v5+T2oE1HjZTnv24Irvuq12KpAWx0xK+ZEVx/blD0UdUR71MM+c6TmzRRDLi
POIARhLOGn5uIC8zRMc4W5Z5LXTGXtAVBESX2eOMQ5I2u7vg2L/tH3TfsAoL
/1s8YeQFXNsIRGfCvSeTKFj1SRVm7MBjKc/r1wdU7V0Wo6n4e+NE+62oBQi+
DFyvj9qxaFoAcxmuMAdw9zqs5PQbI4LNtuzt+CEQblrTrerivXE6GqXobTTz
fnfMA8buxLsyGFpHbtje6VTC85cB7HSZwdAysxZ6za2kldbQNGEszka5ml+F
J61kvMLW0KVJRhuQtiFWsdzyWZXcIFLb5vxR+lusYlflH9BHMUvMSgqsBNmo
QZdE/wkzULOcIIbcSwMQRE3G/tMktpuXF2B8EvMP7Lw0UYyt6HQezv+etKkv
z+nR+EC5nQIzLNlAkijjOtGJ1x/mV6WLsmu7HWy8P/ci/ouvUa/P6bFoGM/E
6pRa8wN180k3WJfGPM4NWOVyAGH0bXZyoQ2MePDYqDl7GzVwzYho+9zdvJVK
GEJO9lR+UXroeGQL/KTgvzCaBgZGk1KjhaHnEK5Wi3Dtu7qY4P5W1Zw0G5o1
emuGSEifKjpGiCIq5wCvfVge/VVwNWr9o3PSKqPL9LyyKJTeWpx37AFf/ik8
6cYESOyNivgmE/uAOHceVyni+oXEjSUQ3SqQUtaOSigNO0PJiSW7pw2D8AAP
8tAqqVSRTgFYvP4B6Te7hMnC1iXZIW0qRhLg69i2LYvZF1Wt8eYjTdC9Btan
Xp9swBWW6Lh2f9Xx8oXwLrE3Ph03qKfK+JzuBmzeRPMKVNroqt4/508zhuRz
unZ/aKpvL+oS2jm9YG3RXvVA+lvaYuHLC8j3/REBbPgoCZU+xpFVRXzXiudE
kS1AgrlrO/ruHHz29RnoAYh3VUr346rtiU7GvrnCRmfYESK8YL16u+0Z2idl
mmXRi8aKZgTgiZ1PpK2Bspth5Tqv8hrPXkRL9/o4QcXBSo/xtnBRbe53KzXJ
G0N0zJjfB7wyScfaSGUIb7FKtfJ+EsyCNxjN75kTQGzjzH/RXloY1QR2SOKU
kiSupAT2gVktkdjWDYk9TtzEDx9xPhf71s/2KDnXd8jRVM6EnTA+/9vKnYUO
nHAGK8pEhyis6gkKf7oZ6lSvNAT64hEUndJLNZ9WwiO1NmIb9xjIyGW9vHYz
Ht8fmomTK3mCmwOSp9XnGbk+qMv0qjdDU+6t3fCa0Kgk9OBlhOpliCTsH7LQ
UcWW3f+3eJA3fzeqi/MFdyifN4Jqx+4Iopfyq7Sq+ldis3h3lHZbLFZ5XCHB
qaYw5svnMBsbHeRoqZP2s5II09/UOU+ohRkHpjADPg43vZRCTSqhg2/86Cab
wGKY+rhVJLmZuq7A7fbjo//Re3iuSnOFPoRleZs/0grrSeDWkJ5Vrs+X21i/
PiFVjDjRiv2T/s7g8LPp+Y+DP9iprI7Rjlngqpuzb1q8Zbd2lSW9J/dg0QXi
hxa+QQ/uhRgJV9igrpaETU/7Dda8wjSFMFmtQzTa/IdgoKAMfc4dIA12+n7c
3jP+UdWTpBXHKJB7lCsJt3hcg6Rr6jELyqBimTb8zW7aOXSJuN0+5hA1x2Bc
LOLZepiqD8q0LU8bf6CcoGalCPEBfeiRo+1ziRbfWE/vDrRswiVp8o1A3RGb
8BfUvKZK7nhqQzQbvBQUJKd88r0UT2IAxEeUQVUhEhwZ4/ep9PH4+WwtFCfD
mW+VQiPMDQ4Hea7mYlHrAkLq2FbGE6NS8Up27ExHwTXUimUcixbmXkERPleT
mLbmA9i7NR5bBupNOeeaY3ieD4yRv1o7G8mHn79w4XLKON+xkNYETjphLD6W
3A2ovRdrU5wo8he8oCsjux1Eo4gsX87xR6cu/oKGECxiqvNWgaBD/PYPlBam
7ouvuz21D0NijApUE38lPrTIZgRfFRZbuEhQ5oC5xVMbtXUn/qTH3ZY3FKBS
gpk/Gicf9lCeh9jXJVR3n2X79whCvXzFQZNXpDisftEL1A2pUV3y++RUM1bd
IhIdh5INOYur6UO9FzYH1uGwCEYLCPPI3VfLlcUGPvQargatbcLx/UeVyvWz
ED3QdAJ5hHJ/F2bQynN8WSP3BcdWcEqxrLdFZ83k7MPX3O+623BJ3E2GUpo3
bCHLbURYZlZ77kmJ7G/+GE5FokoSKYdb0BJDWYJiDQwbbY0bAesNnQPEOaH1
+bO7tibTB20anOJGPLwSSig6eZCUcZ7wH2qEAKBvdp7GCVHGnOoWlDZ+7zhO
MEs7OxDczJ+5EXJv+c0Eq25xWEGEg0R4A62tgNqgxqVm4Vh1WeiZun7rgu5H
Sai139euy6HMqKcvqNy6Tn72IlSVNZC2+ns16JbYBLMwSOP92ufhHrBn7X8s
uxyZkCE30Z0SssfEMrZ5WaQW1/AL5NaYQID5Ugsmmio/k5/hA95+wh2GujTF
QIwxItF+EkGEAWE5BVZOfm6v3Sd4KtnBSns/amnYVwwcb/6CjJXtiSxo9/6p
aKZYLHuBTyPNH4z6AoFpMKZcjyChaJwGETbF5/u8tGFAkuloKJaYtW/Gf6Hg
ZYEZ+xdDoPN8ITGvppIAPylAeVYueGiFWECW67Kf66y6X8r/A0SK2Xu3qgEd
Xod0dNnOnGzTE8CmDEbnuyIow90m7JqBl71U+t7ECAn70CUJx6uD103wrN0D
EzFS2VLHBVht08QYTTLnodrAo9NEr4+Xc063sU5Z26vsQtd4ZrQYS80Qei4E
84xgf/PZ2LMLXH8nulG92c2tFIC6TglBjw9hknZk+VCj5q09zCYB0e2/DgMs
wf2/iSFFK1naH6UaXdu+czDg4BDc6fzxzxRtcJpijXGw/Z5vQ1sagqCYLR6Z
mbwqwq+WTHs+j3XdWjpXIPG85vSTN9SuHz4h7SU0YvF+ly6XIlvnuApZuS7x
lAyVH/Wstz22XIxnZKldxBhi6YeJRMcMsLwjqeUb9coLOBUO12fyjpF44bCS
nY02FFoLrp4H3lQ8vTrXFKOj5Whbg6eCFJ4qfUAto9MVCjMJx7PM6TrwBirr
MXqBJW/tygRuBUm/oKwGFzJQn4QLpj2D+XLwnpqC9LKvvIddKpTbRRUrb8cE
RyaaZDyx0KtQHLCI/oPX7A0nikJmLR8mE12MP+ZZizvwtzLh+KN0bKNs8v2e
eBse7uD5rbsDvN9MZdMVHE1VRuzHBvBkOvqZnGXky1A3+/EXKWzSyj9lQKJw
qnZ83H2eFI3L9d2hhEGnbC+K7Al3ewxR+lEjtwNeZvKkiV9V6dKj14g/QQNS
aXVj4CwgCsubfA/yxuSxoxC3nb5QSokMe5rniUsDGfPd4moMgh7mMmdpWwF2
gccqZLPPzzASnjw9HQbFNTTK1MPQXjvt96lMY7OxVFrnzNyL/RfFaKKaKfoz
XmKOf8hk4+90lhywP+897MfhKYv4W7FsDFjJGX2+dA0KqXk2Gv5DHhpo0dkk
oWMbLeng70mftQWppjDu3fxzgklRGE2Cnl9HPnF1KXTee1tUzbZueQVvydfH
Pw80iaMsJhzM0UuugL9OKK/05fdutjwxMjpBX7/Z7Rs0i2gbJTxnUBwhxisi
XpSDpknP5y+t7b5tsvHLaY88kghTW4N2o4hhBGV4oNItJgYb9Z5vM8Erc0HW
19lDzv3qE9EN4lAOhcIcsHm9YlZ3uAcvCbF9I2ihWOlIvG8t98fguaBZgKM7
58o4IiyWgZkOqCTkNjzpcff0Lny2XsiZgJaFLs7JPawC1bobJsY0FZMJj0Yl
Z6BYKTuA0EGxb4Joz+R2jC+y5WnQGX+zyHAS7m/OOl5WerkZpRLaaoC97WKX
kuTVsND+MBNPru6IOEJzZMCNY2wCQeA+0xepsYcTGLxjK7kX5IrXZjjTAei/
7FMR6SlfgAxO5KyC3e4xaazzjxxpx2DtzNzXHUdmNiEu4SRU3CmagwM4Evaj
1dhdDZeIdmHrBVu7i3NjCRbBJUQGhYif0FrJefxblJME/euXuo33sV4i0pWy
w/hF1O8Vxft361Usy6kaTxeBXrLi6RUCO1p2SVgtAIKPJu88VXexcOIsdosb
wmG1a64+ZfHwi4IdnPgYngfjmqFwzBXAevfoPoPAekmTt/M+lhmw7wMNvDt1
QrKXkc0BkCpCd5idy06AGeFSUCDgafdhPFGIvi/mlhOa0A8Ua3C9i1Oztn+9
bag80Sv2q/X392wDxj5qzjW9WfrY4usplU+1aIY14AANI+0wFdu2NtaJmmJC
zyL5oxuwfdAYsKHF00LS7DTyUuThnmj3JvJ7PwlwukSeA7Ds6lRNjj2FzI+5
lGphO/g0MgV/HzmVHH2res58jaewFxR1l4sNMQFwhe4OOpznzddrWrX5c0IT
DKAXAlopuJfoBtjWJwqC2+Pwozn6dEPZNeJNrax+W87efqALnErABWaYuG3R
yS0NIKBL+AYDnrsQBvnx0xUTlM450N+AS87t6pvA5Aw5hO7j+7DeD+G10dqe
sR+otQYzgEAuNwEA0aOTr/A51WjX85rGfrzS7cMscUX09NaCumMUvNuVZYPN
BK4EV+54PgnLSZyIPOyGLzGN8qZaySoF/tZB9dw1uWoc8jXdzlU3585Zsuev
XxxV9RvqNH9ADIRQPDx91iUIRvGBwzmnxYMh29DgtskFb//lzRbmEFZFsbHh
acQXglfM7vNKXXMrrwjvyvV+f1ycmFVIrB7Cq1zTPFvOa7ld/UT26tr1aeX4
+UkrsPBiwMBZYGG79qZGM2DM2ZrLULLep5113jvKwXmTUH1NOaGd0UPeiaJd
fb/1wLhMnAOMIZRm4DETXasEvsGhLPkP6/2iYE5rm4J4UFSnJDNLtQr14Mh6
q5fjhihMsXQI16tmGSO2RvJqemMC40lIpOuzymplQF6yJ+l+C/jr55s2I5i5
sCaMrj7jGRU6xrpmAfy9bARTUQ0bFiZzPxYAAw2dhWPhwEmNqZgHXKg01esP
PnGiwvE4tTfnJ+t2Ip+MoChuNmKxut557qf8W7102WVi4VTOtwK1qLRfJ5oP
zsEgNV9hv9DzWUeqGVjtbZl98dXL0cMNT0Fk19YzkWfAMw1/LHsjlOhzDL2H
nhXeyzSm252JlbotSdpp1tbzpoiADYrrX9RKRPJfVWhvOh74szKUsYkDmrX0
RoignWX1XoYTq97N98sPuRHajYV7OHp9hIZVrJ3fI79f9abfiYZRdX3mBoAq
QkIs3z3swAKJwweELiTtvATE9p0wELFwtUyEobiBGEiD8+gk96bQECfoyQtY
IYTwdpBK8ws0tIDaScScin77rHujSuHXOw9oPVPlj5CvTAPfnP9NmAHHWVpf
qxtEIQP9AQcwSg8VKaN3DjHq8k8HXzXToq80kvTwrwjg/gwxvCW35IldISN2
/LmReUtqLGnQPeCR5r4MSBC1ttQPyezYN4XylT6pC4gBUf33sVwwBElrCLw4
b+rwqrY39HvyuPrjlQlspshN8s9lWardAbxvLsRPfgLS6YqEHi88CPk2eVYJ
Vmco/h0nGnSJnCfd5FEpijNm3N16J2HFvCaaHAh4uapBg77o5aQhBUNqPg+H
fuJsUCQK7F6r7xMZ+cQlLZOjvvoOPspu6NUvc2RJscCN4E4Et2CmSaxplHU1
YPfEO8UQ5YnBbBBbV/Em9H76Jz56zMqoHBzPvftMby1T7kQVoGyWrDA1A9C6
l34UWNpr9tg3y2IiMdoMc0WQIXKCDIjBQY96T5ZUgDI5Ufg5Dd1sdn/aktEy
mGZjWBFKnd2KLUCNVRzyRGkZe/zQUbUTobr0bazCc+OdCv2P0FceBaMWNaqP
+xHxBMmOczFo186AvCH2eWvWeNZ+lG6MWPDC3k5JtGoCt/rHcqWHGa92Mpp2
ghDGKJbB7W+ZhqhQ/f/uK93VCgwh9GIv6Eu4H4oav5ciqtgSmYN+1ILrJNOs
oHFmTluF0MT7m3ZSjPrLvj5hrLRZwdAyZ+sz7aW5oEiE31/twNI0JfClpzCd
io55YXFB5UmLc7UbuMsEy4jzRqhHidInwxCH7XNxLOKimigCmTOFbPZtkYmv
HD5TepW0Cw7q41woxaCinFcNa7GaNZ1CZd6TQ0kYImYaLtBgYtDGMqq7AXS6
lH55J1/a11Jxs2wXvIPR6PUdY3dd15i4CuX9EUSyBdhpKUWsKZgftxNKm4Ab
JK+bhY7W8FD0BAHWWJgk1ImTdJyy9o+T6CcDfgYZdoABkcsI/T7IFG+Zne5L
3NpVet9t4NEP4OJo/jD/O6B3Ug7/x3Hlsv/Xvz1LAzDRm6/zxZ6wblycgLGH
Uve74qfLohwWrqf6BdMEzziPevHOZCfKTfhEN7SoRcQGgUtC5V6cr8rC8KYJ
0G8cshZwshtIH5Srd+KSsCwtqxpA8GxSXgzAEnKI7uoxFuwJelLYgrBWPBa9
4Mzu2/l1C8aeNqtgOiv3RXql772tvFuRHLGH2XhgcyF7m71aBHhSLwJdiUFD
ZuF9rw3GrP7su5DaqpjjaiSWGbWwYQnLCQeK3j/+Vn9Mb0fZlmMxYeE5sDpk
tdoBjxd3JqvnYYoks3tL44naE1Wi6Kj8pBgienElW7H7YaEurEBLsTA0MHuO
Znhi9XXFzCu3s4dcbI+JDet/odxi3NR4i9CwNOn3CrPhkVc/03THyfyK4Df6
CnB/1ciAVk9QJeeFRAJkddB3mg952C3APD55X7IfJMNWjEyB1fweDeGlFV1C
Tnp3Jgqs50D9fVb+u5SKhMBvaWHB3Mb/dQW6Vv+dooVc/youUl6GQ1CANU8v
4iuA5khffsLyWtomwzb93071WOVoeA+rMLCbtrILm6DQmrJXi4Uu8gPQ5Tmw
B1nfHDAZ61v+Y5B7TTilQKL2fPStskzcWcrJ4ZxAwAIrDUFbWeqmJV8jExW7
YZbGyJ4LZjlJC81o15joBHCc9cC95u01gzeOkKoIGulvd3rDAQ5AcBM4bUCj
UrYbA6O4aniq6zlP3gya5gUf9tTzbYoyvU5et1eMIA1RkOZo873SjeIaHbo4
MFSRuvR0CHorfAjYjE8igznzWbJdTUPwBuF6oldFBaqhUBFIBFM0e1u5/h2c
ACQ7LfAl+o3T6wL48SGHK3nsNnkM40yTd6vMRpbyMcZnZ8uDxdek8zGtMDwP
nJALNtf7NxMb56bB4UBsgIq8JT3Lib+RKemIgOFeClRCZ5PIO3MMRLebZmjW
CDcPHUawEHgU30mYgpotPUbWIWy2vSqhDPnSnlrj4bKKYhIHmPi1oE+2ZHFE
hr1Ig/gLs+nRkS/0hzlm/wg3u5pcgIAhKwducn9W9GtZxv6WCLAjCdY1L1Zp
PWWAz8jNdI90AlR71VOmdQ8ykT8bRNGcO/HZ/pnMtCQS23CJ5jt4mPOX+jJq
kegLEXSD37Gz2MBUcdcGl9lPfUrilJthSwX3yThpv1wVbbGnC44LkkpyJPaj
CXyW3n1g/Kpvei7oLOlO8bzFKl/41Fr0kaQpToPryT+wLmzOdv/1OM313Whg
8udm1GbHPNQKvAvSSWSHDmpXopd2Az25SWLwl8qYipw4399CPFEVMENPqUWG
tXhGl+hLb5y0dSSgvupA7foV4Ws50eohm8jucP2dfaypFJ6NsZGHJQWYXHWD
0Vdf8HmIaSfcazuY3FRrnrFJ1mzIywE6oFxz6x2yXwPQXGECVlm0w59rBsSm
CZkBZfOixPsf2n2xZCh727+mJEix+PlLwPEE8MtLxhJORRi4aUBiFEaxXPST
SVscBYOS8dkXPAByfxQKZcgsEldU2NFno4gA5qpcogyNsX6dcJbdA+9Npo8m
g48s5gcUzWUibKtQI9H1k+jPetEpOK4YJO3WeqcB7SyxelfbyG/eZJWle1Ii
Fx6teKKghdd4PIdze5mhU3cSZkXFkxLmmRr2tUIIrhYOQBxSbM4lxqdhwmeX
eNT6uBDsGqCwODCC1U9nCksUYfKVxzj9mkFGxHUokq4CWWi1lrM9EBZjJZsb
yP5gg9QMq7+ctcJJcHOvQEJJYsREWeLG4c1dfMek978FEUOn590xcTNn/zff
EAZ37Zkx609wVxNvTaJtadX7vLMjnY1dsauHCJ8+OKSqD9OOQLJA31J9uDe+
h/+SOBdxrX8N7wHKxMp+q3w4Evb8w3SWsxnrOXqcEofM7WfdJj9vWJwQtDRC
bRkvHv8mAxJnKQmfawLZg9huQl1Nv98MqCXBRuGY74MRstWYTGnbcAdJium9
vGFVbvK/9nJEURykLVwKcZS4QpUbIxQGL8Bt+i1qZLyJLO6VSOJDVmebTQgS
hqTUnShNNoKY9CU1KTFDMlxVE8z9+wp+gEQfrQGQYMDLcTpNDus+ZbbRld84
pfoYutEDAD12/JtVg3U+j7wI9xyl2TD7VMeKT9tV4OpEzAY2brE94hTeAGGt
yglMd6VTq5mCwgmi02hQ2sHP5XHkqqlFxEoX2tS1+l0TmM2nMZ2IqbgPuQ9h
btyEy7V4h1AqGTnUhAA2ujrbHX94CiQmMO+vwh2RK/q6wliy2LsXMo/VfslE
umX0WA8JqHCiSJVDWbnS8UiNOVBoUYBQaMUn+DfsQe3bFuue6JcJszEHsHe4
3vnyOJ2smJWL/3rR1K33SMyQzkR1w5ILs1kRZDByJIoCakvNunKG5WHxKT4j
lCNvNE+jko+qF6NgEfT6CEgKdEWbodPEIiiwtkOJLt5ymsvvtYg+LRWebLWP
yT4+txNyZwfDgRfa4rKgQw/NZeglsMiVzWnCfDmdKKMb1T9C3rZKhBIA8TDa
j58sNyMgyzjMu0J/VUWPPxpgddyn21KWTJoJKEncf3UDzEdIj6xsnE2ryIDa
ccA7yX+d5Wjn1njgWVvwjU1N+U7Z1wEVqGvJqZGSrCruDX4kDbnYV61FNnOZ
VFlde+OwHWjOiTpgAkGWDvrck+M4GslJrsG8X4AbD0PEt4rAGpDcd5PyuIiS
x+4igwpvK6zWsN+jxxa6GMvaMmYrtJqC7nQRBHnZZzF28tgYQkALkKtH8ff9
asA6BlLctqB0SC5/ltJmOzYbV1dVPHrGbInvuRr8h3aR4ZbKiPtGtrFInIMJ
wnJkoZAmHhl19aa3Ti+A5M4Ncfd9GcDWxS9D3h9ADiPEyJonjWeRbOE7EZnd
9OCXolh8ZvT/IHqTb2UlhgY/Y2thOfMWvSbpGI8pJ3iIGTbJ5T4z/abcRmvP
hpPjbzqYcr1Eii+vOUEwR/LjLon48KcDm7OaCyW1eqJl6hHHxp22ODhvjVJd
ADvQqN6fEi8hEhF2ZCN/5Nb4ahUjf3fmiA5U8MNJR171T/oDtSspP/BwOGM1
kb73am44MWL689o/ZkDqe7Rh2dUxKS2z+UO0cqx4u4vXCvJTSkc1Q/DfdtVc
JEmFpPq69VkqQZ7p0Z3UyRAsXUpXDr7RR1HpXyhih0y8vin4zp3cEq6/1F5a
kCRGbhdfwQKLVC3IpeDwlLMdk9MLXSCif1wr4mntLey4ny+DK/ARkuaqUZxK
5Du3TaYdS6xDgkXGk2pxNFrB+r4irCudrNmlGhocbTtNf6uIZ2SWJBRpmShr
gaybudmCqtytGSWk+gmqqWAOZmIDZ2zkqn6fMCZtXSx/JFjjDoNN56dK0zL2
VA/AyvPT02hP5P1W558m+mX3kb7S6awFaexlt9k9A8QXvJqVYNbIoKUX41Om
c/evbfrlPfFPf1HouGh13isabYRa+lZ4GDfg/wqbto5s/ra7uiV46VvWWeb/
aD0EmQ4C2+hVSR8tbLGYm1cUY0NRZ98B80ZCXcyMhHlfu4zhhQiN1+WcitaA
nbxbiuekp2jggzy2Lq0/ZQcgpRU7rljaJNKzD6y4AmjgdgY6fT4DeQ8x3eu/
E0+ZmqQO3HJ5wXhx376oy+/hmlpVhQHGs5wslBIvQDTCydPythGZsikcOCqh
SopEwzHKd+p+sKzKWR1D4bP1TmOC9XD6GVD6xGxF24SSCQIO90czyg9WTN/i
5hFSTmHTItR7cnIWKXdoGAkvNTzTGDnBRjH5+V4jOqdk4RyKiSbaj9ppHMBR
lCrB1OD7VNk0RLaVGZiqZllNUMCU/JS1Yt9raswcZz3F3gUVbcE+o60Bl7VJ
jkbnsqJgINrn66HQ47PuJWoTLJuOttZZUMqyn8vpMGUqYQJecBrQvAShz5hF
W4beoRASAN/Hm+SEgX0mv7KLKznyiOpNzMyeW1LPdmOd1iBrryuhqXTPYLA2
hYMbi+J22GAJwHMsagXy9ztB5Hmls7pfy2gIYYgTWatDgLBkm6oc/UjbdAAm
g6jJhp2qxcSliD0Y6vl32NZoIeXtDguoG2+7w+I5FdUHynRdlpylsJUhumBg
Aee0aiUMuHjU7WlYROlSspr1oBfCV1DPnCa4hVQECX94pYl7GlWHCBYtjN/4
cK/QPNJAA32ynl7uqALkNf3I5e/f0gWWe0yZqAQwiXJC2iOoC8Xizcrads6k
1BV5bFLN7Xs7QFzPAR+1u05TkEj67i9MlZRLRSQF7i12kWTDCNb73NB75OJi
SkpMuU8m6NpAtY4xhrM3m5AFZqEk1XPQ5PzUbnt5/Jmn5EFFbQuFbHUG5yjN
rvSJtXmNv90PaWbbivmkYA8DZSnabRNTOh1r/fNMq6kqy8myJr1zvrhDaTCg
VpwGOaZlQYiK07qym2Vwm+O3mxoLFikuqOogBHVZviaOiWy8DjPOPQKlzdT9
TzQMGv5n+PkZmzPyuD325YT7WyKD9GKqcHPRwbriWtZULMok0Su5d6PEJl5G
9y9OAvueCLNu8vhkezJF6/M6swjOhnjtJlMJh7YCOG64IZ7PxkgmvxtoyeNH
CibaeVoUSKStafbr9vT01sEb2i/jqf+Ai6MOBDDJdbf0kdl1N4DoyErHtDm+
Mm91YOZ906n8Lz67QOgAiKBPaB7+/a1+LlVS+BuspsUb42ANXbu8rZxA6juf
CyD2nIpHjCcR+KKbNT9mNMqpgMWblkTEuQ+bB2t0oiMUFC21/2QbusGzexYV
AlJg1LgdOu/lmDargItWxkfwiZAHLPAUvYfNBxEnojP0BWVNDfU2g+OZpAty
VE6nWlCBTt9sUe1I4b0bqHjDQeQFeb7wxQjobxYInj46bNzpFLGaxqi8ZlKB
2vPnqwpabY23/CYSyHlTNji89PETMk74giEx0/ioz0cghuTcF1hMc1pXPdip
zz9j0jqnEJsh67sHDBxRq9B3FEcnp67bXHTNh9oAJBRDaFwmL6J8s+o6Olrx
fscByTwHRLrhZkxLunH94fgTBH93qthhCw2i/2eyO2x8NIa2iVugDyOHmgbG
j7mp/3pwranb0WLP6KL1DOFpRJM62NU3Bbb9KBpVR8YfkntPGubUIC+7Jhbr
8iCbl45KMoAVuUmyaIGajLcLIarkdEPljuD2uS19fOZf57g0UEQXqgfRXCnG
63xT0x5d9UhqGei0ojPuI6jkmAWiFcJdXE4og0cOTdXpmxfhMzdvWidbElKy
v71oJYZiXylGpAOuD2m7DjsQuApOwOiXh26w2t/40SWjSy/ZSrwMTcXznY/7
ZkAgol0Nf6Y4QoeVmio5+EBMLIt5pMDyo0rw1GYSus8S6fQfWx/tiSJnsv7i
JrSfLWxSyrjrvjNEH/VhnsyataTYKa9FlW9HAcaMsKTkrlEkGdEmB428ZuhA
dIF0jf+wcsIBtbUuZRverf7V0jB8YTbKLiGqZRIqTkehGlmJmsQBpL3XiCf7
tR+sD5A2zie3wSz++hILioksp3CwjKWIPToPTS/cZIGCtN6MrP2qTs3dV4F6
01l7F498r3DM7y12ORm4ERzXCfkUtHM66kkoUwAspRNSINPMJjfw9lAovLyg
IbwJcFTMz+OzYY97CRx3qYU7BT80kGjUFPn4qodOJ2kM2FSHUiC2CfhqnOcJ
G/cmL2xOvDmcY2bQ0wYmxo5oFfkuLYovl4CEl2ERZhnJztOxOtHsHnK8myA5
zQ+WKcuT6UHO92AplJWWTx2mUr6EY092ghZGV4bMjjhaktWwtpObbb47J1iZ
Lw7gsSBgAd+QUrh1XCJAnf/kc/UaFpJs83r75hvOPv46MFJQ0LyhYOigSvvI
30UAVPYTSNUl4JuMGVs4RMIF/+vA4f8WFtP9pyLvodLyC9WTwn4Rl8Js4SP6
cviPfGsbPm8+49qS9z6/Y1VFRjr4DTC5RLca0ws1oMacVJ5OI6H5GLc0RsQI
MG4Guqot0ITh+i3+CMf4gxu6ltKhxDNPDG33lMH3g/GoLCXAiD8RvroNBSo7
0SOuyZnN5X6bxsOG9EIDfiYMhYHtau68ZkwdNtdSggYdvaix2a4o3BSn9Mmw
xETuUdy+MAC6tMuqphUN930qDPh16zG49Hij5vAXN4MCi2/KxV8mqmhTP1IO
+pNaBR6cd/PownHv5pKBlJt3PueOLBNOwYkOSLh4L3J7LB5fwDklh9ScX/If
wPkOvF31KoEw7SX+eOtb/xWQaCy7N65kChFRqAeALANQRVBFs56ECrKXhtVe
aq7Yi6afibX41xyBzy9Hm7qh7fhxtcR+t84gcrrQ+IbFhe/yoLrtTVdVj0ed
QKjEAu6fL4z9N5f7fz8IRhypNzqKrwlI7LolIYAHXyrB9BO7ArZNxRZCOi5+
vBqnfRXAqudkz/qZTJBvGbjHEWcj0X1ttAIUpolVllwS/+GDOGZcVeL9Gga2
RUNYI1r+tX6H5JD7iabVvY6/qIfg3m6HXDG2qPznz3VAVzeh5iLlaXyvaIlz
hWZkAUzNFPW4CViAv/9kXjX3SkpXYJ97DD2omvlq02xZNaa2QCl5NNqJfNsD
Mn/s0n3p/AEDsZp/nP6JU3L5g3IkiKwfzvQXe/7d7Mr76Vtc9dFgaA86eLM/
rif7NXoQsyhQRtrcVJNS8AAUN6DqPOIbJE0LbBFgZ+oSMQVr2EpZ3TYx8ssN
GnLI31hGAfJ6YMdcc6w2bYmq5gJgescDW/fijaGRDlIcVHx95pzN0p4Z2SPp
ld1ofT6Gg+6azzzZ2JjNjKXGQTNScKAGN3FVFn5Jkfh06a+aX4wQhi6w1Fas
ECRBiqAIDOb7p31k5ItwU691Xq74N5quc+hHXxK0MPHbozNqzm48RJaHt98l
w3pkpPxatb6MymdnXaQcwLYwygz9VIwQkRPyMFOxYL3EmuQIWEDnP5p/jtFh
CY+O+MRFqYIUcOOtfNteKF24xN/cfbbUxw6/RcWUHqHje0aPiABeAifGOnBc
0xsV+QrcLOQbvGEcSUy+Wor5/pmn99UqHoYq3O/iYC+JGMarq5Vj6VArf77j
XOQtvlfPOX+BB7HWHb9LRK7jHXrHMeXoSu+AxGl/Exx2wgFqMX05/2BZr6GK
fixnO5QpOwtxBRq/TzWPyc+BztuWS8OSgP8RxXWxUYdOl7QtrsBxJO881dYs
pKPoxK91ogcE8NhqxVo7zllpX7GzDhPQAFWPA9YI5EMMqZXT+fYyFolwIBqz
w8+pFGDGfXR5PPSpPRxcWMmqogwdIf6yk4qefeXmoK2hQSytNYPA4Wn0RaRP
2VGh6oQBavjZIPB0ub+H2ytf3VZrke1qu6paCi1zpY06kQpVlEK9kfP148Aj
CrWTCCCtGJNsUPAE5H6u/kfWUBVZVfM6b2+rWDnhD9lC/ncnD2M20JMbmkRP
jbOMbO90tn2ecaC2xB8jwAszXhmWJCDs1rtMwq2Xvb1lf1ro6dx7uKi5BZlp
Ngo1wkH1MBEFGQakEm0idzIU/pAwFdtiBXw4Nl1a/M1RFz16fZ9ohtFD2efc
oBoC6wGkDvNaGNgtwFCvruvR8lcUgIKRYq45b58/JaD8Hef49bMwkLVISBDq
kaT8aLRhYb0RQ/h9NC33rrdgsBVcftkXTkqQ+1ppuL1rWBtBIsfRLOSLtbqk
JUl2OxuI0jumnIm6aKk6/P/677Qe0+9Ml0PZzTMSCSDLCq4rkb5LHLGLdJ8w
hSEj/n5xcF0igSTT60f+CbHAvKrtzShX6Wk9zPXOvID/kf4QYnDBZNyK1XeO
iE8Qs3kG2zb3W6DrbkLvGPaibVVV/ucA2XuOM1Vjwv/Lu82HsCksqL4i8gEb
SUm07EMs1lzt/0LyU38527roqGHml4kKXZNt40S1T+RHslhk1v+/sOouTSCy
fdom2Vh6lGmhsLCIV9thN4PMUrRqDSIxIWqCMs5m19h5XGc0Lc71v26W1sKe
DXsl3jXxjPePMl8busgewlC8RpBQ/DG/kL6gqZqYIr2fGtYl9oPmM4G73I6A
lC40WHQZFzsRi5MSuWCo4frt+6Jxs+oLAf74JHWTaxU9b2OQ6eDQxWfSzsht
m9OA4DP2mZ+QRPRhOvUPN7GBJZgk8KG7T9B8vWubg3JgJCSSGFg4tuwH8sii
xOFKkW83Gu1OTexQgXCDubTfdqMRIJEGTCL17vd+yOxZCEQ6IIuQ8L8djIub
jsKUl0/EbtP4J8cUz4qy8J56RiQlQyjJ9qgJFB/dI4JAeFxt35q79JFb6EWx
VBJ/dh3oto5/uniOromWKZfV1MdXZ3B6+QD0vKmkpTov7kd8nh5Ut4a4R6aW
iGJ+PSpaMwOc0YlGdgPYrQOhdUyrS7p+dcOw7wd2BtYW54jGL6/yTajiB2Tn
uBOh/XkQDM5uK/ioowg3DGxHj4CmSmsTw7mCjmYKUeVGCuBef4qEJqt69slB
luURElEATd88KDdWIy/22N2nVf78KtqXrX8v/aMxRwbY3pAAbm7LrFRYpbxU
Dre1DuODRSQiQcX27jtE7xTPGYMP+mx/NEaM0/69Dk6xJzir/zy1+X/WEb8c
NmqHEtn8UruKWoSMWJH1BJAnFWSOottkwhfinxrOAyfbyl7FAQIgO6kASTe1
lgpUR8am5PWWb/9qRd71EJeUIE06dz9g28S9o+3PvTjzO1ckt5AAjBSDv/Oc
uAwJESVvxtZEGlS+usyvZS/dHP6GrGcRZ8D1qyHDF6FYmsD5yy3fcumUhrR9
AamM215p4+UC8h/02k7DZ5z7F2VHyZqgjM3VOUwXqH2T2ekyEoBM2huAfHTj
UgfMa9yiWQq0oUxAfdU9bsDJmkRVTNKc49S6xkXxo/3y8fK467moep/p/tha
lWMhCCxlCxabiJoRYnadHOvOCJk6dOb17OSi/juhdTyItHYOmv5/4IvwPDGf
v6qUBs+Dmsx5S3+U/a0FTjsAb42KCjKQXwJhXNBbIRqHVWgtt+vB9gBfSEYd
uxkdl79aioIXiDALNeKvX7JkXxZStGddidScU96eDTOPN1fcYPXESQuIFXX9
PIGBc/xDAYrUitg4GXrioLHUOIO8q/ia4sw+DWXm1uEKF+zLiuK+i4q00R2Q
wRJIoMH7wEw6SzkQu3j/TuBN

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfQ9KeyGj4CzpJU8CpD56MhjVMZwhZKNaRBc1oMGCWbIYkjEQgkqMJL6pjmfaqSOQj1kLvKkB4/ni4gwj+YEcPbyvNzwEwYk4BXf4o5mPyCIcs4dmAtVPbn0Fy/oclvMzSpzuQmnlgVsrG3nv09tiXcb7ZrESqPLzk6DwRPi/hG8PNtQKMdSLr1EuR8bdsw4ovSAGVfyWSu9pt2bxGTkx98iajLojw8axcm+yXcau0ntJlBeuOsN4tajkYo4BTi4UXlpc5aqhV6ORBOpjuDeL4Pk4q5+GAi2CMoNLS5XGECWcapHGP7cutuCDrlinBqC2WCg5s7Y6hJ87ZESOzhCDDB36MH6YqUdXje70AHD1s0bhVBF5Qo4/iecDL2hW/BX772bRUnmFFtUalfvxwmYzcE1mnN61dZT43UcnzDTaItZUW3qhziq+7NrZXXFmULoPlhdIWC5aQXvVl09kEVduZ4X4kQHtLRdsGhRWEngOC09XDj8ER7MtNIwjEn7UfbL4PeKbHIxVcVYkwNgIYkqaaZt/rQ90eCfodDwid2/leq02aq063b8/LhBQqn3VpCzFaka1/odmbCXmJp1YbQ4EYLAVtBTsXcKehNjsOv5oLr28jKIqYmko5xy+bJ0dJHMx5SeNps8q34RMAqeiG8gjzyBbRT34zBMDMY4Bn27zx/wkLWwl3yGE6ZMz/yQu8w7aVIlPjsBUzOuAYZoatOJ7XGWfjcWwZsibUm8y0RYlfEDO6n8CW7UHVr4nOWmuwzlcXqMgcrq7n7K5XSslUlBmV0k"
`endif