//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
r4sSL9cftiPh4OK869tzMO73VF9HINhfqw1yeQugiT3tVj7xKwhddZmqn7f/
lsIy1XETKsVyBjfSY2XAv2HLBdheesUIytpt1DJApxnK93N+pydhee0F+7zB
iKhFvH2joo9lWvwqEk96D2EiRYR71koE+qcTX3l8G6k7Z1dj580dsPLzsNh2
Ef2SGK97375REOnWuc7qTiJNCch8C5ZdA8OI4xKNcwALDifMjz8RhiV/KXeY
KPiMy6U4+ZTUIYx/f5b5/wOVqYQNcOIRoX+xo3Sn/pAgveLFZ94YO8gAesb4
NFhzhhMEWtVWUN6grVaes2tqJbU6FSQvLEeJt5PGlw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nwCxZ07bbsrEKcwv4k+inXFRP1rQHEIXksY8wN/y8EYu9LDDR9rUxavjWmQu
DJx4EKTCy6Tlzv4fxa08UhYnvmxNcDBponuKgzr5A/FBeVlAy3FjjFrexK83
GEN6upLjuVzssGqIUzzn/kUX52/Lx8Mqv3QAYHUdtmxJGnw6ko7xfGvX0EQ7
Y3LQkbPdIrQnBFjlCDJWGTNBHwgddmlbeRW12YT/WRFRlfur6MZMTtkvzB/v
qZplxc4yhBRWk94OJkofSN6j7XzoTAq0B1hUaqhUz/kJxhdy/3qQaQqCHbs/
/cf+7sGfTcP8qBdHwj5xrPoyeJIeQzw7eMJD+LCxgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LdnmU1oPyh3j2CX8UsEbrxacGNNGIkEXQlp2hf6rdyhYOQSEIYRClR+UkncR
krAJ2GFRcO35o0l9BXRZwtmtkoNIMab5JjIA8ZlJ6fKuQA26FNs7aAoi+a50
cuv5R6s1rigVWsl9+HWqGYQPvPDfGMkv44KRMIPvQYOOyPQG30hTrSeBFetM
fcxQpDCa0oyz5ll27/w4sroRbUcVYxBqdwZCXXTSJxhnebjNWjVBnFR8knaj
47O77sEuHBiRnV4Uu7OnxpumjFP8FEQ3+Q2oA7bHtYFmuJYhmybX3Zh1UYSs
2HuLOtYJbZfVCeR32TGeXOPCdLmXwTv3avFcUzDIwA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XlHtWGjih7MbIKuX6P8IYbPhiMnsHQz3xXfS66oMHEQkijJDgPQqSdLXUXt6
zF8wuJ2DzrMu6+o1WnqPLB+/mvSoGlA/nJu/VCKiTizCII1fqRZgxAIZETLk
wvY833ZV5pEvhbodmavdQbs+UBAvvvIvtqTnAUEqeZCO4zkHfTk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
uFtb3up8j0H73ve4CdoCrInIr2n+f+F64IfU4eaWy+oQ9ohDRTU2TH//GS2e
H6xt3EQaKbrFoa3zJ3941XuaIB/p+1AGWddYx9W8Yy1dCw1WRXcPSGUZ+Fhe
Y18oj1CYzvbZA/FfEzJuwGPNOIMZ7ooAQcbWX9JT173/oZlEDXczwNAhCfjd
uf7DA7xLo3a76rmIco8KZIwQ75g3CU3dHxSqOP+ljfcW96QvdvMwGHkpI8b+
80piLmIWepb0NdDUbWJh5I6m6YiUMCbJ+rWO2ziiWqLEiESSgvA5k4pyZV5+
21AF7anbZlQ1oih4dm82BRkhv93gmS8bybb5KLdXTjsx9n1rWvy3ivT4S7sn
uuAyqkzdnhAvxrr+YXax4+2PGpDflbJJAyiqZSPEl1vYldgBV8Jn7rB/izGC
KnCULU5oi0II9xy7HCgckaa/nZE7Mvz53Px+GTVy3yTHQWO5JcnfPH9PPRfC
RlBmILw7HyJ6JnO4zaJQG+KrgpFEgPc6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ug9CzFpTfobpMC1Ae7lfQjHp7yUnlZH20tXufE2q2getqoTirND3QdD13BAi
e+SHKIjtF0Dcot37TGTwZr6Uytk3SVIN5yaKgfFyHwTqWC2bz8Rb0HgdpixS
KP5whfHiv9zH94D17IRWBDoUu20uOWxRtO4YrzyIHBb1i3VrWb4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JcVgNaaicxbEEVvdV1mUT89eK6Vju56q/KgsGdi5V4Q6W85ZhaMXlkJ4BCGE
4Dvr/VBurGwtrU+a3x1/Y8QxBD85LtkLyvbmKqOvxeTKnqzQ2KvbZ7jVdjWg
eTjsURaof+DgLJCzrI8sDh2Z/6C58Uu8aLEVf2iEOiadDAgu0Hc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10416)
`pragma protect data_block
ECiLhayB5IxSbiyxoXoKOfZKw78rzIxf3OpOyCj0WXgB/fYR5KDnZYOXAdV3
rrQ8w/LDGwaqWxx97UI9sH/1lMuYZVlr/iaGOC8xY8yY1Ogg5L6mFMBZDHHg
iNYYoz2IyCB2krOFD+8U/sGAvKm7YdKikr4A9zE8psBIDhjzpVec8eu0+3om
s+iCFSOcDPfX2O0kmC19+QG1PlgQtOy2DkhR/MMhb9nEpAlhB28vu3mfYdwu
/LdvP1Tq49FkcWe/EU8TGWSzo4EBv7EDUw4HYap26Sk616TZzFtvv0m1zzb/
mnnL6SD0VkZX4a8YLsxNYS4SpXBlo3GCgLCHlBCLQDNS5eK4xONt3S3vWZj+
X+pquIqvgy9mOxbbS7Aj0miv8sLfxy9IRrbh0CzWUaPSBtjeBAsq4Xrokf0i
soW+ZoSXCdbawNGOwJLOMKDWnpDsQ+q2uxDERCD7s+ZYM02BWHzRYjtmfaqt
q7LY8HfnIuly2tlgasE8IJbU2nrY75RcSZ+BqS9k3O1m9wFtVnsigjXQnbiT
iDZqrz19tahwBZgZhI2AgLue5mgf/Kax7/j57OdvHyy9hSCN71zQ5b3P2Sum
Dpy4i9kQPqxY5GxTgv6G0RewONqYry6M4yrrefZ3UDVjdXc0AZzCQ0SdxoNV
FDtyi7B1Eti1lh55zF9quvYfN3p87+hN3WM1cBu4meVnJoJNBkRfQ/YundOZ
ABiOgfNlSSQTk8qMnM/J6+zKHX+o7CNwTapawyiFiuFvyoKQ7hlO1fy4W56f
rxn1F034IPw+m3e/FgEBdAkf2KN7MIPRGim7RJc3O5U1Og/5eshwO05Y1VmG
FBZG4ek3TlIvw+nODF13li9BIWFmvbD8eVC5n3V19vZ4D/O83m/7HwvVTgKc
NupxJEYB1t04iePGBqqW0GzIgwDhiM781icxSS+ZPolUhw91b/SmRt6kZcsg
SVNWMH5VCnZRmV6mp1kJIl/kJqtskdvahe4Mh48c9vAq/iYXyK70Sf1qG4wY
gC5oL3Ykbn+YRmZh/bRsIMsLQkXnXrCNJZGAZwvD1w0rYqynQKFK9DXEds/R
N12VgIDl3nkmdGFLcrfY4ASoLXeLFIkxXY1g2rxZ/dyFVXNYhA6BH3ZTKU7C
vT5+USpPFnen97JCvj4hWUCLqGEZhRImR00F2fg0Ztc71Za3rDo651AKR79y
WTF3Iexrdzgyf9Au2I0uPUubslgGL9r/CZwIR3A8AbPMt2ETzuu8wt3PQuYp
fS2c1L9yIPqXFZlGwFB68XLcvIgQWL8H+kOkg3kRllaCw8dCK1ewp0NInjo+
eofaHmLqKuOc/nviRNN2m6l4uSIwNre3Z6d8eGbW2UbNu9muQsf5NQ+GwGye
mwGNBOUKWZtSKLjSjUYTzqt9UpbP0NrT4zCePjC7ibam/0ALeVfvACuceIRu
B0WU9wSjJTw7yijJFWHDmHPPzMSigc+2rk3a3z8BdumlGd4s0SJ/xwqwc8eE
GeKSd2N000XM3EzA6anfbyCxuDGQdDO728KWVclYjWVDxcbEiTPnvUm5IbRn
pLb+O2/0Ei826tzxw/5dtskbkrxKy41AhOHxBFE3I1QgWl2vN2xLTscEsG/7
OrtLB+yE7dX9L+r7kWEN75OJzyFqtJgTaFWhPw+3PKByndlMimz6NkvULvdL
4UfG203/FzMllM5W03d8s3re3PSi3V2K8g9NBsV+m6jO7deZCZw3Cybv6/Hm
yZuX/ZgkGuACFrww3rEI2OJIyOkVasvUPiiidxJXzgmauUCALCt36Hucz0+O
8zlyCrwrDsGig3+hUHpAmtxBX1MHzc0nMZwI6NksosaD2pqwNbVhbg2ywVg6
eS6+5cVfrQtNewofD0AvJIqLsY6Y8gu6cYtQjA7CfNKpZoWPuA3+BMoRvaw8
oMVKK7IIqh33OLeqMXHVazK9wEC+VRO3UuGz8K3Lpr6x/+kM6PivFdGeuxGq
F71rC25rk7JHVr2BzaI2KCtTzlDr5vE0gFxZnXueCtRoq2xVgfKRLu9vqW6/
1LdM23XMxHhPBl60zoCP8jpl27hiAraBfuP7g9htWdTxiWPVzQUssXiURGr/
p0DXhTBnDvdxAV/7O2CofNMqnHqFjtvVA9xyY0h+DcWUQK9pmBjAsDn84vT2
kZMQD5xt79aTze4mYKaL2LlqSfjeVniNbH46/x+I/OssRosT/pZxwjXdEvnT
mx4/1lXado4wKfpMVWOrHvfFAeN6Oo37f4YWIhDY478RvxW+ql4X1uhwWQjG
wszt3z57a7q6FdZvDcR+b7RKcPjSJy820oNVy63ksNsUNj2D6sAHFQL04E+6
o93fequ+8pjJW9D0KA1GKISYxF7F7DFxslAVoqslDvRIjjiWaxoIQmpSxcjg
QG1wGL4NUapJQReimWyibLb5L7/JUgnwBUBHJXoM2Mx9EMA7x2Yi0qPq9mw9
Hmo8m9KLa3VKSvQeoqoXIkCXaWV0MLlcACyyiPbqzG7IbAY5PrKqYc5D6aku
GQBZDpCY8OUyo3zw3oos6Bei3Aoi5kQAK64QmtPD4jxNfRMVUFoNKfWIV000
Sa5ye0ftzbDSxOPAI7zuhAgVlsJL74XRPqzhDl9LqMKci/6jSqfzQwAq5tyD
sfFjSQH1+8Co3ua0uEgRlGbRNfhRaaD2yejEVIzMlPiZuo1qNvBgCu/y/bxl
8tWj+o4fy/ug6pE3s6iFSfyZL91uO3i3OdkWdKNv+SSBecV41RpyCwg98GWu
EUt0G3VlmBKnz0hzO2bmVApZdSjwzo5b05C556E4Q9RsyttE8I0LE3J6VpJH
ksOoGbKoNq9tBUBmMkB70y6tkGwB7SeWOwO2+HNSxoM6zSktu2OizYHxZJGc
7mCzwCJAjZzUB3c2jKPpEkF7RgTSxYFv/u8aHdmCoMdvMnlJkZyKgIpCj9Nu
+Np9pFQwjQByTE+iEwZRAdZRe7Dg5UW9ZJcND4CZZGco2/N0YTWzLPuC/WS4
R0+8Mak+RpuAFf7pFnnahXA5guETTI/pAHUReIE3hzeyyd16Eb0piXvItH6S
QXWisr8dPTITrvNb0uF0h5IhPvj+4juJvRQZnkTYNEeJP6+D7EKU2yMwZ3zB
m7FUGNv385M2Lxki5LHzk72SWL1QrGYRFnLW8L8dQacP/meglp4AsvnTya5b
WNWqfO8+XwhuMVSrn7gxcLHBtmx6SsjxKGNiaFgF9u+Y2bII2EJP/nvWgUeC
lPdIAE7pJ2Mg+LjyXcSkgz3XCi1VsiTJHkMWrhGy8ch1bN7oACE0yfgu6pZD
AGT8O+6/qMEO2zHTOsgW/ogWYnrkokah7lmxQuWNNp3Rfd+b67apGBwLeTkH
QLMGqCblog9jLYnDz38NwnCcVhDKLZZkxs2M5pGZPf6sdb+JdA5h9v6631zX
vx32Sej7fqf15IfGGzFw9IssGLPjBCfbiIUsFDm+21sMwVN8e0+U5NwvqvU0
t89Ql5mD7q8doy/jXd4+Eq8EtsmvIX4I36pNWwIH40VyUxyZE4FIQRRQJH9l
UReHTlgasZ1J+uECzgafV1RzQgk+iLM3dSHddCvaTGYvXxg/B8QmMYF6McHN
pu5hj+723opvICbYFzz16ZpAMFlh7aif27gFqf8dipH8S85p4Eq1E+lgyqSy
Fto3fylOsy9PJhmymW3GHirFNk0zqlWmcFLUEO+vnjpPx8ikbUH6I3u9/6g8
E5X3PsSW9w25FwfpsR45h58nqcZ+q61x3hnzRe7A/jT/4fVveENHlUDO+1HV
/RAOF+qen8hWA6TmDyEVtxWhz5ma1s0hM2vlJZh2HHkN+VGC9gVR9UJ2nX/F
qLcnnzWlVrxy+7YTr3/sNnTLqhVADGBtm7j3yzA6c3b2EB22VyZmMzJyYsFE
5YgQnMsenCtz/AQbltwsS/TbNcWiE0ExEpWIwjS6P8mzI68jm8Z7yhopCrGz
Ax/tJINntkG78YHkioN0uQV0cuAVKPhsvPQ04ZeHlbSh0S8S7DqgzwyiycIt
LH3o0p1dyD3X0U0R5LsGqcAzfHFuFVLs+ZP+wSQ8bhxcknqFyCd+jGUwGHnO
ZoZ24Yws3ekWPhpZbIjKtW7CJoR+iDJKF3Wt3aao/YNHJCEPA9fJd4GytnA6
w/HbuxJpjOPKipWSU5lkdXTNjDQkS2ku6Yck1fJEFV3w+hbQ3m3OuWwCeSQ/
9517j5vQuscK1oUD87TxZw7RppKZSqIywL2cJI8Hd57tDmoXZTTiW4uitzAf
RXWkQxM4s0uvkojE2OFJm+vcMo67I/Hd+ByJPiNW6NtL46yEnDDayUO0OZED
m8CZ35p+LoxNOLBgnkneLOMRjIOhtIT6tyGBLcbRQpYg89fVewmLFLg3DcqN
wH1ijnW+YO6Xs1aO5XNOTLVHxE3fjhr2aJsD2xWftbsCIhxKnsMlxNM3LKul
8eyHd5K/PaCCXjUezF+hCRr3MWGgkolISz0Vw1bjoTPhg51iK6OSuSV3a+L5
7BmwHk0uD8jG9WHcXN3lKPT4KqRlph0A3JHdYgUhJI3kMtaiSa8pFHNQmsJf
MEvIzxdhlYccrvTzfxRcjwq3OZU2SBg0F6eMtzVowgQ1yKGk1LVapGVv0j+m
oVGK17yQky3grxR7Jux5chiwzop+OIE8XLrEEcE7/L+ZMTeHlsHi1tvqAx51
tLD/mC2YDkR9aM8kwCXJUaH6kTbL8kuCGihz6flgO+W4/vmY4OV4WFAvRZnD
MZXIJbxI6AifS70G4duuP6ksQwvPPrvbUVtJQvbdHUwKLlwo7jP8YvZOzrrK
iMpiWDP5c7ZFe1Ub3Pq/6SNwHWmA2/a1Vgddd77rsLo6PH4/5t7q/wfS3lVU
1xjSq7mYQqXUizj+c0rbbzGUicPcS1vV32FE45V+P4WBVnwbV44fD2Wjw2Zb
lxX45tRQS9jgCJ0HU+uJ2w+kjplaKf8tUTHpsWoRhKPKzUcNsIJT9eqtFzGn
HjrBMf3G9V4kndbfgUDif5yzmGRhObtRVEPm3LLSqOvV9ME+alBOYztaUI35
UHmT8qOj3y6oJk9MAMk3oo0eiFuCBh0HKfFxpBI11RMo4z6O9coL7GRfC3h4
REenOuysVPZP7q9WiLMZoi7DEc+FAkuzne2Etj8JYRjmZ/AAqo7Z3zJTuEEd
ToYS7LB4uOqvCLBSf90bobsEI+HcFEOzxEUd3W7tTOq21vt+BQw2l2V93azb
ZI+qaW+5Tw1DLiL909/Z8Eh1q2bi6WMLtpqj4VeaYaPwRWiDI4YXfRkbJTpC
QDc3Un9IobIBLuxBRLj5Q6FU6w6QEnWn5aJZnElvA9bdNG2A74K0kUQ4OdjI
hWkuLWqITEWL78CYO/TbGBBF4y/BxZnjlTuVQ+WupZrQ7FsIF9lC/gBA7SYf
pzIWx75vrDsOYpKe9V2k+El4oWS6DEuUTJ+wKBdR3O8YVb3/BwrgsSB9vdZZ
z1xjxP5nOXqGfcea8qvl49nWo/v1+4dy8utJjl09p87GvRndWPiRNI6+orPl
MpsD1TUjh9haqpPKCLjPOGgNL2G51koTWP8Gk8cJlkwVuYq06F4OZ7eB5NzR
XcygpwMexm/tEglRAh3YoqFELfmgf1jRaYuVzfF8vXqjGAN4TXrXAaUjErvb
sNKKb7D0IwHiRcjY2FBXyROMhwPAc6O/KiXKtM7/tMa1vXhCVdcbQ3NrbwRO
cuD1dR/f2D8XZuGLqa4JTTfvSzBBaGMWVckv2uX/BOKgYUCyOTulVAfXfGL9
uHQfK4mLqdu0Bsuf1UPJZgdjTKg/4D+4KtbiwDv+A9qAdmzXZC/uw5BzFVK9
VcpPiiQzxZbCZWA/nKHkXPs1lDWLW43MSjP7PiY2e+Yo+b1AAw1jArhPiz6D
fqezLxmWG+P+MQhLlEhwK4yCOnF22gkGOubj2rhPMGQ7xN7h/NYFBzfWCnIp
6oIHWE8lRAKhT5Ytlc+vNHNhQJvDK199rYxdTCIwlFHIKLEEHL8Dpv8XXTtk
F2sole8GiqQpRNsgCJTaYBChdN5Z8KKQZjfKhBODyQ/1njWPnpaBlMBfvnro
lvKwb5OcYAOQKAVJKFvP+MERx9AEu0zZLeiDiRul9MWcdb477Oykjdyt3vh/
8ezb6yr82/Nn8JVENAVTdZ4B7O0hbpxzraJhYyf16yVRyThOi0nQ2wP+4n6r
6wc2AhQUOncM/TX1EGeHSLKCspWMUnbd4uGQ7Woo9JpXKXnCjw4c1iSa23c1
IYPJA18W8Ps9J5lC9347izXOIQma+EIqPMlSFwIOLFrIPGXKqc5ZD96lgaIy
Ope6/IRyYEDqcgQNYMSl+h/sRcQq1NjNX8PT07BlVUhF+nD1vAvsjr943Y0A
QAlTr5s7Xk6JW3xQ4RQYmfsEYiuBJrJ41AGWBhTWCoBngQeLF+U/Mz2fEIHR
G2n9hQUtJ+f4ZqAOL9HqKJRRXjemgWnEG+Cv20OAA9ZqtH3inlX1Mob/y1lO
SAFDJI/WcRfx1liH+/yMTDY2rePC44uwj65Dq9fnTlHkmVs5QEgcL3OkE0oZ
1tXMkLjbD+S9FP0W3a2ifLam/B2TS9QuSX+yjj4P6hWWGWyQZub+qW0lnhSl
pm/+8JynDYOEUFLeNsEoAftbJG1a7/FDJYyr21Syc+4JySOZCgoQ4pXSRxnX
6SAe3LwiaD3zE8p7ETev4AnLzbrV6kh1S0P/Pe/QuV2M1GiKbdI68tM1P0IZ
iglWwsPQB9w4XDUM/b4OgMwMt43y5cr/F50GflzuPVt4Cu2wg1PTlO845hjy
i7cHKgzFWtzos9mCFeLSuBRD3qJfb6ALz3LTYJA6oisy6W85ZNEo311B6xfc
Y54R7svYVjFun8armA8bUSWnfbnT3Lvl1r5UdlNhcTor2e5J8M/3BltNNC5Q
qcA/hfCNrnUAHyHGuJ0g8BTXiJzZ1kdGk2GO+JwmHEeArxnGWISvmoLwOMzm
x0MMO0sowhFpc+zyT1nrLOKo4TIwQsBQccpo3xHyNPYQTPXRodw9T0KJmRiT
Lc5Zen0TgpXV8nfvcxSVdGb44+CAIf2j3v/ZsoNfrrhGJRMdjYwPMGJ1EocP
naShGlhdW7gQriKN8rsK7JUPwirJV3KOFdfN0KzzK9YEX+4uX03H0Y94uLk4
x7DKkPJj4XljRg+YxtHVArWmw5kXBQ9KNrEHo/tjN78fNIkkNBnhXKk1saeR
6Wuxncagaffo7Ty90VWMMgun5zA3MAeDo9yrZOrQHZHPjG6zQB2eRN0ATB6m
Qlbvgq/wPATV07CC+GiCfp0LmWNtMw1L0qKETlZo8++imHYfKXGaPGjFY8R0
qFfQOEFEYRPPM+bpV1wTvkflIYykOyF7J8EYCgUcSwg8ensbppA61FhtYioh
91DYlAUfAWsvPai2Z8/HlP8wet2H5T590+irRVCRQxEEyxveNgIHx/ilS1Y+
ja7Yo8VTV9lEHr8y5epU8d/Kghfy8ZSQuDEGgDXP4JU7bRbslmfLSeWssk/L
jLo9AZ+79UQwaWdw8cuJ++9MUP+8yAetj1KoJyyNdoN7shImER/IFta66b5L
ieGzWy/TXP1bLpMo3tcbdNwAXYWIhBf1zhDJOXmjBImu0b4amqsx6PVgi4Yq
2DOjx4eMCVVdfuqsmgtsF8n15lRulfUBeGHDidqtFYG7pENzics9pTf+Sgua
h+GIsNcuQ6Zsi0/j5DHxNNPtAjRHI2tHwbdCsMlsznLEkOxW7tg2IYOz2weI
6UXu1zP3KOIvoqCx68uXZjV4G0iMhUk3t51VbNBXe2p+6sZN+7970a+C9M15
DUPw3CILT+JJrcthTN9aGkLCdIPCkCqmfAzwsURgBhO1HTFjA7UQmU6JqHuJ
2gIep3eA0YWqnSli6mn7usSEyEcr1bLmW1D+Nlb1GhNXd69H0Egr97aigZN9
0GyW1YMeTUxndX+ZC1uiz+Aq1hvGmfT7lTZNGs5e0sFZPFNvLczv8pfAFSNx
DSDc2kOILNaEcw7PM3ytX4QxkU5gErhrfnNRqUEMp2wHauei2r6hDIkVftLf
QRPFsRax+Gm3SymU1bSaNwu68T94TL0HtRs3/+vwyWuzb/MUdbqihEZUuhsh
VMyX9ehZ/5t5UEdy24+C1168UaQj6kFSPI5c9B76bNdrCFbT+VbjaTAsLJNr
PdFRILrPynke64rGAxVQj/cO6VgLWmXU96/e7YYb+y8C22uM+PavXWTP5EYA
hf777opUrptMdfIm5g+BKtoBn0l35kFBVvDXj8JtPkRJvM8VEezs3+Rvet2N
HEt1tGDi6RQk/S4GvKzlI4NqsXBd1YPXo0QOfkpBzuvX+ayjesS/drRWDw7M
rtsFPljjCoRMyz6P4NJ/sACot2FAO+qlxcXDdPMQ9blIR2fh5hk1KcVnrQWS
ujJSdgvjf0NIyOp95H5WSU8dSbuoQdJGiYhDELUj5KEMgGVf15WPOfj+zFxl
IE92E9a7t9C0ztFLcgMr7zYjP8nLeZG0dLAOkrk3bAYBTuuK5uYMI+bZNfTO
n1x/EQpOotXGDYMDRCSREFofhzu5fbhDMkRJw+DzMKq9FQAVACdNyLCLfz73
sjfsXOP4XVMSQKg1QNAY2HjSpb9zyjjm8IcygT3RWHolJX50m1L78CaA47+h
v7iq6JkCc7PhfJx0jFpKlKrd25ua1JGIrp8sLJNA0Df56PaHvzIiGoWjcPoU
Y/Q2cpcXssLFvnz/7mNma2GPobwf7aHdrYVgUrUOrN/54FGP0wvid78Dl5+4
OPdNWL174apNN2Dl+LR0BdXetaFykJjCZNkb94ursvHOMrtufiLJpEC9SoOl
tqYadZI5r0bo2zhb5iL2YQLzpiTvtkqdlMSqVtE7q7IBllhCd79nHfF1Si2V
dO9cxhBp+Ml0VqDHlo+WqpvMrDcezf7auvxgcAg219ivL7Ae5yvXtALaxwCn
is+R85Up7gl9hx10XFaD24xuOD35loSAyZRScrh12fga8HkKfOCwv1aStCV9
4aOHFbFFBz8iDlaApqOgQRJ9pJBW3+ODHNaGhkGl1MmbZT9zvJgByGvJ5aoP
k3f2p25Uz8lG62LVm0vQHXHMNu4xVfggKEWpyVuBRcp8ktKMtfV3KTxW60Ng
3QbSOsNSt0DkWlcB7WamiBgzUPRSCrSjY1Owj5fSdZI3+3Iyz2q/HZA7cQZR
4F3ZdQ7XgGWMXJ0oEPZbY+T3O+uIQCH/gkf6BFJ0glHUAYJjoO2nDAwvZlMr
1BL9ARAi6f2OBzJBf2c0rwwakrjRCm5D5aKCIVvxrDAmAK9qTR2ej5UK915w
XWlgLhw2hGYdbwGwN8DuDc5CFNIGVZGFHwQeVF6BG19/y4n0XZysvJnnuFQQ
jKA6peenY6m7gHb09PPFv2EDATGlCowpcFF3CS+V6dokee6hBInhRkOQQvYJ
PE3vmpbnq4JT4ATUqEuRG5gyJPK5gQRjl06feqgL6LNlhuKSyf1Vb6i5spkO
CnBW9toEICVXcz6eQHnWiWQ9SapAlqn4EjVJuYnxCOIgPoQHKGqEloWEU4eG
jgyxKl52sZaAo2TH5gcA8gMCzdBbPNkDlCOyKoJm4ZeClZOd5qZQ5sgNaLKk
EWjz3q0CCD39Na3EOVBE37uEiqLXfzOb4krMSUNEvTDeB/dswp1hKIuv+MlU
YYjiKl3D3sAKDHumHY0KRRyVjsa6EfIIXJc5jJdKjm7tKDTuIeMAAjIwM2Dk
6RLxmXkY+hD0eZcrXMXS0/zcd5NjO71cZVwWiw/wpDhPAjvSzj31ahfwDGzA
pH1s6ebPXjn4NL5YLMVhrpzt/eGwZipZV28K9Vq/tneQoOCGs7ZnR5/KVMff
gJHu/L4gAdUOd5NvNmzu5Z3P8pp3pjlN5bnktb2jp6kt5hjdrvEILA1Wpz8H
/50MiQvCqNxkKANBC+kneGbQZXB9bsOrYV7FewiWPw3hxl0Lbab7D928GaPn
m1gs/8jqx7ExXkfkBPTx9++BJFBD6UB9X8PzHtnbU3LRUZZ6nBMNNOcJzoQc
zah/VJ7cuBIRm/CL+0OBUxTGEOxr6h8DUMUVmnr7etXzjCzgSoK2NoxJeF/5
j61G3K0iIo045UkUzHaTi3ervH3xTLiwMcJfa1Wr+VWQlUi3jOMIu0Kyke3D
hcsfw3yert8v2uILt0EuPWyd8BILvj2cX72BNm6sNLOl9dRl9/eqcybqc5PJ
DRUsDAxoth1Ah4L5HVhn06+YuC+B4KtjZDQ8re81WL74tgtXJjAQSDFjVaBF
G1UwMiohsQSqc8Sy6DS1yOfFekOGvvwS+Xd/dl789KvI7K9Q6ExyWaJZqb1i
8/WCqQDOmLuioN45RZCaFHdy837iG+I5ddK/ROd2paHYHrvahyxEVTtr9y0N
czgrXPwae5mM2bgRI0PnC4ev/iZLmKGL0u3g8y3Hp9Himo1whbSuJ8tsi8+7
xWoKvx1l8VfuhjUmXTVEfw80tGijOV3NNdBAhgG3pi6vlxzzkLLaaMsiWRls
Fuj4VTR27Vd8hax9Fuhf00w4VQ2/t3hEegiBySH6Uz8OCJZY6giBDIhHygAC
/VXAp0nMNvlSVmCRUmLUAvitPHFfwWQLHYA+dgvC3dJEfZj2g2i/TQocyHSd
jCmyytLgyLeis10KVeGU3Q5rgW8sOe78pyjDXGDUKKNtrdw3VgC0NKbXFkx3
e0KgX0suLDZ71HaUdtDZBTDqFceylTFuMBHWRckihwpMT3ftxLz0o9zTD/lH
vk+qDf5a2+l4F7CvFjBuxZPTLv9jiPuADc9lq7G7igyO/qI9TEgMv8R+OTSI
cfshZS93+yUtjNaQu54vquz0CB33etgsEloIJ/qc86ci5ExuBEXRjqWOMl4m
PauXtO5bljDur4S0kscKMR9cJ6iPxc1ieqzdKojjxyjI+Cj7yW0/E9biZOAc
d8hPO/eghCsUGcXkD4uo547WHVU/Fw5wXiUdoP64S1UToaLsu8s0iGhjZCXX
cuS2XV5h+xO8T4qjTXdXurkm5ajYA2AY3bedjRiFUYXRBovVb0KVrhTZFq0i
lsHi26OL8BPAG4qgZZUMy7K1P9NcTmhAycbUL/GGR3ed4ktk2pHISNdl6se6
M7JW9AnDBkHonJqmoFcT+JDb7UvgiaHGBO+vDp7o395j2usWpO55W6cmyy2W
VPJHfFT7KtIi7ZrLqSLVLNEHIuu9rKm2JiIi6qgHFCOVxH1TSenzzg2Yk2to
ajrleUQorqhMY6B8iROLng0qu6vZMf7Nw0clk7ofaTc2e5B0aC3+JgPD492N
gqxY512QOX2dYaXfPgjjul5X/2ck2kNkIzHe61poK1zW7pBbMkus3zPyMNR8
evGNHreHX7w6isz1EiauOsOMM6CPlgSxkwD+kuQqDf0wn+Q2gno2UTg9qaZc
dQxHLft3Ozu1zVLbSLo4fJUtKzpnrR+ctWJv54E/mZ3zuhju/uqQ3PmvFfbd
UEsgomk9L5uBTdLAQtryx85bKtV9mRoryMr8/kjkKZCzuDx23RSE+IWtDFl4
lHuNDizvCGVvgBA9rZaiZmKjPRQZO+NpDhejn7czCs68QlM1Ymy2S8DZ8Cp0
i5UKqD+Yjh+MfeOrUNnB+aMfsi9eu0oq3hcSoSW/P1DIUnwIBC/qcd3Qq8zQ
YyGIySOacJgGVQsHWyjCxAfKS9dLWN7a8Ubn963B9cG2p2a/1N760+5B9tOT
lY0rdOQf2LcoRkqKLd48R8WpcklSSlgD+p3gaZJTlwR6ONAcj1DwyTdfJ4t7
MbdRNboqd9gl23wjE8N+kn6MFyC+LzaCKuAgkd/ODidX8bjhattajp8LsYj0
/E+74SntfjfKSfXzJaio+PHVCRnpoD7W2SZxYKIgAlAq7o5WuCvu7CSCgMwj
dW7StTflDHGFlV1IHySOv4h4HmNGAU+F62NNkNX3qYMS225BdIb9D/GyKL7u
OiBBmFTTc08/vJa93U6NsuAtU5HGZrrFba0LSmNsvrsfBYumWsxNL6qPNdvr
pOMBvRciwc6DqBOSCs+bCbVrO8+I8brQRJxLrZPvY3QfjMkZBpcgNnaUC09j
qgVYLVySMowc/YaLqln1NZ+r1tit4GLBJtW6hyRV9YGImm6evWBpVbd7CygX
0iVp357TRxLda52sCvZjDTYghrHr4DqGTM4ZqXiQpwFERc3ijwslqWiruVS1
OPctWH05rU1Ul/v4EJ/ISdtm4dTYzpuMh3cZkPJ91zas0S1XiX3qFxfeRv+u
7rDnAHCO2PL1tOpbc+4wlFa4K6FNAdn60aiJrBWQPWb64UqdIdWHJNBDqnyI
xkxGyDSPyu9331Cjct2k0+cxe8sniRA/I78MZR5vC4OKClgRdIKHrFgRKTtk
mVe/L+fbQU7ML8zixCqPMJCElMBQvfe4zX4uusblWZBEk/qdZjomi+OYz6ac
AI087BloV17pKyLUvfrPYfPj0CyDU7HHQOntePk/NJwxBRTVpR6hL5KBJMT2
kCHmsCcjjVhKRvo8CiERTVbH/b44jSlznmgBMjn2Lcdp4+cCOYUIIuFeTxGQ
lApq+d+JVjaBstkXNIU29jb2E3+EuEUNUfRsZP57FJohwER11phFSeE4yFAL
B3vgjXXUGDca1GBm4cARFN7LRSgUhL2meogBA04+p2hy13D/uo5gkeutpSZN
fPfRI+y2e5uWb9s+HEFXou0O6BkjxufNqchOx6kqQJD+FR/FFI3x6ZPEURrS
ZO+d5CAxmKPtXjQjmIMXSC/zK/Dls/u0vlFr4bMY+ZK1sH2YEtYwpMHe1/Ft
WCwQVPlTCKAV5V40W8QvQTlJCFz4VzDRbcWv2coR2Xu4dd/P7OvDblxHvWKJ
JXHWYmvSe1WhVm+vNvvMMUOb2U3ZljsUnTD3Q91ehg4S2LS96Zw6Ka8hVel0
iNCcpThkWW6RRIfzSjhOm+1X10YEFpJz/vTcL1wy31GM89AqLzt9iokupQVc
2N1n9m+z3P7pM1G2SV2QsYr5NSghFYUrfzHnxt+vH6fgw9dV4uDNI62k+gI0
OqAPQSic/eBh1rFnIozMBtbkauCG5rJF5aAzO//IKetaHg9U72rQ4LfSmapd
8TmdUsnjXzw/NRD5kGIqfANJClNztSFCwj1fgs7HWhVpzaYzpuGn6lkOA7hd
b1sQKIDpO2ZmOgiBe37LYjSAx0Jnfj8YpdwG9zVV5+ud1Biyqy0RCk7octmj
/7fZkaisTqAamVs71WSxQByey1jKsisSuOCnnCdo6P0ysSneSFWSmmdUtv54
NT0jw2cWXMtcS5wKtxc4/rHbmo/DiCK+fP1Z9a008Wc+CAPOkBuQiOD9M8L+
8B8iK6G/KCL7cCqdTU/sXlhEasiGVgLVD7I9tCrB0h9AgqDAcXBMF/3a5SJ+
hqAjsucJjT3/9Y6IpCxpSWn8j5kxxIwvbrekzG5yoTP7ruvgNcpzS6M8hN1d
SJ13G7Gqga5zeDQpBvOmVrrnpH6QleTaN1aS6bZ/OkaZDJfh/xmGn6C9lEDW
39at10SaD36UorJqbQsZ7u8WYznhBTiBilGWdzMSG7Juf+MAPNDY5vsV5Nti
1Jgc3SuNNd2w5L7HqWgxJQIU0j968p+nWylDfo3VF/XIuNXIqtQxr0TktvDP
FoaL7VlYHln7eu+qVRlxOx+qDhf3UC8drwVVnMoUhBC/nI5m2G8j65VXUcCm
dwkLiKIPOwitVd49oEu86dDl2xC7Yj8dwelFlNHqDSCo7vU61mCVaPu8dSBS
+ivea3Tj3APtGP6l2UP6mGVZg6EQ8WPasebYJ2AhftCPmRzE/AiCAvBBcV0t
wswgEOhm7FqdmdwSCuYTjgf/KImJfaLUEuMYJVLAZkNpbpWf56rV4qCEJAbo
ZKylYIoOBhgejF0NCTs7z/nse2lE

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG1MFcu9eKNrnaRCJDuKa3MrZC3NnA+CaRs7fY6XxoGexfpXi4hwv0/b1TwPXHx17SmysEvxMIuFYzn2cOUlU2oaUQSnw9ICH96v4a+OHk9qmmxH56M1ykajNcZioDaYuqAMquI0aCTgoFnOj+JTQBOyovZ716kk5obx9z7gco5QBHknDtwyIzNXtixcKm4py9Mr2Vo2yqnRpIrS3WxXc70bFb/So8lxe3yyc/rm0iHevgLbr+/v5nd3rCtJ00B516G6vPbA/cAbKq6HCo1A2xzyEWGe6Rsbc5md0Tg2rc17l/HpxInGkOXKnFTwAo0ettoaFfVoyZ9q0OC/MsuDw31GLxJxRKlEaGRBo9RgVWFiUSkHUVTJo0BgNeC8tznEIg0r9r5m6bUmvikEE6lQEtFT61I7b3jGQxo9K06gx3FaSRvur5mhUxvTvryF8iIkd3QLiy9cj+PkElIMHV+00mqKexJ3wqnI1ckhA7PeKcwuwOb4+KqQY7rsdj1+lQ4vgO7cZKsqYvVUamD+n2c30JZFHbfIzO41QZD1oUdgz3uh/u5TxdUHt1YHAoyzMBQqXx5MqExbr3bNNrLmA44iYdXqAUfDiAOIRxJFRf1EzFBV8sQ+1Yl7uz42/XkzI0LFKSiES+fUGUEdrKTOtyV2UTc7WBcHpRNxoQakZz0foQWv99do1phS6xWiFz7iJYuLMR3f8z7uWvXnGJn0pYEESVh3KP//LiAtpFn5wQIhhdQ44iwZLfrNW94u5ZdE5wJM/lwtriHpqIpDNxV5Yp0LgjRQ"
`endif