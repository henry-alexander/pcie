//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fWYs/G68ejpB2FnSiacU8zDOKOU5GV67tDaON0Izx7xx8cl8L8wqCNhA/At2
/b9aWBx1R1Ecoc5vmcyFa9vpoVtMigQyqNzGZa/c6X+2TBDHihFH1KXkaGhH
T7WxpcZVCbmiBOSe6FQlB9FW9z46uhbmPoTUlrchkn1a6acLf9A2YWBmHh0m
AAXMHFwq/yi3c17FzVpj2kd6EY7omjSj0MgwNKkgQBB0i6i/CGpInmlqP6Dp
7qPZ1223hYZWRbqaOzYjdx0t8WKGUt5wpXrxmpUg37ZaZSQMkhW4kMjm8CNA
15E3HwmZYyY3AhbFE5Uf02BzVnk4iPt1g8gLJlSEWA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kWeUT6hBtzq34sJbIcncV2tpY9CCeF8TWPdpqDmpD5W9msXfURmF3Fz/g2iN
dFe/t76/bkzZzLTrl02R0nvPTGL9BcYaETRhFC/XFVo/JoHpfOP+sFELZTiu
zvjit6fEss0Cs+7N0HafnpJAtwJ4RHeUE6JZ6i5Kau2gETzp+gyehiY3pzs8
DRiy+ePZnAg0DkVUqhTC1dBvUlpSdECZUDbWZO6BrK56zdRSVarrPhkFwBbv
A4z2WlwnfYlLYhqVQhX/XTYHiSFznJvhZGc/QskTkZJ+ByZNpJSqXkoNHuYn
XbuSIKv3LsW7Q5tE2mcN8ZFLbpGbTPFrTSdf+YAouQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Bvm2O3AhHPdlNwRyQpjZFRm6lDKY/AbgGPzWQ2L2cC3fb4T2Bur9k4Cy/qvb
ClmGpaWgBiyyEcJjjCMF94rqQ8fMcEITq3c2o6UbZikI8uome20GXgQhLVou
k6AyHpik0MGzhtBzYkz4S/ZESqhGalJ00WzzSiTFDko2jCJpNNEOsjDci4U8
RkeQhH9febFFOg4JGw/uMuR0/gdRrw7+H7/9dfkbDSQ0EB9MTPXIRqCOquy7
dpwYAkXDCY3bRoUTMRA4u0UQ/ZOnodyxgEJSEg5nFT39HJNUejeZ63zv7RNQ
TOLcJP9LJYhLRasqb2atf4zKCcw4Ez/1TEflxPMJaw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dtZQodizh5NlNtn7DeZ5e1mQiUgj1MlDVnT37hAhPidkDuuEZH5QymYoYOu9
0rTJy4Y4P7bg+y7SVaoYDgxMjgaXNROSQccqc5lVI6wZng8cA/aZbIJKgMeb
tTUalLLhYWkJBIvtVKTqC25AmQMgLvuNMBTFi+qHoDTmYOs0KrE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
O35FspRP+FmAxVhCc9FPnXQNlZKTMbjntdB8kdW8E0lZgRoJfXes6iurjJIe
X7O9/+Q8LW90HzrFFnwDSXjDviodddWa72l1G5hsFXR7AOOjluEaNg0zhjrh
Xunuqc0Y1rEAopYrqeAE124jMdCC/qeWRVmwAdZGFsXVfWxuth7bJsKKrFky
spgqBO9lsYCilCn6BrHdUX7Bq8swkYy1RvW4hvoZJmpLkEzNLktn6aPhnKEg
PC/fGwOYuQIlR2JioHE5G0iSch1NvTJ19aF/RdLRxJs1PvjlsN511m/FYgJG
eG9Nry2Ft3H7DEinYsgwhQ16tDLvkj6jjG2ARUdXYFVDm6XUeHL3ZoV/Xs7a
fxDcCi+1X2CjFBj85mRRO21QHd8/voY4pYfKh/TFKKwJrylY1tB3VxaZmDY9
KRqECaHRyQ0FJp7Oabn827PblRz4y9RZGdJ0wjEn7HJ+a26sjV7Vbh4Wu8Rb
coxufan1cwPl6YDCXAfFDJNvxROFK34l


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YPVsz31DC0tzOsEgMUVy5ntnhHaD/VdKHqnCpTrqEUTusND+86AoWIQ6I2GD
kA4avo8ztIKe/ATU3wN4X7szQlSavVbsHRUC4uhfAymEgMt/2qGEjxCvTJA6
LKSaWZ0/n4zIBkH4qphdmkUGBtxw4fe7r7x/DMK7/FSS58QG29M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bzrGi5Ss4uRQ24nwo9E0hK8W3ruVasRicXfUvHQwmrnoK6BQwcSmUdnpGH7M
gHl11WBRiWt/jngmcnRBT3qyTdFkpMvcIqBzevM0483pZLRe4bHMw+K2QmuM
r3owCtVqBHV7kBqJm9J2ffnoFpbsmOZm8D/kFGqs+p0+3vXUqFc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46864)
`pragma protect data_block
ocrZzOolQoY1svkbUW1mK3LGfUdK6mpXqUonokvMGbPaEb9AF3DWa7aFXraE
DVTJLOekMpkyl3QY3/wa5WN9D1x/aTUULlOLUL5NQA/WNO13PURZb+uTr84w
//OpPw2fS+le1IXDhFFlrOtgsvhzrR/Ch/1veTLwnNpsiuv69t16U9ZNzA+X
K8CQdx94wAkzVl6g+H3KuragcGFYvw+sUYJ79ZEKFP6OpKVIpe8Rbw+Ebghs
+FAxBNkxaUylsimC/eXUD9Q56a0ZHiN/zblEXnALEmukglaLtcxFLF2IVT9Z
aKgW2qbNC/udDQXFxuSVN8dw5Rrm9HSb1ODVhJh7+aklK5bPfbpvwmQud7qw
IaSonY8BUK9lfeSM1njqASb2jwjqupxhcg34kl07uraUYK6meSyHaFuQxKxv
1Z2WMnWDKR0FjbXSBVb/fbuka3iosEfLC6OAn+y78ysmiEx299Dc/4EyXRux
E00j/6OhaIowBenTY6gXznv8PpM4ZHDWp4OmLebZX2pt5Gmo21Wxws1q3tv1
7JjM3tgg2E63QTcK3+ob6SkLL5gug+1R/UnDbJ3eoQ35p494LdYbZ57iI7Hq
mu7wEi37EXRaXpt2fz4rLaN+VoWN2paXMLXh7WC7vRfFFDgdsYzUDSfqV/3L
ff4H4np9VvfFVEXm0YmcOt3K4cZAf4bYC0xG5rUrfn2J12yzE8u3LhtTryAn
pz28IJgZZYtlRMaVl0dYG1V90I3oxr1NRvQ10fDzhKvEui9PpvZTXFMaC4OD
qlFOgYxFVbYIdDVOjgMoOqdfmo6tJeJkZuoevAHE9BD8yfNSvPa8wO3Bjlik
LZG+DdVbAUgYnk7baPYeCr1WgQF7Cxj/O6Pa5g0q1oNYR72b4Kd9DKxh6tEd
obHs0AOlokWqU764Z2PidJs3cVfLmVK4bp/4aVx8DIdSjH7fu2Bd2ZDNHBpx
EyALsf88YTdl8X4qKZgyTa6J1isq7ZlywnDS01+PQI/5pWJBwBWMufoW6TqB
mu24HJbLTZihnpAKXvTHI+yZQ6DvT4tp99Xs48u29KrNDxmxdoWV686gRY8c
QSYX/jN3rILR40F7yyvNPAaMOjuxiTwrRc1c7FJOV4khZm9sDdA+yE9TdMP6
Bl3S1zBMBFXdNfydBNpytCzZ5vLazaaNHxabJfbppNPK9dx90LRgHu9Vs3za
hrxHX/yahxtOCRIBalLeeRGYyhn5Fl1CGvSfGw24qT5ZI/fh8ctIrvT5ev3K
lSOA4p6PQ0EQDKpgZEgvXQTTr4OBrWspTeBYi+Zxj5YlGGtHvtmvOHs61D1Y
8QVh1I0PlWkt6WKaLfsgBUCMayD2Wu2N4FSGENzhYrlAs3HyOUbL5eGqNESC
0ykmquFah7E7mMc+9ERAztDJz6UWUaEQcWO0e1gG9W5O4r71IuW21bdm/suc
h/vRQ1K3TpRieXRZauORsDlPjB0C2yv7Mj8K9qGlwq7cUQQhFtMOp8rjXKpU
fYYhHdwpuHsbC49lB2kJ34+9woy4NrqxfG2tRfolIFuvqmHKOzFYigmZ3pZT
4p2cMRml5/xUWCXTXPOkAHYrU+AD6tl8aDWjckHF1pAcWJlMxKq5Talq6tEf
xk4D/7qVw/JGWrU6ADw9TcXYCzsiD6xd3VHGPodaf8RvXr5CEjg9O0d/e91G
XJxJV8AXSVvOj3BUoYyA+M6a9dxGrnMOEqd4eIgaJDnpTM6My/7PsJxLFiSB
ttN4KMkL0ltbRE9pbL95iFg+J8LHU1MD2cK3aXaKFqAjjurGKGvcbJBwSBIw
/vTKcGHi6G0bhCTBCsXs3Y02RIUhw/UqxayEtMA0dOVnB0N9T0lZDVfOx2xo
ud7ZVe8krTnAGLHo/9O5m+mtqMJrZQTTIiSAlp97T3c9Xl0vLIxhZ6LbXClR
hbErLRAczQGckQbIs5OJC+aryVQEBAKM0mL7nomEsMMu5HPwRHJ5fNS8MIQG
5IaEwXCYFdDWn12ed9Mawt2oXJaRPt5elfohGFc/XdzQ6wA0r1FJi7AhnMs9
ioyrZ8EuWO4x0lZc20zDNjIs4aB3rK8Y7Xoe+xaWdil9ZtfNc00CPmz8F8z3
R0EjF7152eGl9U6unJ6R6XocWzEi3BFMZtlz9Maz5Jq85cG4He1jb3G5MOXu
DQpF7Otdzp7lGlZ583CvgRatWhGZ2c3tjiPB/K7U7Ptsu0VzxLXQ8KuB9kIv
LOdEJvPUe0qdbcz4nLPc/VRYnLHFoFSuKXUSDROSsKxfqZQJwG1BmcugdpL9
dtC/VezX4Gtxnj54I3qeHhVBrX+tD1osH3xcx3sbIsAdXwd/E4nedWzumLPX
LEP0MHWl2ToSwS+TnAgCTQlRVaZTtemxS3/gRZPfaC4GwIQhZacjoBzncuRk
LZVf97y6cKkwIDdC+An4nBuvRtLYJX3mSpxpyZnhXoIR1CUhI8bnc35v0+lq
1HRRvX31Q432BEU6q94eEPIXG2e5OECMYBigX0wczFzE5OSfRH4+/C951ODa
eQKvdyXl2s1BL6SMc4g8wiMYqgc2C9u2Jr0NSZ4ViJFxx6DdOeoeGq1ecPen
wFgF9KU+xVFN0vesehJCGa+PHobzf0EfK9Oq5D+7FDvrKtQebWjQi2lK+Hej
mrLajOP76dfzxuprCiDrX1G8SY5xweikuo29YcZFygSqc4Cl+klJrDOQBroq
ABMrldVkj29ui1WTA0w5nFRj8tmVAEPzcELlqxygqMwksvoo275TDjKC4+bZ
GKc5fRnEbxECXjxUI13dqmC0UXibqtXqbC/DpboU7sZ7Oc7E1em32hkhjfhp
t3ZJLTwJorM4ruuoknGOiEJWRrDWGR07ZZDNCGbDB1bo2yaiHXQZQ/guS5GH
VKBd5vLCxAPnGer6R8BV8HKeJqZ0MJUuREo4I3eu5Qiiizh/tSWPWw5tmvSB
q0gw/c1afgnusvPEpV6YiwCszNLSg2sQn5+CpglrkJ9GplQ6NfamQOrUYCIp
pBg7pmXHE7mkLHvgmWeOPPeoKOR+fBeQEiy3QIkpoWUrvaLPEkfyTu6NHH4k
C0LhKGJpIy2CJKKKgf5pfG2VhxBVaeKGFR3d1WKukFWZuqZr0Mv7kdItkgtO
MMs7LMwXdImJELLOpQG0h9GpIkhYyX4q90+bmlc7AOOPHm2i1jOaqnkYUfEY
KlEGxkLsUI0Ytrat2jFYcoaTmuT9RuD8MlYHeQ78cJIGvnMQpJ5Ug2bJlwUd
CUepajGWZrq2NVnAspPS+QGayxGh/YpjIKkjwrL943Fcb5nShDxORPwun9sO
8HMGuYMuRdcCPLal6YxVX4wZfWVu3U2w6PKVe2LbFNd85UDCeJ4NreTdnqti
vbs9FYHjsk/Fmv4WcuKw4OeNYX1tAMLtuumZ1FlX2G0Ls5GOX1MpXlWe66IX
lJ0m2jVFtrjJ9gM+rGf1xylyBQ2H63sZ+6qqMYj72SDBKkDGN+tWlYsiRiVP
RkoDnwxi2o5sXd3EtAJUqVb2qC3A6DICXi2h4Ce4Ik7Tt+0bA0AaZVkNnEE5
6Mv29MEHC1HJ0nKiNvHKo7F5Z8ZXSMRLZEBWeOEvR3m0HaWWRQS95uGRPwnR
w+/jVX619zOvqq5KliQl2BPuawGAUfS3W5nPXgXJR4wVVrMxEUKPoZ3GXC/W
4fYdrxrgF5i5HJzkSxX8S7MGj+6zXhdaXZQF0P2rihAoXVzYvs6dyKxXB4bd
omHK2iHp16YG5kBTbJlgDMOtPt2iCOSkqVyNkUyFFH0N6anRFv/9XtZVhs8L
EMm8UvahxhetH9V3+KU2QrpHUSdRO1Ltf2VhthEgIoei2hR7EeKIfEB61nxS
6ICal3X3y3DawwPdh3RSbyTBPuGWf8E7w+RtB+T6UzTAUuq/iDiUxCJPENCM
1PWCAy6b0zfqNxQWXgogYqJta6uszZezhToCX/8ATkf9976xsicY0S+IFVbP
Ph9T4Z15fwJHoiAlA6+8ur3VBIRpK2yuAtARDTr4U0/dZzk1uXNqs+IzEafS
RvQPfPWwj9626LS6aWellliy22GyIG/Ap71IHNg3l8rvgW9OE5i+8NchcLxJ
UuqWM34YiWJtNGbgXVH03z2gaZRVb8UNN+p47ViGq7NEMbA/xwVyZ93IlZ7o
vQ8Q/KSmSrGkPCjcWplKnVQjx11sGewKv+a5U+W6x02+DhE/o+su4cureV7s
uxgGc0yrYp6fpAB5lPdB6tReBNSufhQtYt/RLK3aOImqepJorS9nkVlADLTj
8v8VsVC9tko6SIiHAgpklrxOkSs0Eq1Ub//a1/e6myFprdkN2LyG0yRdZRsE
dHsis717efJHaN2K2LuktnKpS5ubCNuUZPCNiUFXqU2f0iWeylT4Z2gdd4QP
/H/x2nFg3B4upUv0xe4Eu4/XhfjZIni8K2xDDQPc7rmfem0TrXVOQClbLNfZ
uQc0QxzInwe+DqbChm0F1Un9RRvZUim7Ch0P2b6mHvMRXysiiceo/kVA2OVx
S5r2MtJ4nWSIXJXIptIILsW0Y6zDJOoOMbHoI0ueq8lidFsI0cft/iMZ+VC8
MgirDOwL/P1kAud3yuGsAMT2fGAklZiYL635hvz8lGsBwVXGoUXlZYOhvNRn
g0+y+sXk934C0/kTY6rT84hPDtjVVy47cEvl75MLSrZnqxSZ5JB8xuKBUd97
P6ZWT9qV9PNG9ZvMgKKXzbJc8oO+j2kCHni06Jhp/dSHcUE7vILWNdOuWEPF
wQ4v/y2eIcuET5gsepbbaMolNcKBNIsd+zB5nCHVXBloGg9XonXxVgZJBerS
+Lgj4Dq+OxzTdgEbjUqq78ouvcoYNjiz1+2Ch1vHBU0ude0Htkg2+GqBjpEa
PZvQ90kNCPqtjPKAmgbN9jXWmDZIYVeomrCXS4daeuUoljwzuE/aXRcHvYyz
/DvL/zd5p1ExoNMTaYmGzXQCnJTC4d2ySJjqjZBx4qVN6NoiMO9N7H3qlTUU
EmYUmaFua587apHGNSWud38jXddfOKMPOakFGa2fWlIOLhTi4KkXUTZFYBQJ
PWIoa6LYjVXT28Ii9neLSxUNSwlFZiOJgBetiCloDmjtwAcc1GlUN0by4yop
2aRAGE1rYHib32QTZfjZhMoulH6/Ey+b7B5OQUqs1+ago/vR6xlRKjmwFq0y
72miw9ga1CkR1y5hGtHnxMg+pE/3jxmvVJMTZ05ieh+BgfMt6ll1Ur9Y8UlY
IjefQdyLldHj4233pVir5rOIEG7TkClJ+sPtBRZWg+bqGs/1PVfcdDVNbypg
zHFH+Z69j6tFzk2LErkt487Q5IkTQnQC1Flg/kTNn2Qx15g7u8HouENu3ELO
dkYioQrlZ2uR7SkaBAh553oe9+kipB7ZekM8DHco2a4gkNkmbIWgDyTie8e2
fT0lVMb5f3LiTyFqbcq/muNJKqLmUQToE9U948ixNrW1RKQ4DxIoRTW8FiPc
vncnbwyooY9zPT1Q9NB9RX0WhebomZplQamIKegui8jya4QvTorjigjW50l5
ZPr8OevT4sEHXjjT7bUd/Sr62kWCaimJiRGAV1gPYBLNX2zlqh5dpPIG1mL1
C7z6Vh85M6iyQR58/dkfOKMc+odDcWz+gmfwtfdJ/3fooDM9768OmPL4Mv8F
HbqBUqRmX3bZ6Eb03iTIlgzOKkYV34geVf+ZAAOIVkdvEYiLEE7mNZ7Ua1Au
jkavFz1uKtSOUFG1cHUstebdDBoC0niACiTpt1n0tTABW8sl/G0qsBruWdLS
TLZPZpTfqokzR6k303LIqRY/8Qtxhst1G++gqHvA5G9jD6imf0OXUw3N/ntt
fMEl/AZASwXtFTY93CKcfYi51UeWkU+H5Gx55qFJGOq18J3i73NS/JDoD/Gk
KSw0qs5IkVU1+TGIzJR+bTKw0tVBzPJkFa9c5GGgV05phFL9MRX/SYhkuphp
1r8hLYX56N7x02sz2D6hAOsfKm+mSaqPzBx1zS6P09s78oC6o5vuVfUKi0s4
4wp4JpRpRmWcOX/OqZceEewaCsufQkK7gM9OQ4i6/r3r/mOJaH58E3XWKSVn
kPAcNy2LAnQ37s2zBahSU+DOWAXVWm40qt8bpiuZebUQLWcQQDo2PwxuD7yL
p5P+G4e8Y5Mr1wC3NV16rTHMdhNsq706XU+PDwoynOTdnqmTprBqxteDW11m
BlB15AF1u7OfAdtXy+pOrAJ1tet7ImqCQEjzAf8cPIou3Xkd0YQta+NL6pa/
Kr5GWNfX8qF9VKi4XSaQUC2989e3um4EmO5Cc/trNVicRfWGsHqPeSuJY+OE
fGrMaZ1H0WL3ds5dOeFVKUfrIWf/lg1Ciy6ISgMw+LBBGY0Yp9pmLSVC2Ra2
rg9pEgtreqnm/69IG1PQihKvYGERQHi+IKafVaEsjtJUoc7ty/Y2hDeVTlwh
Bh7JxkuYMAE1zY8Mz/M/16KOR2lMWhBZvVxb6jvRXGFCk1FCSbn5Ba4eI/zr
7JeGKvjbhMTYcYLBvrHTB+xStmMIZL+nOz6jM0SuqcKJsKQyFOhVEO19FVnB
WABQ/EtrTECByPcXgRaeth4HYCP6PRkjxhwZnNMmRdxUWbmQFI4tQN4l3GDs
WCD6xBvzt2GepwP5sZrPO4CoK26RkezNLer3WwvMB7g4K5kVbMhUAXBRpgyk
UE25ngN2QujyUSf/t1j6hf4VLPD9aZeePagBD5b90GhlZAylxUvwc9zbBCq0
lAQr9lvZ9SnYIFotzaMQugEwOFTmPvN1TSWI5jbS7zUdb14cayLexPZZY4L0
mMemNbv2Zvfapm+reHrXs/8MZjhF00Ozpz00phum/vJGvm2JsZnklJ2QBoUa
Pe2RYkpaacK+E/ag3MYYkJ0j+eLh7i2d9kR+uD1F5q7EN0HyVQ+Xv20julMb
uvJ/fzPR2T99RDJbhFYEFwbT8D6cWyJRp+HPXphNMVeSf6gb3QTPOlwFWmzu
TNx5nbGcz8rSEirINBbAufPusuC37WbPylLdKpJyCDbtqtr1dEjBmpAq/cQF
2nrmebhfGEUoiVdPStyJhxGfBIvbbbEGNr6ci2yG/4fUV46X599b3bkXneBC
D+fZD9WyKtCaRnen/lYai9u+5a/VqOI7nGTiNnIy7UDNA0j8r0rNjsCJfKJb
O8gz75lYd2mWqDx3VCRf+Qg55pzbFH/moBU6x+wjn4cg3tw5yNGac2gZ+YgM
o2uxpnLP7SVfHjmeWxZQvis1+LayhONtM7NGKbmWf5Lp1KndVanY1U/S+1t5
PYmYEDCwPlRDdOFddmNZAxfLR7QTUr6mE/VCMQ5wbBvYNtiUBtKqrj6BwcQ/
JyCiNQghMvQpanf8Z8g/t3PWymK5MzAqWhcH+VyiAGxhaJ8qgePBcX7frOhy
XJ10sJbmW+M6DJdZ7z7z/dm4UzTcazaWYMaNnraB5Il5cT0+cTtDVoh+32gJ
CwceVxGJFUPc/L38aGmiFXqRQIJ8Uyp8W2KpDFBOBQfIvKOLGMqSCJ5ViL0T
WlckAgiOS6hb4fw/ZZr4ZOvewwVBPVQj9eWsWTXPKSn7eaM4a6hrfOwz492x
WwcwKm/bS4LiDeO9YsHBVKmRNhoG/D+/uKv7dayAEAO3XVtnyn3nIvNLfayF
BYzvbBiCkyd76CmgvwVwQvHOvKu5R7O05r7Nsa7gO17IrhRS9mj+rKnQVfLp
bHBtesMATt4y8Mx1IMEsocm7Wo/7ezxCRhtJY1YbQn+KyYelpV8/+Z3Q3oeL
vtMSUMxILLGjbOCcncu48Mn2KUm8XEl/dE2eKaCDFscoTiXIX9durGTLpKyw
dhGI99iT26prCwSdFcvwgvapl0PJgtSFlJ91x7oUv7JQFqj+5G4NyC7Jscy2
hlFut5u4Ch86IGC1NKzgoN22PxSs9A/PhlVbNlpja4QYfFOdcOOIb5ZV6nn1
YCqsDe63fBzWgxm6LIyC/0Fy8gTzdaD8+KNVZ1VYbnNyiMSlD6577ynNBbDh
aAShVHQm/vWxDOefdkmNXtz4Oj0HxaOheVzUprTR3N5WNDbWHL2u+PsgiejO
ZkNeT6Ui+u9lOFOGoJCZDlMz6YFyO5fyOKdVGc4bbesPg95qV1ni2fTPlBzC
oK8g8R5zlRW341URgzQaGUmNOqzCG/fpRMDoMOr6cErQ/QF8Vffz7/8uuw4u
VHRxbsCeMs8zUx/YZgaY6AKB3Rm1lDsKVxpBRg+opCAzsD3AcqbUsRxr5CfX
Sh9uinhz8gSZul0bJlErw+RJ39jST/x3yII5HQIKpjHLfZVGI4SMrVc8HfRY
sV/i2CUz2cOB5EtqHlcEHn50cjyf8AxLQS8NAOBuHHcyP0jAOqJ+S7kV1iKz
U3Wdmb3bH2RF4lnQRH8/j8UtOL7YbSHcHv8SwzeEvkUkuRq6MRZS7M5GU64x
ckh6292TuFpwvuBYiIF+QLVKK1R3TIJHfleZNhBuA69P3E2Y0+qQGzW9tBB2
52FnzUUeSgWp+8THGDJpOotcMqjnxExMo7ivohD6GnbC7X4LforZ4vWVouoH
IP0iXEOApZ2CzBb77e2f9CSboiVktjS+wNucsfvHK5UCV8etm2pJfWcn/EPW
vhD/95VTy19g+PD4zropex4dfOWOOPN8QuznxCuOCAX7IWuritttJNxvM0Vg
lTlnONKZW/ZKs0nXIkx17qMI930cPVOpFdC1jCKewWK5+yR8f0m7cfv9CgOT
UME/Z55sFg+CWibCybDTw6sCF9SxebLPmZoUh8qUM5HjRmAZcSAlZO9N1WEJ
QujE8aaRHK76GGIuxXom7KM4zhWl2d30oTESVDr+erg++V+5DjTWX58HLhqL
w24rPc1LGBv8LneLMD0rhPdHOdMh2wnmdLSac0okdUW0aktKqdV6Bcu4AUwe
n31N0udlkIkWu8aeVl/zbkUjHLvwjBggluZttOB3jCRUPH19y1HrOXiK0xG/
UBZHaphJl9Nx+XGXRnZ7au8HOnjIr8xYA3Ca3xC+Tvq4NLklAL2iTYwIaNmh
tqCRdiqKJkCO2//TJKXr0MP8NcdBuNNNb88Ldld8UzIZz1AV4rTksfaWBqtW
CckrumMng6GP4edOaJNjN7szY+dPJWW05Q/QxsNBipFHNcw0DIrbxxxzJa/S
GWItUcFUmbsajGydAVxBAEfFbkZTLXA23FI09T8gJXvbsiTA0GsaT3mRFNKm
OQOUyzZkCa/Ar3VYgtdtnQFj8qskMq98DO/GpVagzQdlaqnlBrmSBC3tYoTe
suzCMqF4e1Yyv55mK4czerg/eXAi3GiefgeYL2joEMKfbqWKwrNFkLZAgB3S
Vw0cZ/TiqNff9p4ojsA4tEVRIqK8oK6X89Le9rDcOvjgjC+gd2iYshUPQP0Z
FZD51JHoEr1AF0uxiM6B8wjYKuvqvRy3ncTTUqIhFZkjzEby5zsIu6JKhpQ3
/Fnz5GgFh6mCcKbUi4GIf54cJ9QIl9g4LCLClHZXKvTJU6MClG2sZN3mJm2K
G/vBIH3QFMmUZEXdQ6SnW9awJ/v3jmjZIIKJCzJjPuB4M/lraHyvHL+22QuY
uLXi0idgd1LO0pF7IiTeNylUIbdehXiMS/ZqnkQVQYVyFwUvaoxj0GpRYprR
ag7ErIW20GostXdKxIdmYG4has7EY5S4APITq/h8JEf8WUnnsEJZe3nJzz8p
gil02FolkAk/7Y1RKnEDlcLk40X7/8pq67CeiCjjcC6wd0gvLa4T/MOBqpc/
W/lzoby7ufM9QOdWHQ+0urpSmDjIaxucB3u9gadGYr8u8N+9ig+xd3wqUeb5
FOF9903qYiHsYlms+fjD8RL3TjRk5yNT9MbGAFpfifhIEWbpHR6Cbgxk8j25
4QJ8XWGnT/LQFVcG+nPcEk7Qu2z7VtmLO3dgTWILbGFApHy9DIIyCEy3U0cG
N1fAbHwS0CXuqSHEXF+ARv4pFjyaWJ+UVW76FSMUI4RJYXe+wAuuQ3u7zQcr
rHwC5RsSL0v92hBHXgDMfSwkEVJmYiDbPHVeZcAELF1mbZASe+I9wcVMQHse
u8KVXPwdw7sJ8qrvJ3VEyIKMMGQLFbatKOIlfR84kvHBTrd1Lm8fv0FsX8Ic
x8BVs7bwnUbIUS1tnhd0T9Or2m7WoF62zrK8sZ12IH0NR8k2lJ3Z0NeGaZZa
aRq346vTJFWnm0lbDMdl4QeZrVsscnDQs95j+5vtIBlPeJEYaMb4ITk33xyI
mohoS/wZFjQPq/cS1VDqFKmfi2e7j+laQgdzrwN8tViO/zEvFUiOvakVLaRw
QfL/S05ZF/t0XqeNcYQ16iXJiOhNeMLjlm/MDG07vm+c8xzBFWSRgcSiGfzu
xh9MPqted20pF3obj74lH3AQ99BqsBP46LA8/DssWNX1/6IX94KbydJ9LaxI
7Zg43vDFcg8u+5HLp3WtXYeJBjykW7qW129aCg+ZNHRAaxFRdKxABAR61ych
9hxmzL2pogzV+RPhXP2kg9EaYVmDT6ttPphgSeqqLoiM7mU1eqr1X+65SwaR
SRyDW19HzB5fJOhbvxWe+1viK7NTK4mU6ypwqiNwP58tPEj8KNTFVtOvxp7m
PLqrLrLXz4s/ezQvuDpPoAOCKN1xFT25+xF7KJb0y5nYGoMPfmL+gLLuzS7K
aBV9dulJhIWOOKGEyP2cbRdFKNUStjD06btvyRjh4gBptyZtVDuOvF482slL
rMDP8yxT1uy24ukAR9R8OfVRlx2AgetdysVkIhKDy9FVQI/ERjUARlTykQkG
FaJoPwU6YvqtuM0zWCEc5yiHq1V9BuoOrXbXmKAO8xCOwfOwi20dPT3guMc/
mZ9ZxNF3x83HO1kkHswYVhLNIihthy12qYyiRmcgtUQ8w/PZhqoVVP4m2v7s
cGG7Fd0XIumA7DaR8b90vBIazhHyYc4Jd+uVJtJ5z9eDvddTtD+EpZHCPiX2
FGlJ7j8E8EChSJ6gREEq/Z8JNDThl0pi4skL9VzdRHdwu2vLsczIoSdLnUnI
fXs+0l0kAUzib9Ah/6R5HjKn0xAiVPuE00c2BUyHboXBpi3vU3DFDt5zXdtf
lVglz/OEnmZ5RJMTVoIW6H7Y6A2kJ0bReduHPwiQkkSb/PkLodNN96ACcCEu
CKnQS+rxTXGsIfD8kz7FivZ7+a1Op2pGMqr8+H6ZcC1dkPfD5E0zyApuFgiQ
ymciG5XhJPUBZ8bkB+73Evbmv97i1WNU+Tv3q6SZ/yY81z0BfOxmdYyNm1zr
OLsF3G7X5EcQIvbU8EWYKb7LHoLDKXQILJt0AdZZnO29agyBptY3luUj955b
kJwSu+GA/NiFp5rfs/Bh/vVVw9lETieExZ+rzK/da7i5cnQvu16k/QuBtjyW
al2nMGoyoRtVXPqFfGq9RhwX1bRJZPPD1CQ/VugzgbmWeoLzVTMt8r53HlNt
bZNypzjR/SRYnfBwk+W19UjHiOnR8G5+s5OuJC7p+2N7uc5k/CcrzQDvNSzH
9c865t8vvXkSXltm/hao9EhRNjTYlRzkIYp+d0AhVMHUbXhK02oWgKMT0R0d
dh/aUBwC1hP6rE3OG8ffoHdu4KytvzW1ajbTCDX0XX7BmSkzDP0Blfq45IBq
SRfxPD61V19g67AL8wswjnilB2zuZWY5ye1FyNK//Rbmzc7oIOgFhuVh2qTQ
iUt9Hx5qYKWcT0ioN0k9u8U1UvaBS2fmmj0ikRHe2kOgj6hhNnFItm5Ct8Sz
qJHffnYx34e834TEOjAVoSG/c2ChF9fSh6PjM5LMAEb7feEUP3z6UX3cvh/f
b3XlynvrmNz5cy2C8cSF/Yl7E24eE8M4UECQcXG9cqRmEjtJXTNwpSZGHfL5
AsHRgir6/Buo2l922TVEyZW8B/0JpgPXIEiLhFb5Df6Y21p6rTDYBTJ0drMA
/skmtPzWnCV6EJhYW70ClI0VryVu7d1Ruz+ry8MnuHWR/fgAvM8uNZbarv4a
6RuQoui44oqKynKFZmWi81HL/XAxJ3T5n5tel4AWxMO4wohHtNDdCDN+luPe
YiglZ+ARGFXa1SLGCyk1NtLiHtjHjbLkO8dohwbsWuG2zji1xtRCjSV9HoWn
wA6G/PkUfIiGVY/VZTDrEMpPM9Vp9ctnghgJcmPOokHfLr3/6SM3ro4HWHNs
DAgQZZOCQkK/glfk20Ml8aS0PTbj23hRkfSEGY6Lk4cVmGV8m/gW6Pi+IbpS
j+i8Syzml5ZOXL3uhec/J/TgShTe4g3SUKV7/b3n5XKgjH9tRM6I1e9BRgsX
++SsiY1yAP99a8VSd6Q+ZZVCVjneJyH76eSYAvGs3BwEGmDxa/fJCVsnd+/x
wNpiDQz5A1HFnRKSiqV+Co27BOWzJjekU2+jqJylr6dutdYkWq5FriOGIFBP
Yh65V46MzGw2PNZkHyKTmfUoJJhveP8WWwqwMslJENz31eVsmuuTTx/tGWTV
ubhP/ktxiMD3ss/tP2tOvdyRttq1Hc/cdP9omCe49IZ2AU3Zfl2M0vyxkq3w
F7Fxtoe/KcF7+g3WiP2Ycs5gIhdtOzaDMEo1z4i8j2ohcUJasleob4xLwsGL
UN7vwF0/erJ+8Nuia5rLwtcaI6lq5krIrS/EqnuM/ispSpY9rUh+itGmg7GY
hNivz1hoEJEkmGTs+bqFF84A90rvtPKKna+5Ze8SqSNVES7c0JUySzU9GSUM
bNs9jIbhckzS9MJ6E79vFCoo9LsohR35nAADQnBo3UDqBCoUH3lSIgfNzOa0
YZbJz7ez51vwQjGvCcJ9BH2DQTJ8GNNlhcGtxd6gA5AHPqt/7woH+cVabv6F
+I94HmENcbWQF7q9nqzesjQsrpxVyPSyJp+71S/EMSp4i6J5+EcXDx0DJguE
Ix9fSafdRGc2miCaceMtp26Ki7kK7tXYnzWpwUYd+uGPcVsSz+O0rw72jRyk
l3S5Euqw/6KahLC6nYeMhzLFwt7gEVX4reJGpYqmg5qExyO3OUyoUwJi5SrF
FlX4zvSJ5O+gg4D04SERs0U9lLnFs1b32h/Ql9wv6dpJjo+bGqI662AWD/By
CjtZ5Ntv+Rt9inUDCdCvZ8+R12jxvHphbk5cCF9r2Z4GjKUBBJit0q6JPAhX
SSURAUnClBOldlRMXPoZGNFuOwHHcYzWF59kGnzklOBe2Y1ygXmJfLhPEiFF
0AtnfLFekPCEp0bkU49bUriB4PlyGSCtOLWbvP+O/aBNH5ZCAdGkfeUi9MUr
RQCnu9cXOL8QtMQxUdVXTmNs5fJF3sf5JXtH5DA1Ww10XM06VqxioRyFYiPZ
H0cSh6bQ0p3bvY6WjsYqGjDKTej+PgjoY89yWXWwS0wasBculWbaikWWZhHJ
KC7DEeATk7zm6Gv2Z6PD6RDeLpb5p9J/XFJcQguywKTDQ+FPHrt8p6RbG9/s
KfEcljm43xmsjk+vZHW8rCfggtHoOdd9diNVMhMlY9sDihlu631XQadlFTf8
z8rMlDwRdyggYlaVrXaMeiAbLW3wTccczuYOdDoByx/wU9w28VW50E5YQ/yo
qpHxkkEILlJNKoomxBIYWzMPndoF6CEKfFe0LEdvqL6FccavVpBZDuWPWzhU
A1P2PdUtPiKR9QGa2YZcKYZ00SHOjdx8HR73Pr4AYCbPH5Ucnu/h8yKbpAc1
aSX1Zl78SguNL3pJQviu46Rj2WJ8vgMs/YDXfjPsaZrK3PcoziQFVSN26czS
mxZrQjRbQaVS6123SZ5XcWzhixQePb1xU9vg8+2zLMMtT0YkTqmUuZtOluRb
QROZ58mIk/A1Bn1NRskZZK133M4GoQRKfmZZn8jzFxg3IhJNZLCTsPtRhEJg
34UKlENsBSTYy3t7yiq7drhvELf6SXuEl2kWZ89OkYgwzVsPdsc330qRWip7
wdl//BBP0c3HK/XxI0qo5XgqhSvsOtuCZj5KvquQN8eGs0VY0nzyH2T/FugK
SkXDoRnUs5toYr1CE7DiO7crVcuRdFbILa/GmCZuGLf0qW9jx3bhZF1kdEJF
S5PYtTYCHSNYnwpgHjwxVRY4j7zoZrIGenadcEspk8NITAZCvizbwQNTfwix
crKw2mwRKXDol6v1KQDDK0IXXYBw+Lx4fR9OSdM7ni+X51CH2+oZOqmiOPBN
nKrIMmEu5LXQddRbIuHvIITbc+rfLl84e6/DmJ1Xdj5sy4gM/pY69M83OLst
wR7W/6ZZ7z+JeBA7076hlEU0voZjxZp7uZ+H1PDpAikfjBICLqiynmYMUJaY
sUKdDeZvenRVjbuV7jLBU+nQbVDxMgirGD52tmUiR1gzaRsqdIFc19VS1wI6
wS3LKp+//CSYGeBX0aqx0Bzxg/lsW8ojZEFaM/LkVmfhdMmAgLm7IWGW59nf
MHOnXF50ZjzsHhvmldIqPZ2dfY2mF5Xk8aVQCqIp2F6c3isyxtpXzQzy/c8G
nVn7af17AtS8Jh/mDNO138dI+wtGlUy5u6tuIj3iOel9cSOGcdLKpSys4aGf
8/cCF6CLHtQ//s5PjrfSwU07JoTJoYifopJHrGWZJuzCs1pF0sHiyiYLxohF
tAOv04wGC7w2dGg/Ki9vo9eLlafqb6k2OMVz4zz55qOgqVUQh2L25FHCAXur
/IedB8pzKbbmG/FAVZq4WcbZL+wc1H3xYV2YKad5ws4vnW7GQx2goJXVXm0s
SwGLJKpYxoQGXCy4rGy0qELVEofcYPgQ0nLh5KOHwIXW1xE4JsrsWxMVK5s7
zW23l2tzmDIK7f9SJaKkvgtcGh4TZAdVkveCTcEW495y4NSCOvv3i5upgIXS
AtIcJfZEYP3FBC84jXvYYTMV54hBp88iytmPAPpabdi5SNS/oeT53ecT3zNE
8MXF1aQQChwGaAFy9A+fhILltV69mdO3JjnBMTWttzsIvfQXsfp3Vs7K3Tk7
2MIMKuMFFQ0VjjNxXHpa9tMUi2W2AtuL4IXef5O2BiOQ6n0nK7PdEWufxiBo
WrNIry3mvmudn9cIkJBYN3hKqHTPD9khf9oSFLdE5mvJEWHH7yqKtkz0bI2d
NgBEDwFvNGgsXoGMAphOnF/Ji728KuvN1KtsWo0klTiQgUREivs23DIsClpu
XlvoLASGLyIlyjRC/Toe7jw0D6+qH2Izm1vobAZGID8DwUHDMbM/XqVJMTWz
dBHjElZnPUwZIqSIrsTPBiXAVyAn7QzXdOLWkSlEe5B2Bax40hEZDxEPXXtJ
RoxHYttLVoSDkKI77uifDdBB+N4jw1lgzjGezW9meWGVNszx8CVsdwjg7c9c
WtjGpzFx6ROWp3+K9v1uwTKFbFH7dtuRboLh0WfOaXV2km1ktGUP5FwjQAj6
6EZNlOhMIByOn79QsB2v9SYjn+IN5r2LvxMdzjiMo/x/jiNH+9xTkb50vNX2
ygN6QdfouSB4rR1m+ljvIG+joQJ/4IIHVAPJiCtIdh2svqd1LNr9iHCUGk5v
LIpLOsy7PM7T4qXAVP6LYxQYySXTy12rBnkfBQ+xgt5/78nlLPMFRfU1Hlde
NSY6M/3mmctMWrFvm4/TTF39RTCQFYw4heBBaGl5Uc6zs5EXXrPteUOeFxg9
/XMR8Teq0wVrbtzREd2vb8T3USiNkpOqzwIF0+7TgjrYZxkTxWAKx/CZhH1e
Es0izfuayiDiPx+WBkWipu6zyBTZFsYCbeLsNSAZZadL3WLpmkK3cO4YZz5j
z5xNijU+dSBNuW3xdm8I/DREPDxz1Kz7Jzvne+XImv0D9TVJWTxPozVSh128
MAElEL9mcV6KM2RbQ/XL3VWYWBlAsknzo74Fxd5DmL1rB4AmXcv8fmdUW3vb
1DyPa3ewAftKm6rXKZv7+6TYldj2AwAuhndPP/PfstcZTZIu3PqyIe0Mt4Zm
La16X6Jmj8YRdYq7MjiTdrn6bTOv60DVMdsiB7IZqlo5/xkZCJ9+cinngCgq
zYI1Ef4xAVSq3iIz4BCFXnGOGxkOOcpMw03cWEcDUY0i1YFjYpFt/WBhJAZY
J8x3rw3ftkTI/U42lUAZm5o1mxtKvhFptXuFJBZfHkFYELsaG7Clh4h7QKaq
MSmDYK8CMXJ6TZAvTXJfI04XMBzDxEwwsVii1HIN3J2xp+ltAOW0d2CXAAlk
NuTrNwfrDjLgFx80opYXyscakmbV1Rt6wyhzFyAYtXDK6ZnzxoJzlaQBC5EE
bub8GBTJLFslgtcqvej66ZLzbrdnL5wtOrUVOrOc9LcngsrDAuWf5GN35nXp
PjPgIkTlFQfUCqvwguhoYtIrB59yqqiEnkvJ/x4zr0VNPFCWEC3p41Xj7Kfs
sQQ4s6vTuejOr3b/FajqkC7iNS8WeUqEayceilW8jOjoL4fH8fKUIKxkS0ZN
5L27XrMAU9MxNhPGg5JmQmWk8tJH2uSfxzgElq4SKOimifOO+Y2M1wuWmWYm
S1J1keztZR64DvCjgu1/sasBLHQNJCa88eaB1eNvjQpCb38nhgS0KAva9QNn
CVrEDD5ly5advUJbEOwGGEs7UhhO6WiqsZK5yJagfh3Os6hbcw2qa0xQot5D
l+31i2qT4kTa2pvFBf4Sz/DorngvA75mswU0xIOD8cfVacysQvFdQ2A28C4Q
C5OGBPJqrE7vOYwpulgO1bVidbBrRPExkV0iC+EE4PfDAWEzXHTaO54YbNkt
fY9syLuJgdIxElvtghDt/S6JQq2NIWjaIb5OdEpTp10YZ3/CINszbNYhSuxy
KSJmgzIQWVHQuCyhMbJodK3MGVUtaGseOxrh6HUtgNgj+bMl7+Q7fdh1eoUu
MdqQtCse+uYxix+GvDwf4BFDhAvjGKI/W9d5Ws+qRqmlz6jjwj9n005hxGxq
MBo7oWFzT0JJOsFJA+9o/z3tOhXMkSaOtjycaHpND4t/zJ1b+CWuZBS6/NFY
gWAOTFWWt7GJRhduFisR7nabjJUKADiIpVLH1o9B2EGzGzd0a1VyCxKfGqvN
//ExiYUOthCfHyWM9dCVQvxaAscE1m31wYESjdOHvm/kLYt52aUnL/aIRMg4
5t9lbK9NmhmZfM9HkEaWlhop2L7UHSoSxNcPF4f+EppZXiEFp3NPNxWzjLsf
kjGA93OvjMzJBG4t1rydgShcW6FL28+8qu9ZznTu8mkmr8rbdwi9+z7E3ZWV
RMBZOSBpk2ZqEEYKj+giCpN5oduL+l/ES17iswpnMKrgyRXcYSMyP7Zo9hg0
H+0oGAXDF3tMGzlrO2WXvLbDqqh5ajxd0tD+2g+asMsJqv89wESo08lzrLVQ
EipOce3CAZsNFzzA4zjqMoBiMrMwlLV7xwjpUSr4Sps8Q35Y15LFTWZdkYYZ
9Bd1VMwfA56FzQiLBgm7c+FZBv8oO5zvL6g3Af5wFoRUSxKXvSPhTSYAjoGm
FiwWX/q+hAIxpr4EKGZYekO34AFe1GuwocpYukMzkioy1/g0UGYUUus0lJKl
tUKG4g80KMIfxfK5NkUXti4cicjRNVenW0adneJglBdBI8P+Uh5l4cPP6pLv
ePUe5C9Omq8bt2Hnwtyc53D214Fbs/iM+lVSahA3hR1+9nmOrzBC1iuVGcD+
1MSLkOeSjp4i82WNOzy8ecggWGpNKvk7LCBs6LOIv5zmRcON1HP4r+fRbTbX
BOuSF0ntQy/R2L4jmDz+mVgIDQMxRTM4qxEl8I5/Opphlefem8ATszQb5GiQ
NZNbSkuBlWkfe5k6slFDHCnvijprBJj4U74nkLp0w6GJrxVRqeZciuJoeC5P
DJPvTHHYjaHZF16DAK0RtJZcFmwtTftN314kEtTgM440w9xjr/14m1BwhJGG
Zae7UafDFHXxsXZ627dks/xDx9EfT9OSAuU0oYyoZGguEBOl20fWnu24Du+A
9Rgd2HyxoTpaUw4787T78bpMhHqKXXs/meU7eUbyUd+H/FKYYDtDGaSMj6/7
J/ZGwEnvwRVrRpHf5NHGVTBcL+kQbAi4dWNk+YLt+e1uJP6+eeskOoNfMvtj
gFrCS/LWhUk+ILpHY76/4FTb4Wmmgz9upSnDz1sMbT+G21yLCkP/xMczDm9f
fz1JwYBPRaRj6qLkOG3Kw+p8CZUB4yUxHcrDWEvFnbiTbD6lBNApPwhan4vp
18YzurIKZGG+vKDZcOnxg/DP4vZ50HMhqqAbxI2s4FM4bEW9Y7Zy1P8en0T3
rmdF+0gwh7j5vDnD+Tmno+qvLQb46Syskz+WwnBFhEqNm/TRhpAQmG2jw+lU
nsUzqxa5DZAJt7BJwUqpLrepSxL8hfgAxyJge1nPUH6GptnIn2Tpd0LPYDGs
7dOw5K5byJu9cyz5f/krq2HpH0kamVZ7gI/6nPBFSrkKYSG3LXuPYqoHi5p5
dzxqigDegskwQ58Y5BgsGyPVkwOhgToowQ4iy7HPv7Gpq+49mHsWhSPKGjrU
XCfXREzohIuBHVxvoLdOxXrkg0JnV6KqaJ9+PeGIRv0V6LfbiGcRt7RtMbyW
BE1LjmmY0dy8uWtLgK3wEQM4Xv/jJfJXjbmF5naPLRiBSt7Dh0pEMovm94Au
nC34vlfEq4UyedDcVespBrPZU5f1FMNPIsRFE/J9bUdQ7M1qtObetCNm2Hc9
jCpdhU/dN758kJg/xt2SSzXAvO8qRacBNagdn0W5se+4C1s9R8ajtSuUj3fG
HefbnvW6hbbYa2Jb9tVlTUnwnGFOUR/pzyCbHyjK5UdUdzoWGiyeMzWmn+3w
ioBzsWrI55O8OIIb85eqHKri3sxfQU+T4BQqAssFZOqsA0WV9Nq3aH1lPt3g
U/QgwSXLoG8x+leLSIhmdoI9S10DPrYdnXVmxaQRvp3p6hgmK2oWXNEd8mEK
fz41ZrQ8Ir5h59t48alu6cBoazc4sF8sM7716AvDqLuR2NbS/NULfH3OzZmE
Maao/JbVrQuaBDL+JNuk4Zk7K1ERZvLLUw8fA+msMUzaaUW1XAZQ3Z82QwDe
Da9PQ21EFw9xRFwjQUa7dyuVuUS/zj/J5h2BGkPQk2oY0My4aKPZVR21eXgc
r22oE5U97d+/SZ0p4BLFYMHO0T4et53DY0tUjpkUQCdTf/pMA0LS/sOaEeLZ
jdHubOrnAxKrDbwGTu4EE5SuM8NGEGTW/KfJzG/CHPVh5YQBmyyOXWFcnu8m
YIozIsqwD97q1xVqNl50wtY71nJJgYXBdBxbNZardWuUHAl7awxriucaWur5
B9uN0/6tIX7WF+JY4+ytdZQ6QVMJATauYUC45Wte4a8gtZlZdTtaQlFm4PEy
sElS/Jv7lShZMQ15uJTd9WSBoqzfeuR0uL0i4aHw348IKR+QlT6bGkfmQB0H
AjAd46eoVN3uKD8vDcbCe2/1rSIXDg2+uslRnvzLYnjmKfBOJ9pD1PDsyvQo
kKZxpIZIFd9ST40ik6bBO37OGzsqOW3YYE5mmDdIiptm+67Io6YpB+ifNqdO
u/KetNysHv4zMaxzB+czAWS/L8VQcl6vh5u1KAJM8DoitJIPfdcO30K2YOOW
e5FMCopERFX93lS1MQKEuoTVEqMByb9xpK/LX1E9f42ERNvhT05ZMDMLGqcf
qWMEgTyeyOTXHGPWMw0gfd/IuVJDCztstDJkkcJ2JqAth3u4wd1oQw8lLcP5
r0XBy7w7kzE4/K4aHnDr3v+5Ko2oMt0kprvWqThaPy8YZg/oXscA0BH5xIxa
/xFYFhM0lOtcV9IbKRDOjji4ukvTA/g375H5S2yc5Bz3hhUkqOP4civJSbX/
rEubnc2aOWVvpjq8w1EKSPExFGaurkbvfIcHuLhtwNt7/FN+Xwohain+LTtx
iNMK8tZKs6D3QcpmO/z0TLuVrnGt8TbIEKg4J1OdVDreveeZWjHVpoMG3py5
tmMVL6qwO6ir890x67KYsyLv/xawrTF+dBVtwoM0LUD4UtYP/+hoOddmaxWG
sko3nrPCjPdHxDZeaaye18b241m6059kmSyGryUTSsmpWScii8VSPa3yHBUW
zcPkgRTIW8yIWLhfJfOODISS546/qnX8Xba+atwZQh3WkfPFPjxxyPDsKWO+
GwQyCZ46E1t2KbBPL+SpwqHSZPoa+r/Xr5pApZJz0Mz6UtZB06VcbjSablki
+6p70RrtcQYkQ9BDVOAyFph68m4U1fUdbL7gl6gSc4QeMmPiZ/ASQPz5szl3
948VkEV27is5pAVlxSs3ZjvtWgt/gFjnX1bTg/9jmi7xXiksjdXzXlnaYIqN
0LGrZ7Rj9yeY1ilW3eUG2vQmPNn0/PWp2VGqvLHw8C/bAk13DmRitZsRh/bm
Be6PUO4WOc+/dU2G7l0+o+G5CijAb5Tx4NERHC0i2DY304Kleu8iMD++gW0I
gDEVdMEZYA7d5MSjKtQStW8fcsnkb76MUAqSez27s5FMJLKpACbRhOLhOCHf
qQxkiFcwTuY+lm2XUkfRZvd4wAI5rmJFCWK4noCz69GHe9KXmEvWHg655465
9ULDXWuLwi//FmtMxSmiRMpkKOefTMUcSLNR2cD78rb5uj6U1lwB6qGVtHXL
pI57GHVwrWdO0O3U+ViTr1w+vO50qAAMj8U07hEhmIsZ3kHG3++CYDb+J/IQ
LxVLypEYbORlYo/QlJAHRyjs9kYPghWOVaGOV38cNKzTHKK6hVlQ6iOz1wcY
yZfuD5WwMDWbgW643B5oPf3i4jW9Tb+eFmIfO22zFgbkhXqCIXtypMJ5SOPp
bcovuqqMnamTgZORIT03nd1nKq3WznmZEIn1LDVl3KJCCXxigVkATJPy0/vs
KisXHrNo3JKA/VFwkI2fmk6k4HWJ9jpME0X2h8H72I9K0hVsvNgo1t0gYQoH
1TFlNK06d/6BKXAh/n/lOSFebJQUZ+8ITNsF+pXMfpqnVLVL3xN0ZdtyJdJH
ZwgMWmrVgVXnAb1LttwYFBOWW4lwUmu+QgvAi/s+MAeulE6JZUnmr94kY5Wx
KztGbm9iZdYVS/ws6de54liHIJM9r5gxwDWqrNhoMSIIitxVnMMkwTOPzZQu
TIk8OEn2ZFPl/FZFRMxP3wgBn7iCTvmdm0Vrseo7aExxab9RBxZb64Vj4M5c
eRkEAStK2DrHWy3bOIf7COxQSVdo0EXC4E6+vHtKGPEcn/VOpFLGw36F/Nuv
OpaBqdyfMi72yilmB9D/PUe+kMLjgtMvQozoN7i7pXTAwf1HqjD5aFP0s2Mn
FRWoZRpSWTdjMBkCVBU4hu7yzooEehrCO65Nx9hYD2fIgAwcKUu+w3uVml9i
DgGHacPji68JwfL0/p01QAv+fTSYtncwgFSMYOYnkXNdIAwACL33zDdFKbuA
Jvbos6FQm16ZdFxYSr4J9ovqN9EHHHAHWcm2aYVaG5P9qxJQ7xoQrCgxb8PZ
5Go/w0SKR72LI+xbzbMyXwaV/X4AvsUm6tnuRviw7HQnXjoICLqsMgKs4gm1
Wxva3KR+3/vB5nbSK/5LhJWSRP3g4CGZ0uWZz4HzM9zvWcccXBt6iITSKS+i
xZtei/NWix0vPigHNjkyIdj41e+syVLeyN5tb672I+em+d2AWhdBqvGfOi1M
UpvYpAj5MvM5O4iNqt+UL6uHiLA6ZvU+lq1RsZVDo9ikn7E0roxXApwPE/XE
kUIWZLbJNqSOkaQEujdFl3F9GkgmudkMsB8wSOPtwWKkglKcKsHSo8+WH5Pf
ytM4sGr3T2f3Iye62tdvpbk2wy/AohErz62CndAXllQDTr5/1QfLCp2KsCq8
SX3uMk3k9T1kgQCeAh8zwztDBxzOv1xvq9px5nckgII28/QpkJPRETs4DL7K
HmQ+6GR/zS89XVnfKFBpcRzcZuVsi/H2I7SitOp3FN1IvcqnoMzpmMzB+W45
TDaK0xwEXB7zBqyPD2WbUmIeT7JLZykmzuIsdu0jR9ytq1XwyzPxNeIj5JKP
66ir4xLoNOW50+5GXWkMOxMFLmxsEfLqUCFOLQGEd5PEyy0ujojQWUdv44EZ
l1GIHhoyyVTdDBrbwtHRiFsc1E+X519+BKMniUKK6iG7+eG+OpmCudtI1VLW
aGunNT9bxU999ukqv1ZD4uHredO7+3I9cd6YcyKYdiACK5vpUybeh7WJ9tAB
rq3nH6tCasqvKHMagh4RvL+EuJ8kLwOfzUssXRNGEeynCPHybPBkKBWrKkmZ
0XYaen2IEDlIoE+f19vP8R/rKZ57AS5XP18a2lT+tuHQvsoSkXxMmsVh+iaX
qXtXQ2fcyKif6uXlDTsx325Qer3K/KCeD1F2lzFd/GoSOOvcVd+KG4v2tCa+
AAjhvlEEECH/LmH0bZ/ND2Wo8UjjG+KUc4gFc/MbVsihwRoC9M9qxqdd03D0
v+LrvwnLgDg+UZ+GP6McUKaPCOVgUAw8vKPPhKReteD7KH6arGre1Wevl00q
kmVl29wJpMpT2OFhLczyTgkMlmRwkja63HJuUAqxz8JbMbw1jxRURxN+62Ye
ou4foJicIVJrZVcAkRKt6l+eoiHEQC5C7kgtEGAfZbyHWgJmfLRUaJL9YJZ3
lWJxzl2tnB0Brs6vT8uyu9OdK7L0VzWvPc9qcUywGujBgN/kRKNv8o21GcYt
Lg/WO3HK4XlAp6InlYV+cpqRVGiCRw5V20O3T2j7iON6t7z/v5GrfuBkKbSd
HkMvX1c/1KhG9kL1tBQ6MioigNVpyMZXALjVu3G/a+7MsnoyKYoMDdKj2APU
8OJko35VjHUDKAa4oTJskhorKaTy2S3uO/WzqkE6XAQdHPxB6M0GQ4Krr/LS
Nq+QTEzT2LZe4k8A3aHrXz+5TkQ70okS/twJ/65do/eetx2RHIyU4/Zr4eK2
3vLmrCVfvhosEhBOjWhSnBhXgjA4bGjYR+oEjIL+ctJ9BcURzAMkH8OBv6qH
QmGcaa1gqequ5nuT0yyG4wZ07YefOWENYAUu1njgy+CaBq9tLqg1nlZU5q08
4Ft0S1RlMhdfnHd6CbqKMkYNknR7qWuuJDKcqBK/QlQVU2IbsbTTRY0Bcen+
czawE8x+wLPAX1dAN7EPWMOkSOmeSCwwbeLJ3p4ASjhmLd4atz/O0tQXsrhB
uxroT7JGVJ/H8b3P1IrvNRLweN+CD8jMoOHNRfTS0ST0iGuOr9YYXCBmGoh7
eeWQz7ie76qFuxWs3MMkbBXrt8CogfrcTK9lIkpWvjIYqNx3FUZ/N0zBzU6R
poV75BKvIWDsRNS0aGdEBsNNVrMu7K37Vu2NZnV+6BSRizt/YWIUH7NdZHZa
zw+lKJn/6T7ijz/1CBjwzrFiChr4NRaH8g9Bga9zFiuWE7arXzEn1jQ69YF3
+UC/NfqXfu2PPa+qib9U6RO7MiGf0BiJyhU1+Ypko5x+1nWZQOFopyNjx3U0
IVkuyUlKJ22hdHCJ7Kyqp05WH19PE7YuvmjTmBfHH2j1mhVdAijgFPYNVLi/
WCTC5E+qAL2w0KVP7sxrExUlBhHcXY4FmW5sEOws/+0ZubEguwiioJ6EH5Pk
HBm4d9LZU142N78x37HXVSucULczQ2gu5aYvMlaK6/03xKOOJeDiXKepL0rd
NjirppGgMy5n2xSLiASF7QS4FGDJXB16vqBMn4GX7xGDgMD2yuKer2cWla9U
d56Hsz+LipphZxJQAaFpueDDDNhzuotN/esT1/9eio2n4pWaYO+ZcJ55JRyt
PgjiCyuF2431rTGi0Hv+OT7b0NfWnck91eW2l89xVTMZOfB0koqWtd70W6Uk
ZCH3olnzggccHcG6/bEwQKu+Z2hzqfsmpsLg/a7WwW/MsBVQtuCXtHnM6M5M
xkNVGfG5ZgwWigB8kwlY5Q6bjk+no8aXaw6vrRgUgasySqySYeKd4TFaZKmg
G8EapQ0K4JopVRz/qpY6HneSitXUpOHddRfeS/9tx0GdpZg7gYJAHAsYTJND
tCOL2ehO07pJWmS3aSltdVPmWy7Ti+BhahRL1WKYuqSiand3/1qih5/GHKBI
NB58DHBpPtFo4oR7lCpbFqafCLuCefjef0OBuP2rosrYN0UAihLj2XIBZ9CB
AmUNpYtu8QzW1VLRkucYBk6yEEq/PGFCyrozv5pJKasmflPnSv1IWkaY6j8n
m8xkgNUWuV6bQ524udERYime6CfP6PRMBJ0Y5XS9plhsr2kLtg9/PBbtQhes
ZwY/uOr8KfO4SyTktrqN0zf3poVLlOPhYg6aaQdSf/cFnQdGdT5pmZRN6iNY
mS9zlOHLgqkPJ03rZthkNMsfa5gm8LC7/imtWOSkSOtO5eMNJe+0gagUjPzm
pP3ukEB2DO/4vu4XGmaCw7EOVh2yk2nvcvrpcSXvX/CigAkJ4PaTlh9qqS9Q
VkQGo7cwjBrEI9TfPh5otkTCFDDdn6rpaGh2yhbJslg5YY9HZgWCiE8tJi0j
OugKWhthsBE99BGA3KZIyhF+MjKRJ9NNwO/UcNkhrKRF8BSp1Tszy99ZXDSk
xuQyngdOEwUOQnHV5OMgnsH6QhPNqmQQRR5episK90vz9W9jAybni7414FnZ
u0z7giSeBNvhzaShsoXJFPZhZrIKsxik9nikd9MAyCmBlB8iXPHM/HfG3Ayc
vqo6uP828H8iRfVIYZ/FC/3MI7xMpRF5TkgCKIB/XFED752S4yE/dJ6VjQ+V
3EpXT/bf4t146nOBij1QSYdOJ6woDtn2Hcd+njTmjJp45lUZ5qEjpYWd1SEo
oy6rtgaswczFqv1p8yaHcgJ089U1cxIGdRtnQ5jPPZgY8VgQS3Cl3pwwG6dt
8yFMrdB59gK5EIBazifpZSoNgSp/6G7AytLMU6ScJ8rppj8lLrAL0Kl07e7r
h9p+syAjKIPlYaf+S5H3c1320mSTMBovFNcoHpm7fP8eNw1xG74t2KtVDSLP
9ir0W3Ed9DbBBcVUIGXeWW4ng0zFgCSeY+FhsBZsxtP7c56NM1tNWoUDh+hb
zhXBVt6xpf8pcedC7RKjCk5Qsz4qYIbzUUm/jhHpcczhQS5LkfhTvijf1z1+
z0HJTypJbfcDw2uLKbCekQVL8FdoW2WGWSusJjCYeSqcFw0uvie/Thh5SSwA
CWCahUSPv9oE6b5aNTWODWRpKf25HqtkFMaekIEAP2aRXpq5WIBFSYQAl1ON
F3ZWjzEKDQuEZa84T9AhcUXR8HDfuvzr1s0+N+eCuMRe67hyz7QHPbZXDb5N
rW4udS7PJkkOLm5/u+MQTKb7dj6erfNCrRTqDS+3XMsT9ebwgtIKaPMyf/ve
7lpyE14zV+nQWg4glfE1fYsg4eBqt7Uj5h3m6nfRoEBrcTb+wOv0nkDI2iiA
pTBzvSe0qaXoc/wVwTc5LT9LjydfXzwUCljeCoPxWNdnzyE/YYdC3mwttO/s
ucx8L3Qw9nUXPXiLj6rQn82PioDfx1xG6L35pHd3AakFssmau56KeFQgXhoe
RE1vGYxuE14gRTbWyXoOz79YsOri2WBJh401yCfPQvaw3ihOaNPxuzD+mkPO
9ygdjDXmjohBNnDPaeRHjYLCJ8bJSfLNkLKmMp8OZwxaJb+U2wJRVBNyNNW0
uGbKi7upcmnHQ5JQL6ltJk+QxtKoWl3B/N+Jz0JaIGeJ7BBLXMRouyHoiBfp
p/0VQPZFL//kHz7obw1+w+nPfYIzozAJpE6u5YAr9wBW7RIJBF3ADWP2y9N6
0oar/lAkcmflQCRs9K2Dr0YEl0m+TrXPpMJck+h60pDVsUYwHytMd5WV+IF2
9XItbSzCiNvO4m86YoJLvZKLnceUpsJS0V6Jzoh0p5OhwfJaHro1dSdG+X8k
nQFYX+vL5k10f1J118yoy35vNHibjjxcYWwP5ErcjrC5T8BNjejg+E2cGYz/
pLGO51oOtT5VR02PKxqN+xc9l4tcJPgxTyukvIT9arr/bigC1p4hcDEZx8OD
BHIq58+/8plIVxPivhPU6JOaOpstfY0lmxGKwFMxu1OFMsCe/O8tzgRzz/zN
FUsbnLBGCUqgqenjP/jAGvRcu6EezNBUcFULp+/mjZGdY/5G5we78UWOYSdl
FVp2Ngn088xPyu6UoXvcyckKO7RctCzDz/KRQ+fwqunvH1bRv+Wtgbidm33O
8WUx6InwHrMEEsrOqLjL7ZYEa9wSulhrOjiW4IVB3KqlZ8Wq9bsACrj95dTz
a/QugJl2e1yvpbRXAKl4BxGKtfxdRViJTxf8hA19AaHi612q26hvwScpAdop
DS/LDUQmGhT9V7kVslFvyXb1xJEXxNCMukgqJyZOc1LuCPGccwjs7T7fDHaS
nFjAt4gwxxM6Mo+nIwA7dzX5QVVcHQxtdIluvtbBksXnuG9g18rQgnWQdPa8
rurcq1RPZ7RIG5gLO+W25ClR41OOZSifstYjW84pGPey2wplOTz7h1hpbiDg
16hK/AhaDqsxQahMSaNIgY0OaJKT3jzwEP5QU9K3EXtNQCfI3ayBlS4ukIkZ
Vm1PTEmVtXOtTkiNHY/pMKzJiGZ+SSHMP0TbZs2ph/1LeSqu1a9x8yqIyVIs
+zrR4FttLPNrlZiftpxFN4S8JtX+2hFJF45Uo1XxdaotksCyqwIK3zFkYTzy
b7CvEfU8pSbk8Y6FPNsa2dss6bEdq+JL0drhdcS7vE/QAmaT3+6l2vxO2I/l
v9GlRda0GF4ALMZ8NIVE9VNKgch3FkDo+846Kg9sZIwapVNH0i6E44d/rhG6
lve/xdYuvBNcGOz7prh1FYBnKye07Biv5+yvB6R2LtXDh35iCXHHxC29xf08
oPP6Pyzbruu6ovKMhOxgD4Em2VVckYwHk3KQ8zU8vKgv+pknO2OpeYeCUMvt
Sm5b+BH5lXTAGchKeVGYssXiRtEeMaz5sMYiBBtE0/WC9djDV8q7oFEXoKF5
fhw7DBfpMYU4bPwh9iRwY1w4KydlZ7l0UvKVGLTTiDE0J6/5+ggLMVgJkyuN
sktf1BS9LpY21CeKAi980ZhezrCQhrzB7qDvQtzoen3h/KrEDmzset6G3kdU
zFeEQJCdRgsTR7DXgDlSbimJfu4V6pC7zUvB/tPdZGI9+HzZXzQGfq8qs4Qy
POTQyJoVzbM1kwRtCfPmIKFBzl2PtMU/1r6OrPjIZ1MJLpa/frP7tP/RJTkB
Jh8PeaISYceFGrfikXcy9KaM8tfU+FX5sNVjXRJPziWP3Ud5OFGcA9NkRrtr
fcR17Jr2CePM8kWcPu/s93K8wcIxx5FfyGeL212h4KMh4L9oebQrPafQeSU7
9N1ghAqYh/EQwuQ/JyLpGKyD0wjT94aAYvElklpqNVXjH6XZ9MFXuDJDjj1T
wpLlApoXJfQk506UksmcOS98Rbsi3qU9NqC1C8RPoNuPLSFGuSezsny4gyLK
INGvXCkrfb4U3YEBZ1qKlZGROxZcc0WbVs081VvXY1QVkTbw+1GEL4VG4WSl
28pOQX5WmmQSjW7x80RlgGYrw1B9jhyB1f6KtVj24og3yyKKQTgF3OysX6PG
cHNMPoxVUMka89uUDdoqgiLBhwcH1sbfoy900WROLuiZGZNkPVfKidJjGnM9
l4Uyre0f5FEElpKLL/RdxSzBkdSg8CMlKOpksuWP0c9JZTBDqTtm9Xmfojyw
osabhBok5Z1YYkmD0dgMBTE4qVbSdeEzVZ4PB7tEiZFCG2dtPnrrNE8Ykaxh
ukcTCPJyBfng9GGiYsRDvOhTxf+xUhhZf3EpeMHbQBgVSJ4Eo2/FZW22l54n
W+xT7z+wg34uoKLjpRvjwP/gf6uyu+UMVOnTOE2wt5dIZ260WEYGAXjJYi6A
9h69xkWr/MqI4m/umGH0RHaqeMQSP79RjgXTckjOUw78MS1/eXkm2yohOfHi
Kq59SP3bk+ZWO4G6NfhIxWl3H8m5tP1D3eVZxXxaPr6oZ80a5DhgAJScqAY/
OF65IIH9bbeNsY5/fRwTt4KO7Jnyu9AO9O3XdY60sZVQY83YRX6wfgswcpIx
zYfOekU9UQvEUsg4aTKS13j5VOsuFLBstRXzl70X6N92BLLj01IAKugcKQts
OeT1q0IyBi3c1Fe1jNdmeohvjcol8NmfzxRm12IZ4L5anHBYL6Cb1MAD9ygU
X/8LvcKqjNKqDWc2rV/nhGYAoCjKIvh9WmrvYdFxxiokHXsdOzkjVv4o+ytU
mLrDK68C3lA5oX5M+DJr2ximGUJEnbo5F8S1uEFo94Q3ASujs2nR1a+PKlq4
hp0JppQig542kvE/gwouZV0Y6Mp0C8BB3Z61tiC1WTX13/pDN4BamG8iZMJ6
Uk9N74m1OndJ3cyC9BGIn77zRi6JAGOXRBuPF6vggZBaivko/8/rcQ//pCd0
SQxYd3jhBTf0IaiSl48a59ECYvHpA67XF5Dqs09nCaI9d03O5peDdeKMsGs6
nx1++BTLowJeXqpq8/c1PQgTr+TsfEe7OuDoPBIzdGILEBFrqCkmGao/2Qpm
imSlcxlV6/s+4Ni8PcJ280qtlLRc4d8264Zhsngke0vmGMiTm/cjwCiy6WCq
XRqtWmTeBJiWySUy/JWY4gmBpnRVR7MqDJ+XlaHTD8uHScYuxfgZfIU5cN7J
9nL3Cj5d/1s72Ov3rMZW9FaTjFqYG2BbHicDXYaKnzirHjRHGZpmDJMEsEHw
nLNuW2j+qf+sovVb7JAT1tD0p5kMxBuMiHj0veaog3x12dmOkAKWJXejjwmo
7OyWIhnGzzSiovrEx78kECMYwEQAT9O6Vkk10NW5WHFGyGcQW7ep9gLJlBPq
RW2P+cbfOLMOmlGRQ0EqCKdxSaMFA+bO9Ek8jHdWLcHA1uwYx2CcnZKQ/OWD
btqYsc0p5QKAhEcjy9VBYi1w+9RzicHQpNUB13TxkVp+aa1PtMEtgSNXZ63F
NbtFrEjAALtoUfAhZzSYHpGGt7z8+q+zZTvoeO0nMf+Onnu81k3fzNRggOJ6
QTAJ4HmsVUJ+wXXAYV734Wp0FAt6AQIkusn6vxMnaaHVsizJ6G2qvdNQPigV
ftOSEgGg+ebGNTRu/RQdgnawm83OjpENKAnNTTJs37TbEQ5KsESeNvN7KMRu
fGCERd10ZQ3FJ1ioEyYf6JtG20SNQoTs3jR7/zkxMo/emuyYxq5+hvzY4DF/
CdXqMKgMP1AQjbgTa+ZdnBaa2dhreUE+6xnIJIJoFNdU2Iw0QkLI2YCvsFkz
m72QGCXb2/19g5sIazs58wKf7XuuWL4eiIiRlWFN98gfGern74F2RaV8tUiD
oBvD98nkxLfGz0czmIzxBNXDBnbJI3+6Fz6ZGotRcq9zOG/APFOCss8jgNmW
vS5UP2svsntskhu96A4klwaAdr+Ag+gBNpN4pE1JuH6ab+XYxsDM5xrTHDg3
CALsY8V+HNguvMv0JuVNk7JKT0Ohwt1nEVeBHHkK/9sFc2VvAH8H9Q1cqycY
WxRPDgjaPtekVLo44r7RXIaa3lMB+lBPJJDKJjOm2v/6oypKp+suSxpZ4oza
hWbgtXTKl8dSY54zG0YptrS6RXhDTfQcbzh5fPg9bpeRnvGYSk+qyQsILYvz
sk5m8CFrrxX0gdyPGVF4/hspWYbE6dKTKtQC7wNjuHJHzFUDRYoN8+oiSqKk
j13ZE9/ws3Va23E7RI1uP3sfYKSqseSaCwJbUl4uyLqrDmUlU6QyRPHqIERv
LkKp1EitECUFMLW7StGJy6hVW8GHV9lqnhOWX9WofQgfyfgQ2zylGWMejbhQ
OxdgVVyAEra80qqwColHfyW80SFtGsTmRB+uyjEDIcqVCVryrM6y8WJceh7c
LcTZ1Y9VSgKSZG+ZiQzYGN+HoTS3uCpXIh/qb8Akb8FfDbKp6GEy1z0lhtkN
/q9jARluFF2jYqMCba9w88R8eLObyMKpLnEY6TYyFcmIJq98IM7YR0aVVuZu
annlrId0anfV6+hDq+GxQd/n32bHmedWWcNLrNbyigC/I1yOA05iB1yPocoo
JhtcVQrlfL4Dz9U2y1ooLsSVhi+f1dUWQL7ZpNadoxjC2aTMxTscitobhQKL
uxXOX1mCZH8jjZxkBne3HlCL46FUwiWZEQDCwoI0Fk+Am8MSWRddz+D69e3O
FGztjGp/VckdRvzgr0yuvqI+Yd0oVnM/cAfJaKnlY05SlZtNpoBJ9/AOsQ3s
x/5sb36jbksok98B0rVUAUT3N+wTE8OYU3K8Sh2Iqum/2G98BV3TPY8bRwLi
+5JZEzRa9zqgbZFdtk7jtK+dAdcUaAMYKWrj8frQDydhJHGsJediL5ebPA3E
NAB1iyZiBv3xqf6ISPYECOlSFp4bzgmqJ2TIpqDLH4S2eaCBZt04YqsIrpRP
MeICq6oFdFTOS/+26qYmOEeB54MugP/zfnR3hf+rrantWs83j+n1BYFs7lJh
DtVbbmRO+efMIop4BlCc6JhMBb/aiGi01jgJlKXbYs6IrUIxZxbcfv7D+VkS
tobkti/OWsyzzUKMrcaGCGW0kP3qFhNR9KQ10WNGLt372W9JUEmFP1uy4/uu
SLg0kSus5zUzWSFY8oq2IOS1HxTJzpPVaF3Z0fY8lk35GLlfYgFhfGTEuea8
IIwxil+E425GAUL9CJz2xvdXm86uYkThn0ij28LKGbKE2a2/I6DP3gHXTxL1
igX08gXCGxRjTGHFuPExi7cPMzTmkz3NCOmOSzctGnJwt6YDuxYBEC5WMoUK
3sDJE0ZNViCYNyxHPuZ1VKiZr0ONuZULVzAZ0GnYQizxf2M4sP0WXGdO5hBQ
mudvb2EScgYDEKn+mzt5Ya+4d/wj6rcrxoGDTr0vbD775fMSb+f1OQU8WrKE
UFUi6kxMaRVZjzsJi0z3c53SfpXNNczJ4tnGO5cdBWemuHXN6TcxKepZCxG9
PHlEyJ3lV3RsXUB63jKaaoYFTU1aY2NYdsQVs3kzWy12lbw+HfuSPUCCtYzq
nfyTQ5xxj8TYpjFb3MvLb4C06jL8kIoISoIn6+R4/OH9bY8JHSiZe9m47i4b
E0y2v46+Yzl9xg21QBU5FNSbL3xn7yuEdk1pFRG2vh0l/n+1H+3NqgxEdTV0
Xflkl+htblgMOwhWt/HQjaAkLq9nUIxj0nVzhWaLZc05h6g/GiDCResif4Ph
lQrTanKmrFZxTlCQiVh6fPMR2cf5+xIjPt7aSPISCPvQ/lKKelJd41gV7YKv
fg6+KbVYGjBKOc4I19MyVWM5zaPQPW3qj8IFIxwmefb6beNfHHumY1FKqQNE
V6yNumfnwA2/cgIxbeG9JL6ZrgnLNojFODQG9zx4qc9QncUTAJCg5kZbp3pj
7gLl92DIwD4PeHMXwP1Yr15hzX8hU4ywE59Sl6jsRz08yUeJpTEHu5/XWCxL
YFF6mkcQ47AXfXUB/E6wdPA1dapcZIJGiU9W5R1E2QYtaK5JEE0hzZ06xb8E
+l84CqIQxqIaYgNcnJIBvkWf1aln9o3USF7f90qlpSo/Ue/e0jbCCIOG/6Fk
9i6ERB9IHJmkOZCyU0HX2qW3zWLRJBYKyYRfzuPUx2UmT68QnBqFbaALgWXD
udoyTm7yFVTnWQl3ZM0OTHSZ7NJ6o/TaG70dUWfZ2fHetxY9YRYP6xT6H6NP
Gg/HnK8KzVQsJ8Jrg9CfH8b2HFFbZkJHKPFZYIiwRJfAg9B0f3Z0dOPEr21y
0mSKAYrPWePkP7gBRE2z5EhOi9GhAwxLEoHzqODMZrPFc3P8obk7fj3hQza9
tbFpKW2ljsyzjtM78COEMup017vAfZpJlmHD0CyGXmQcuZfQ6161ndbdHdTp
wSZpHLPoLw6A2EthDzsKAU5OU0TmVrZQX/i/ztjyBXQyvUVzAubXma8tU7Iu
WXxpAnFiecaLg3rmzGqlSG0RyMKNSB5a+8/W5Dn2lD2/KGZs0d1yuKUXWBl3
icmCVCUmGOaWt3C+jqDYAsdvAtNiMu/qLwqL5PvRtfsvl3PtlKfgXcn5NYgb
AAEDaKDpuMj7lSM37qtCNeAtXnisFCWx68kWCgaPGQQmtwLNa/4BAxW4Naa3
4wI87pmGa57mQ3fRngw5QCm0aHVK8WyByh7W2dig7j9PLCOdQOJfS2Sp6K7t
81MlxBJJYLzmCqTUJfi3I7gG5vJgIUigWh8jGEc37uZi39z+v78EaF8Atyuu
NlJCc14L3qnoDjlVNbKnAhVSz1NeMkNIrjX+nbHr+AxNzfSHEYqUHwFANsCn
2T3eBhTAOwa8CewkQsVmktal0pDhEc4cwFEBVytyG/gpJIwD4MTWptggPUHk
0ydacCTNzD/mxt2z30ZLU3sFEBWx8D8otCZoWahT/AVIHDfDmTUrie1m2W18
nrW1NuCPqYuUMve+VgVIeayCq90rnZhYeZuD1Vv+t9opdAM6MiEuAMTuo/k4
kbXP8ozKZDmIanZBYBQ46bV7MKdQcvvZPsj62aSRx3tCKvZFKJf6gmJz8VCd
fPo0YKAc04XbgOh/wP3nABI7f8sDCOoKSDCPVtipxxO7Iyvzurwhzu3Cbt2I
CiS1jDHZSS3CH1Ix3NkbdVT8wZ414VSAbnRBnV1u1UWxCwnQbIexk2xHaJeq
mJWK/SdcTMUhuk953BVyrEn6Gdnr/BK67D/QTUBPdhzqoqzsgdhmZgfaHJRq
9kB0t9Kejp8RzLgJZ96vniB1OCJqsZSczCMayc1662N/0r3Zz+Ww0Y8cQdTe
oDKohIZ9GwWejC45QiWrchoEn5f8ZFaKtOnYLjLfiqH7XsGDGD5LAHimf8HG
NXt2Wi1GPs2Rc1isJz8tuaZFkqYsKfA0qRPaNYVZyySEF0a+CqxYEeBcNWnh
XQIxAPcA6IWEkFEQsTmErCnwLu3D0d/aUPAoJMqsehCZFY1DS2mN7auMurbl
wmdjIO1oEYRT7mOZIb57grI2cPdXtsSUnaQCuX9bwq5sIK/lO6PVrzocBryi
AfY7zIyX+yHFeb7yZDdhrdv59BcEVaox5aU70QHiYeIPd//28HWQl122NbPW
KZXXwaP/fD7N/lqdc9AiBj0zy8Og69B0hmEZxJR67erSBFS7Tl+pUk9wLXkN
md70MIV9i0B6nkpdyC/WT8k2v90/NdQcQwnVOHYjrsg+wxnKXhU19D0gQt9Z
JiYDXJ588dYYW1Qp5sRZJKh3/K22VyI+oGO+X+DTnjMDH9ht5e33FjtP5q9e
WsBWjq410iZWLjULQw1wH/sgxmw21nVemLHbb6DMcYBfFa44A5NX6bYZJz83
jq32Dquom4a4exucTbDQC1z2JCh8k0yaBM/86Sd3ouXliccw1VJpo4XNwg9J
GuiUiPNpXAUgFeQtlJzcjpH73V4Xponqmh/SbkJykNaDLp+LTZi/HN+kdG+0
C262agMvSd90Q8pfljogcBlbxbSeeLBq7qplDg8RuGmiZHBvZeYsywz6INu0
0/p0em3+YqlWAz6Yqs6b14D8/O+R8Hr+5x/I4VDN2VUqqbwA95R8ypDRApXX
K0j3C5roeuttOCq6YUvYudlwYbohb+VrIVcB5VsVrYKHFYCFqgU/W9UPCpk8
mYSWwwIYnUxMIHdbJ5nSLfPMJBTYgNKTzPdLcRHszT7/HtzzCQ9fVyQ8NwOp
r+RJLl7iubpbleU0EumHVoUwwBG65ojgeMGyCT5RQHzx35JfZheqMmGCiuYd
DfhsRdGODTurfvcQQgc2by06pxW9OqLbLyqp3UtbIWpK1nYBD8O00Q8NHVdI
Lv9BFduqiz+OGPRC3HrUDK/VdYmbbihiPSeTCQZnV0n3d8KRjuJc3vxnFBvX
/3wr2aPmKIHVhrUExPiugaGjfmxXO1N6sc8dE0uNimC41uFOQKulSiwVizRs
Cltf5FadqbKpi83gD8M0HckeW4mOKfBzsMTKKy5IkfbBJYDjHMQsYnAPpvOd
9CZZ1NWG0tVu7eYPAIP7zuqL2rd76iMSH6t/YWO2p/gsF8lCtgCcOwHnPGjm
/LQ+kARSixz1M7u0KM+D6921CvDy4wIgS2VXU/8Y/2QTFZUH7KKgVBANS5q4
mGRYeMExrUrTUXpDmwDy9hoG020WqpECUCAYeuDcmcQwJMAgxzfWi7VYD90e
yYX47QgBdPqebjQ2cSk6O+WjrCVIlSCpp/IXa3s4xHgqcYH7qQU4BbshkzgG
beBlsuyKo20bijx07N5Jy91CFj8DsUAaFz/yi9jssb9M7KN2+v7hUYQiEeTY
+wAiQDDdK9DzBKfdzxeG/SAAaBvOOXrVuw+OmyDAgfzncyROT2mv3hc8wqBM
dmCV0nOmYQJ6mn01K+ugstGHo6Zb3fveQGyz8BNa58vy1YgcqdFbTZqCBcSg
UZ1Ro+8X9ap/lBckV9j5ymlmuJbYPZlN0pc+I2iSVAl98FcD+f5lRfZZsYc+
AUpMuikQCwS0mExXU7PRzT8B8AKdryhjMd6qxOZpWNWzkOSPCyZS9riJXMIs
JO7yfu5K7cbJ1LG/vjnKDi1SQX1iT/KOIn/95271PlFaSOnpIkHTKdqpMyfg
PBSIZDzVuJU2S53X2nht0a2W82HcbSFU67PhIE1x0uFouayfg/rZeH/4AEQd
HtNkEUGFyZb3DscmFE25Fpa0v/r7dtYQWPnsGGhthAsOjTksXvN0Q3c9/xrk
N+sln6G3aaogx7TnBG9NX3Y9OG0WbqS7MM2Gucl0DJ2zw7ahDpLzXlImxaOT
hUfj8EgCqiLw+8PDAKxsGg1oI2Ch5q0W+ACzHjcJQcOXyMOJ0dWOMxDLdOLt
sx7jv6/e3NKE0Vj5DYC/k56Kp9b8S0PG3H2HLJFFmYpPdbJnBJ0f6QkzCKGt
yZl14FMSviB1Ro/0W/RodpwLohYXS5+rcmin3CVqm2FiwQBual5rGLJZJR7S
1pcarIFsFA1NWxQWE33vSdcjPZF+tCeNIn8LYgoSQQZDr2TNb91EdGissAl7
cXNLPkc0IAOrTyJr6qrjd+/nahqWBq5ICPDV3lm0qDtRVmRHenbal1tKHX2d
x39mJNTA0CZ4qnPPrb9BCmdEqYlS2dmTe30+8FTeoT/4E6pQN4fW8ACtj8ti
tzMynylxWp2Gwe1TKckztBAgNe6O86g180MW7zJXSAZ9FscJrHvjoCA68uvQ
Sfj1BktdUhHHIeRE3+HkxN6cNHBg8rEYNLH+MUXet7zLEbIq24OQfr5WxQ4I
7onsL0FVx0UIhILpQYss3ajzijyLatRQb3d4eM99M3IV6/8mebIzR9DHAmVB
gjQNFBR3v1D5hEHY8jPG5pBgkxgARnJU1c1NxO83SAvVUGoJz3mOab61c2kN
SePlT0VdO1VSO42HnqETSmoS3fj/bL5h19p0ZPWGZDiJBJnOW714Yc+wezUF
PWWQ8EyRgFeI1XK4gb9Ps1VZe/gPlATlmt0fklX44CTDPdpBwxLK0giXOhca
2xtXDxuwrwanqoyJ43+VaVaYfKN94nCNoHHdxxbmvJzaLJ7PbfGynJtpUvKv
9t1yhhL7a8ZE3JeJb8QcCVu0TrKJIbI7dZb/XUrni3TXCakV5W+Wjn2aDQRC
vjE/iwHixuUQs0QGgTGDBH1e7z3rrubcXFZ6af7ORrFFVzr+r9KTWJ6+dWiI
VsqqMNuvaYp4QDI3mejaJM2E3nplk0tj+1WY/c/GRDuC4NohoTEfqJ8Iq1vu
UaJ8Tgl69ZeWZu6BfnTCjTwuCXhswuK2MGR1qmgFO7EnpzxJyteC4vtwH+nd
ipqFhbn1OVPTO/kFCI+Sc9aAYVyGYuWlbMWP7o9V8mRdSJiIooZn+1uAwNVo
wNT/8uXroivUCHf0NXApAU8qzFRn4/hAwEOaAe5cbBi1XJ7ghbIoY1gClO+j
JoUFmphJSRX5cDeO72Nk0zzJfaTj0xRnTsgDu+zNAkH+gWuxd5K8emmIbCwT
3OojVqDH/s7IGd57HlaZrJyYjxiUFrMZTGHnT6ptYdXK8RTgohllx203owmm
f6t3v6nhkIj1LNfVL1+xADh/5IHtbcsXDLHDBZeDovS5vss4gGb9QT53BJvF
6vhL7MK1RcSgDT0cmoJkyDkTuanijvCAPC7etArqOx0tgW2BBP48ctfMuT3G
azS3UhlfFBAGoTJhjYYOoGryootQRufCq0Et4I0WI5H3N0+EcGjzlSq6pDoM
mNJNCsRRtqVaQm2891HxAu1JvZsV9R1Ec8nXOHvIduan/W6I3PLBIvBgggTr
hjYfnM3cdnRlBViZoNKdY3IS+m1BsfGgivXaGX2vQUfIYRX00FOnPESUDXhP
eOlN6WRraxNYM2SPsAsOOhVzNq43aUwWjAVyC4CbRjhI4ZpD+w5KkQi8KDmc
VURw63Nyoh914Yjtv3Kr+mxtA+n10NZCz3menih7LGZ97Kybeuc/xpiWAuJ5
BmlzE49Fk2XKHceU8BrglftcifsKjPQf8+0swq5jc55PtgLhDjTktaXl8tok
gYCOWbcJX1A/wr5kvH085mz0rtcWELrjh6vXH8vUwRXCXQfTDOasaRyMZSry
Vpwg/KAhr/AJg+IOIz6Zld2Hr7Lsbe1/nkk8v2mj3OE1i9dCPP0bVHA6PMVL
G5sug+3CGsGJ+hYyUOZj0/Z/nWLz/uHKENJb6Yz7NqMPfSCA3r7lqDzEEmT7
pXZepb9WACrAkeaRu3rBuNN11o5VR5CHnOShzwQ/Iu2zuvcwEvTKP2MD1LmZ
O1RisnxdSBeDCsIJlD/RfP5V2WKXTJa9EuKTCdtN3Mt+z7b7FcheTHUhHcrP
jO3EN7DJ3+8UGG9G0/NssnKY0NXxwfHWHg/rOWmUob0cXhPMZmUHkiaiwxCB
nO9cCsH3ouxEZ4JihYquJC7faBTucVreep+fl1orudhcdBO9KpB+3GNPYUn2
uVTf6XFF+EDIEbq+YOUiQPkfqwMjDrYdG9SEr0G9L8nTY8J7hENNCEu6asC7
0QnnlhZfGWAslA+h5uguuUn+ouCkWetgOS0a0kt264XLj/JBXB40JdpVcXN7
ssbQXiowRlHFg/1qmOW9MM9K8Px3kSr8fR6TX6PCuXuksZPwtuh7KAqKMFsN
sR1YX/fJqUPgsgLIWh60xyi2t/Ts85yFUTthlHW3qaPYNF5zly736Fs1FHnl
NfNUbZ4MXe0caoYdesoqugmToLg+H7m/GnSLmIvvnkbl6uLp1x+bOyNiM/aP
9RQ04fLPY0MEoNe0SgBbJXtlfw32Ut6Te86qiPwegD1KGwOVLK4rQ6URSicw
p3WpyDjKDoodHGDVNr89WmQ+Aa3jWszS1GC1un0LK2q6rbFbW87YkbYjFAJ5
CQ4RyU36ieIejaQuX93Ib6HC4jJGd++/v+jTiPKjOUEJObeHJ0nACd51myLv
sDeRO/GwxhTWSaW3Dx2pgFSDu1SOJNTLxqC7fQix7Wg8s3O0GjuAPe4arGHe
ROr8wWXYnNKza0J8rgkt0ztXqhIvCzoLfC5QsUxx0TZcALhRq8uen8VX6eeK
Ho2WmyE8d6SmccO1oWAYagtXqZbZhlmsaCTy5i7VAx/nFgr3px2GpYZQ5LfI
WW79VXMTP9tr0jKr0ETfgaAEFVvQI/C1LvynrskNCjaFmTsFW8yTqwAcg9dU
CD6ppJ/vJI6H4ery8bk3esBTtlIVKEhF1BMUfqNsxloQvQiQBLq5RfGGXh88
6mARWVYIT08yIaq5bkfiwlx7tdv0TAAQ8c0yAcB/gRKOnwBYVKXzY+ZOZBbN
6IOjuDiORRPAc1LZlt1sbky3wWn1wNTKR10ahqNU2oBy92/T2ddUkR0CwkEF
wiE4gICc2Oo9LtdeGZ7QmC7t35TKHvdWL+CXInQ/nXj+x//dgtyuyrZHT/rx
TWVRzwyuoDVYMPUk08TLt0jyTJVA3jxGpjMRi6q2FOCLCtmtkUaqyKPNc/qp
DKOXY37Cy/CdhWfuEDt3QUhOqx9Dt/WiCh+6bhgQDNzLcCGHlYunutlmSp0g
CPT0uo1VQqoHurwnMkGC2wu6w++U84pjty5eKLrLN+1Pm+5ebtJszfFfKCX3
7rGCHpxbu0PJM/G92T/B4xyO3+uq/j0P7PTuv801lyKoHElpKxOvbLjwsytn
+4jcAlPk/Q/ax1Ko88mE4d33hStcyvWscSTJgDklaPRfUqhSlb4RHLopoy7d
GKtp9Va14m8hryPEmSLF0+AtJ+gVF+KTd3FGg6wz46P4dNHUeYieeJ9/4tDq
gndZFqnWfhBVt+EsETXDlp0r1z610+Hq9ajiI2jGr2bRj/bOT4XrkI6N+KVR
1BDT6sAQ9F6sINnHhQ/4RVtvj9N+LgU0ZS0R4OFuxQHrl/q/Iz2rKyYkK3vm
GS8oV8ykUFfLgJRMFy5t2wkD7CrZ2WR43h9sLfeQPNjG8tpuAzMSjyRMM42U
X/ekkwzNCRpNOxwcoG3VJ4UXjW5Az56T/9p06HtHxjC781TFWjwTfKRj2yCg
7u/YvB+7h159Mu0cVLOOdY7mrEUQd7k/OrTpCU2CP3QKgcPEZ9D7HtrrhgE8
vcSVRlvCpCvRXN1mDLgA215gL9QdnoYLZrBt0FzAYFyC2Mj0kHSzkrUtl7T5
tnLGQOyepHPk4lpia1uXWw4yqbZB3IF18wQ+9/PR2k+mNHlATGcjMgI1lBP6
koHbCyl/Ew6eBO+kfG5fb7rSdFCwqogQtsURkETpmrBGRWl42sBi79mpTYwt
WLY8XklVcleu5ptB3afxgRkfIcXrIeI5lKrQEwJtgUxZjheIomJqS4h9x4eX
Y0eAExsgEw57G+VUhqJ+f/GWIEdJHsd+7F6mdd2TBY8pQ1g78c0GHgQli9TF
bQxf4ENobroFP0F/wfyNwBKEhBMqdW84oiauNbiuq32IB41o8QuJVMo4N78l
OjzTGjkEpurE0QlsZO9Gahvdrmi/OPKyf+iiPRVjfGzo4L4v6chTIZrDKRiR
eC7No5EFLCxwlR8AetQteAIyGOeCfRGlh+9wMEa5LH3uKYxFX0VQVr+JhXzu
WvFT6Z2fWYffnh3WJ8pI1pBf6kux05NSe1v0a8i+03NinuLvKlw8WHdDUE74
BqPGnYITh3G/vOoN2ct+82vvRgPwYAQDUOTdIyCcx9R4BZP7vafolsP+6uqm
8sAhTGeeXOcx/nVwpTcgfqB+q6h5B1yHgAYeTg15XFZvS/n5/HteZw8Ie/8S
hObua6Aut0VN4pgVibyGDmvrU8KANW+S0rWfoQkkcNj1mTLKo4YIvBhhYRTY
zaM1vq7CLPfuERNMqe/7MA55H5iIXLbqCmulrD3i3/v84g5mJCH58KSE/xPT
CwstblJKo8hzKXnUrpDljl77pir9rFI6NJqILTQPYHnGc+3EnDVWF2ME6my3
Zg7S83ATngy1RsLDdaP2+OIfiBpvE934QuhztB7sKyt7IuID7rfMM5umiA31
MAUgqGmMgD1LmMRlChMsP19iI4reQwC/Ga4nH3E26/5ajRXCG7UCDDluAdpr
mrQqe9NWqWqBa7JZlF0uno4kDwv3Fvd5yW6LplCDup3FUcBR1VUYU9iKqFMC
MdmqGqmhSgPTmKdR64cFfTJSZeQk+DP/wvFCWYu/jZbyZiL7zRB0/A6NQgJA
uMQofONHbRny11O3SfRDgBdQ/14I3H0trCl/NHT1niDcAUuIfTcXUjBMYYzi
tKHrY3oyew6hUoA9Wqum8tBw7eA9fUdYkczF8AE2l7ATXMi0wE27klMziuhx
UYZgY0lG8JAbk8OMvuSGcViWEio5E3+xumZXm+tkKsPZ/6goDh5p2Y8g6vuh
tA8id5jIBUFQGqs7ml44cFSCwDRrVXpuMyN+NiI+Q7xxIxupVKjgk9aY+Xgz
q3bBaEskR681M5loiL1K8Ckpq2fLzNuZRPZtEeXyePwXF8haq3pmFVk/HYJH
9zSLZ4iO5Jfnp8l31AxymDmsvjsZkh6e/b+tGYOeaW7ayaM9r9DeCoVjITJZ
S2mdhyJk5Vq6jMGG/ANB0c4gPzhttpJZ4Yx+n0SjEQ3HLibsm4Ce+tOHq9Bt
QVmtnv9wQNA5iQEz0ECa6Q+YPDPBRTQ/YCeMTtc71QsI3E3HJa+i6YYf8wUL
5wtXuCbPdEOq+yJq4atZeHaZpw/CBG+2xFXHvKUw5nKdgr2ZyovmN0IO6TGv
zyzdGXekI0X3NDCe4kEBJntRDxWQ5FdEPh3wNoqqbtIX00XgFxwkDE/Q59X2
5ExM66AGGRYGt5sTKTQV7AM4ivuKu4JdwFz5xI8qVYC0ht0wpzSGDLNSj67V
g5iFBclgMtCW2UNlWBa912ZDWJsTB4NWjbs6TjHbzkZezcaph1AQYXqGIZJL
SKgVgc88hvPUkCf113K1/5Dfau+MnXMXPJCi9rWRpYp4RPryQjgigXPrq4qb
t+gCStTj6YkkVZdomcu83guNjwBGg4CzHOl/kb5VZblCo4cXJi8RXZrMZtkT
dJRKdywMFWvU0P0drX1AsoEGl1BkTUoWhMMGu5i5iBAeKMvBdFBkOQ1sDnub
pv8xi9lm9Onjg8N/3G5BXWmtuCOthjgcaria+UTxmax3Mjws9OZook+hKnbL
i/JwoAs97NH0k64DkFcZplkl1BB8ebUVCBGo58Rhh0xcG8+VCzjA4F5pjf6m
xOnloZemyqYcA6HApTFYzjhQihoClirx3I5oFlox17fhn+igi0cJAz2ZAIvZ
45JrrB8CoZ/qd9eE2nSXWm6JfH5lPUV2y7WYcNwldIpg2im+Vivy0O0A8Xzd
YaKeFYKSiuuVbQt/2nf2xpkZ1k0yKj5Ll5ksxlABBO/r6CEBK7Qh9lcqN7qp
zxnt6hWL3DNRrGKeodyfWtDch4r2SS25yiLJ6Sih+d6cvWtBWF96CZJJH7Mb
jjY1iSnC/cJO2saeJdagC1hyifqzGKrR0qtmhfG21Nzv1WFjVm6lLtwSWPvj
RPClDcBHEDSQpTvBSaddyJvsfRCxl6XHyEXOMghzG2dD6CiAhhuaG27bU0gW
btEbK/gKlnHdPPvJ1VF8V2YcOdwE3F4oLpiwKBs8Q7fRuYY0npLoyKZ8yVWl
RL5vxAqEV2bPy5GyvJz22+vCiz9LUx0unIFJ+Wsh3ZDf/GDFLNXr51R3fw+g
UCI3iypHiDtCwYomzz4TI1R0L0zreXgJr3bBXVlXytfFUJu5qR7AAlXD86u8
cUFWZFSYGKAI5Sxgy4bA8ERwDJPpt2TF4XpYPvpgeDeNtLROKGAIwzZOlkeF
WsEsPFdOIucCjen7uPa5vZyO23JDBEM4nRPQ/9xGO2rdI2O+SNZj/gHNzXdW
sWYXUBjQSrQukM+zU1ad7UoHKiYXztUxPfZB+zeyg2Ad3+xBQ2OsXAea4jQ7
RAryKHR+NUw6HcshMb7lUO/oCb6tr03RTOOKmWrSy8Jb0uwUtHYqKChyJtVD
VrLJIFnTo5qqlkwOQBuH3mypTxD6VV7cRGAbdl3sC8+qQUtReDuMH8HIDMbL
7ftT7ByTK+lyM+I3pXtGJBXId1afNPAqDUl1DfkQaUY/9cTQr4wkzNu+JuVg
OalN50TmFWAMkTGdELIDYcHBph/WcKAeXm9BoQ/+8cfF3oKKLMB48TgCVk9F
6Elh/v7f1NPz1efkAqTH4wkxBCqWrHnxNVMJ6zjY9siTF18oTHclobtVrbDa
lsH+IjT3dsLyevRpY79pPltBpoJq2IaNBmcT9adPfdT2H095EUSOfdxtfF0n
H9QG+Qs54Jq0k1dkR+vbj2ct7MPBVd3qy4Ezrs6jV5uOVi3VR4VGY74ZVp8V
N/6ilQQTwkA75GTOYzraJHYidhm/1K/NQ78xPb/69uchKNjKVCCXMWfa/yUj
+VaL+xqyrsOBjMeD6EQXWDuiEAGMOMMyg1NCD15CYRIEqcPxsDmyM1HIrqXM
JanidFGqUNcEVz/xo4+gF+5NWOT74aXak+qOz8f7gVplacZ0pkErOjGhSBtk
cXhOMo2/eONKnmpJBaMUNfK0Me3bY6CurEPGZEvMKFncmFvT52czcoHGYWpK
mXkF1ASsoPaVqSTwICVVWcAeTYhNq+KrCLJeBF3CBL5WTJmbRpODIcwdJgpk
UHIgZnE6wZjEGxFvzxIC3zfsFCIOhiPptv5s72V5U8XXmlNRX3Llcw9NqzHH
TNkDKdvk51+DugmSHacLqFpmaq6u06eJE9BlAdF7AHwnwj0AhEovJsgummHK
dXs7IAoJrMzDJV2TRmSQgzjqNvDK3ZQlJCDInyD0i96CwuJFLxBEl9qYzcQe
yHkcDy6fPTTQFQ0E2HStwLohIVcFW8anAi+ORfN2IBLxq8pej7yRsse+AH39
9gxZS8Bu++WnZ/uxRo/DBMe90kgfeWeiofc53DRCjtkOglqbmajd0RMlbeHy
AUCQfDiAXtkeupSVkTI2lMVuh+bHZleChLyDrAps/avyMyzzGhOTjniX1DFr
y7Ssowt6V/CvJn/0D/ntSeJafmNUzuvO0ZyvECJpJ3HAAa4dcabsXjdn3MVC
v34jcvxP9Py+OM3lib3Ri4X2WeGaNuvYgsuVQwt6cUUshoYrAtBUnySSE3Z8
S74x6Bt3oNPZhChfltxeJvmbG9iauDXwGcIAsUwRj349EjgzL8VdSdZgCsP2
ChjRs4SwCK8iRQepcokLqu8YcE6JDN2rdWXWonqFuD8BXPSgfT+9FsJDjkM/
EcK5J4bbTsn36No2EQpEV+CNd7ipPzRuVHdCmPwHYt3cMBN38z5mtfbrnfsp
l+Zklh4Piy2LJVRSmjeLBEiYEw2yC0gIBNjyopphFb6+e3HSnC5klLjebI9V
poIkzfXjTIDOKA/z09BxlbeFlowGXM38hstbWFASy/lqA/0H60bPAX1aT53D
oe054ei6oi/D9OLf6xfzfSMC8ePtkIvawJaeiLwcRhiOlKPgugfcTTuxt6PX
SwrQicof5yj66dUhOrNZnf2RjSC2mBmJXB9XbSPzb8zG7frctF1aY9VLjAaR
dlPuc24imhWQ7/iukhUKY1WYoqxvsDl75dMtvh/v/BJ+P2/eYuSk/k3y3bN2
4BmEpPcur97A1/6oP0vKD0QIv+eoR6DdzU2owXTD8hNdtyiqtO6is5ZDv+YH
RfrZ7SIx2jxZhlL4AIDruZhuvyXZ+akqJOfrpdSYh08Ree5N6xQ4dO5IIDvC
2sBLeMfVskxLWfYTHgd4HN9fcINO9T3W4kWxBdfX59TBMyGmW6U7R3mAi0Qz
5jCx3TVmjax7SXE12QUNlrA4Tvz6xNifYzxpi3PEUu39EPNgOBkLyr6BVMCS
uG4M5bxVgfO+hwEncsfGJ3kg1CVkpDdm7C2Wj0AOetjthGd+klzFLF9pB95f
DDGDx7rIOs7ftukuQVCPlVI/A7jGFsOhy/HA8vqeiAexHFcIEEoqbTctTByO
IUv/6LdaiRVLFv4uwuYKh7VjD0wNmBtyLLhdkyV9EK3zv4dHq9QqwXo9XnyJ
w5175FhT4fK9yx4iYARlW4NhgtaACma3kz5w64+2IjL/GeMX+q1Ie07yddri
SU8V3TSO6f96i3vWahZ0h3IiRoUzPjc+Dli5WI3kBAJCj3oPVWTtU/jmDbjH
mIsLTsZcFAU3vaT1bCr7+lliPzajgvnAru+1fAlpScKjpB+JNWXNjd7aU9Am
I0w7n4QwswD11UxoyJD1DRpxQirK2DKTw2BbSN4IVD2wsUGn5vLMgySCJ3/u
lc2f6IdwGGWcElOKMif1n6GGlM0we/gx3Dqrc3F9YSK7s7VKBFIoraCe0RgO
chUsWUi0MyKyeqAgVhTqUA4T5fNXeWWUbXMBzRIstOtjAQbkJ0QX/MuWh/9X
3RRafkTsjpotw4Rt0/clqRtndbZuI1dZUHZnf2LOCErijYTKxLRegYYzkwc6
TkSVXtg95n/DD9/lNP/PO98iejfhotUxF9SIrP2Vl9oWZuFJSM0bHpuANsgA
CTFxUNRcOThYbaGiuabbZ96wCpdA+KBMfJDbr54R8snn2FhtDVdpw99C2m1O
0eeebygQJW+1Khfu2g/qV0QjRDifXENPggs2aRQOHys/IXCR448L1JBcG1gB
jGvsI5OcvI+QRB/PwoNJ9GA13dxKZuW5wgkdMU2LpqrivFvKmp7VjxCtsixx
eNgBqlH2/lW6klwacBDzAuEoFPxkxZ6cVTDNoWjkDNkjstfTdifq/9BAeagQ
7hRONd7XvECYNQ3nH1eJCgwZGFb31p35n6muRH1y5RSmQazCk4HcKPAuGruL
gx5Yp6mOgMj6RQpOjCugA1xfqJZVKKSU24GL92ff2SWfSVtio0I++awBVf5L
trEVg6Uepc18GKCQnf58Tlua5O9fplPZiAd8nWrJPCCghTS/7wMJnJNyLhw2
bLiH3R2S4W8HsH0dGI4hdTKtvimnnpwNadlkPzzfMHUeLK5U9T1kYTqBHv5l
RzZtKHWEUfLqMwoxZWu6rWXJWwDj6bLSpLQ3DTxwHVDfUGOibgptGb8YebKG
geNIr1YYGoum2l2X5QfSq2fIb4EfR31ihGu1oSTX6MtNM9SkkLkCZlVngn2g
EM8QyLzCPrzA+F3YUPr09tA5FxaEVVW5C8uXqJOOC8tfKt+z879KkW8qJXB8
0dp6ZUEYuuFMLvLlR9dWgiZXgJvUSgV4BRDp+b9UeZ+l2a39ep1YEIRs0cB7
oNsBRjpKQsfkOxgeJg+TV62GbxJsuNZwdRoWPm2LdFTIN4npOzUGjUhC+FMR
454dVBNDb7g9Auegu5yo3ap05TTsIAf+MJwKRBsH3jDp4RLLODgP0/7mRs6+
H3u+8xLUVrEZcEbhld3lr6Hze2CynRw8NKhb2HRWrbtoYHttw2jHmkBw3qYK
H5PDaykVzF/6W5dHXTne6XNAN8a+AgcXj0su+dH3/pAituqG5oMuCO9nYp/z
V6WrEW5nrX/cksB+5vnBq96wBuFrz0n4LdM2VJfeogNTCXSQdIxJ2f/SC4/w
ZHity0ubQRmr3rsIvaM81iITS2fdidGh3OlXdAwQYrETYsKP6fKXBE4Oqyem
SO5Hciq8WC4nvNG6piv7x6Vb61mr3DjUh6QYy78HxgBTj7roZD9RFAw1rZzp
G9uRg4g+Z5EpwZhXa41WbupECHaxj+HbGavHIqDGU8DALUbCyRLfLZgcRhek
7G8IanuFHg9LzY+Jy+co6mX+vWIZsUCgPaxv3/vwTmAKjZUF+RPkzjRKMoiL
22u7thOuDza3efTWKuM/2/NcUaCGmRO7IBaEukDDVMDF6mHVjXcWvZxXZhBI
38bm8sjUD+lNZXfnori//KRxrOU1anmOt4nO6lLXzd7Dfl7PHwN0wLtwJNfG
LelcbXZx7TmVKNk09CZPjpBzvJ1V5tE2pPwaqkhgb2xzPt4n/r45HUzDd/Wv
doghkzSusdo15LAzJtlZMpFGho1BibDPU3wn4JS185zdAuEAH6/zHI4YLsBc
d18Xx0zBMAXqnolaL4yojdsot9RdSWOKAVzAk6WpHOJm4yr2G8Kj2TYjSCIk
inxON4WLXT33q7/OTPlJ8+S5+Ay6WBqzVvsXDz7EASVyUwuuloFXOC7UCOZF
aFNNsJZBVfVCjRva8tB2QO2qWhdEFVb9BnxWv1naWFBpzAm12aXWgcmDm9GL
FuItQuPnjWgftHX+QolHVYnmFhuQ620TCYr+v/O1lluORL/c0QVvg48lReem
Z7Us9GV10B8XT8Qz9tu8+rPnlFMa5FR2jjzDo9wuBxy6f9lSkjOo3f+OlcST
U2ThXJc5PsBO4iKpYMdlplbMhmz8jLO3Qx2CJE5OHP4e4kRvFZOg4i94p0Kl
vTpkpmS0zCoajWG2i8i5bySRWhhKn7DXvQ6HiWss/BljeKTAdejxWDrrk42o
rHmc1VI8cpYhu6ofkNPaFZv6GKQFAm+QWX7PFQLSs64Sn5/qaMxen7G2jQsP
ZEB+t0UfcFfPlQ742ikY0RdO+091MwnEoZEpr4o22tJbs9H8sVA6JHUVqc9P
eBdsY2cBQWGB4/gOl35Vss7mapVo9HQWv3S3wfvPltDW9wODiWkQTsWJP+wX
P0IMqg12IKrphWx+s6s5QaghyD4Qbp9DYm6zFZdWfXydq7mmHopqwIqGA3u5
rsxFbNTWbTdTulNy3nSOTU5PH5jfNYCQPEZ18BgAqS55HqyAq7c6KGic55W9
Im3yeoACPyFTnKGepJjH8DTsuPhZK9aBEO2tnmBWfCCOr7/pa6HTnve7wAML
gZFbdOym1jXMfIDcmciGZZ4pDmbI3zHAGrkIy41DfXm4Mkmqwse5X+Jp7QI8
NGLRuo4+roTF8flD02GwMdGEyaWNvM1/+qELVQR0B81kci+49jIUTeOIKgyD
LJxBnFT2fb5xYq6kz3w/t82vUStKS1J/x7dhOXaZp7P8cRINZE9Rr9WUWfoM
Jh3PrLnAOpWRLhvABwA/Gd0kYeCSvdByLKGf6s85jeV2dGTxqvBnmDVot/vh
dom7s4/p5O7bTV0n1D4qEKt1SSBhX0ThfIleeFBKc2SSymdru4Sw3RfUXoLx
529wI3jG9DHpCOgyEqKCU0AI9xjzoR9qfy4na+P09iQTeb5lFuyVS5LjoXwd
YGcvKSIvfdT6w9vYJxRM38mooEWAylODKWZwC3PwB7zCeXOTaYIpaFgK0Zw/
+qQ4rU5AD7DhXsJE8ApKp3r48jYpmVqxjP0viOjT0zS/hPiZV4XHGE9Qj3Ok
0F7yyq8jY7b65oFnTRRU4qpSUnFkGCmzwMpmafN6CtLrgGsgTN3CXAnvILRL
2y7MKaRopl+KAOarLmjN7PnxDwKhmlDY7dcc98al9kGEr4Lq1JDMoy7riHGX
yvT7QAe71xyBfuxghrQxfQLvGAQhbuhAa4B9bLGM/Whnv0lD+ABP+K0JPVpH
bndO5tVu2PsG93j/ofBjr9o66J7+o8xKd2AvStSrtqVItEnJqP9kAmcXYNud
hS2xlUmPcgyPMuJJDzuOsX5aSpUvj5ZvpOs5A11MHFVMSRVFfIP5aJkl6Qfj
aETYFMB5zs7eC1fQK6mAf35yCqnv2INI4kR3d4JJErlsIo038v7A0HDgnPYg
+caRp1kvwkRa+2kkzsWZxyhAuwbhCvURM+OpGBWW03ikYvSGhUIX0fZR4EBy
GcHKfRIHGkemUFT+Jg+UUo4z5lOpHBfI8TbSBKuLKR56HvMeKmSZzO1DrGYT
e9XGJsmjF5xooT4rWxBaipiMRgM77QGGjtS3GQMYKcJ9QNHNis2rxUQ5dSj2
KPs4QhO35vABgJoCR5oeEQ1jEsSevp4M+opTJToSo+6xlljF36kbDw84PYH/
w9A/K2ZaIm3057bdoQuiMrbvM7nlWHO/U0wPoWSyj76b9xL0haGpX7aNOlkN
DTaHkfXqINA6SBw/X8fK8govlvjOfT94cb2GJsNwQ18m+r2h81tg+s4F2jWt
9sQsaUrX3skOp6zN5bIe6+yKfMZ0WQDQOqn7oL2gt+7fIeq0h4i+aDmtx8f0
sZbaeVfxhB1DLydd28Ai9mVyUgwnmZqflYQYF6pOkm3FiRlFFXccag2ZHhx3
cw8vzbCOiZOjR8G2SvF+WnNFriiWIpFh802MWKmS77DWS637RpT9j91oYGj4
d3oqVavLWaAZUqSSu79yYWfMCZ02X4FLghExcN7TD7QSSdMjiV9YtpzCAf3u
1Q/s+cNVRisqtgx/TrOczTG7VcvBkCIs+1FkOu7kyWTrgr320MSS90GdLbSl
b4BAO7Nqt2VFV79tem1uq2tKEj7ebcnVjFFe72+KfSG/Xr4m7yk180g2s8Cp
N1RApyTzhK4W54+E9lsanBJDt/Sp0e1qYOR+CXBSfMYbAQa50/a+8qGQHWPD
crQ5v0jYGR3DeEV4aWp4YexF504Am/XsmlpPLLSjHVsHQKpHDQulstrj2S/N
BrELnShxnagM8k8O1/vx7kZl6EAleTOTL2UNzVSAPXQWQzGE7v/p519eqHt0
OoeJbmVCy1KjFIFIJUVPWahzSMpIy9xGak77w44EA8HnXi5053n1EGK89dju
1QBYA6YlcjUOWbGjuSk5gj7n/bjdeHgD/AMCqEdz072FKfUqK3w29t8v1seG
rSWp8+8up4X3xDjGxVBdsnB35WvKnoYz1eVsUPS8m78oVNpAzJqtXwgmmBsN
nsMYdzLi4001DiTNfjnDTM1U3cK9IFp1IfLjoxWP8HzhAWzkmeWcbIsYYgLj
Ccu1/1N111OfYgTPMcEUxpb+iM2PYkswfM0a/7IYFPKLCLcs4gMVXONYTw6T
JYUsa6StZbhdW+dpf/W7c/7YCmG2bpNxHWGeMLNy77Gsa7mlp2qROsKT/P9y
nPMnQnr/5CmKNFj42Z9HcY/+Odkj7VZQQ+B7KU5vFoMRYqJdAn0N4XYKRY48
nyvS//MKDe9EF2d4iOTb88VHFZbRNuuCyhrjMq2ApFRcyPKdhTYiYiTf+Fqi
Sow+5hn3ri+MrFgesnHWPWSL4B1lN5cQOC3OksN1U6nRLXaF/6x8hVFZKLDV
bErBc8isNFCfhWlGcb0H87pKxrHMlxzf+amCmwcrG/wd5a61UcwCY83vv2w3
so4CI4xNUxWD8t9Rru4G7yZBA6wLGtEwqDLgw/N51AJ1+AjUBGX3vsUTEhQS
+WYBRXygFmqC+0RCH8zSHPVf/KBGJ8gR0wb0OmfshWvRlst/wioTqW4JVH8P
T16IkdTnE0Rus/1rOlkve5QdXSvr/yzWKzVAL4dE/Q2711T2/2LXZvxpyI8b
jJG9p7lhLLjXquuO6mH6nPhb0RJZQ+MTNBbw+fH0y0s0d0YebD90EARerfeu
IxsDpHjMb/wYLYUGs7/QtpRlUKGaj6MsGAX3mM4a+U3wUK0FKkHb6SR4YVpO
nVQFz0gw20jcn3asDxKdlImYobyJTOYIYwSs5Df0Nu61dEv6di0xJbh7ezKT
Yb1SIWccf75pj+8WY/o8vNM5uEVDGt2lR636C4trdMqW3dda3QNzVLrozUqX
Q0KoqW+cnhJFiTrbVucgqDqD7iY08nMzsnbfqvDYed9sD26nU7LgMXXxn3rV
np0dAEW/VVAll2SJLs01/br8I2eDBsZJvAl9B+RVDrjSCqEBrpF/t4vGKFOT
+G93FdLatv+25ZvkMcAMH02AGXtaxTdjeRarVv+ymj0inuxmy/JCdCNRW1II
J18LPu2+CVtSs9WbVJXkNS7j7wPElkREoSPg8lmbY1QHN6vsM5WFXcmmksfj
4fK+aCwM8MTMLd7LDC/FB+eZCxzkTz/heVBwhtZleb97o/PCokiNLDMtdv91
OKoBWVPzsfrleyTYRKok+3/9GflroyqdcLePnlBVOjrEY9WjvsWTfcKubyf8
YdSRMxXpgBHxNKWIjq4LTbbiNKUNX2rsoPOf4ju9ZDZLOS8kMUycV0QyqZLT
vof3BGPoVN6wya4SzN9Wv49wWOmADQ4KUQycHEGdED98OEWogzV3ZkprNsN8
Fr5vrSkfEGCw55tHvx0WmohSv7YuYOCpeUyAP+PuBGGQ32wn2pyXWKm+z1gw
iYhSsdfcNIUrKt6X3n3VG198KTmP+YYUytQ/XmBb9OAGhnMYktlUnTFHMKig
XnFcl2XoBJcItrc+87SC5mi/+2kpBxGNy+vGqvFnXyiGH/O83/3s2mA7dml1
wG3SncPgq8W3NuPdg0okyvDTPeP2+SbpMEOPODMut5EM/lXtmC6RD+ELrphZ
lgm2VRhazgyJLtJFuYtNDBBvqwCVBmNIuZuIi3SLb985ATkzJZlNNzHezL69
DZg8JtA5SHyqWUbYNPgXPJi/kk7jzgC63aFbuY+kePXtwKCFaA/EH5GhYByF
27q5H7HT3lk1G1VfENmsFekdn5NSPiKZ5fPJVN9yjCq78K63hyw4X52Qcqe1
BAg+9Iu7UbT+i5VgisJBEo44dVBKpf5TfzQIKw7QjTrsEce+wXzPXrIQNa7s
PcKY1kuPY88IdVz3iyisEoroQteQdKIIBIGEfRJ1idwU0sAnyaqAdZha119T
NxpLAlIwnFIO5p+471TO7koPoBZ5reuRVaYayaFBFwzINv5rXLMyb9qaTDZF
0uSCUxo+6rnS8WWCdLs12zHcvkuvP3+hPd0QFXn/3TyDqKuON3Ay43pQqtuE
Cbvm3bddqzDbsameb1fVNqnh83lur+i39jS4SYVfI97l292MWaAviDR1FGZ6
rRmZrT3TH8YF5WjPYGXFAnihBa1r3Dxa5aL6N6DvxqsqsJeF5jsHID0nqwWF
NZtqqE3ODHuXk6eGyH8uMiPWWCySOqkHs+aA+WVBVduYYWyKUf7aGCfYg79W
xwpPsv1okErEUl/1taQg1T0Na+Mmy5YqLws2jJyct/TgxWIUV71EZod/N/IO
xlhnbqVWnmCHUAuDuCbTRDSmIybx+4NZJ1dOftxWfxFngnZ5kRjB6L1N6MXA
V4w3yjMaXpruQNjmyNG7LM0R5KW1QmCajinuUjRLSlBgr1f8TgAb1szjERLL
Y8nI0DpJwgGIzpot7NI8HL6owLjlDQnrTMniIAFq/0yRjoOqjUvS8msSzT1h
qHEABbjF6Hti1edNySTJbUvrQebdCmeB39mK4W46qkR1qxalJbfAQCx8F7K4
iXNBRDf1pCqrMgqrNi62W7NQ7oivRJgYN9N/MSyJTuY8wALUsHWbgdgn6ZHe
JQ7knhPiS39RVY3vwnRwvox7l3z6HFvxGUi/EzuJiuIjfzdBvg9PyRw1z+tV
hEGD4m/Ka+yZFSf1EzO+g4ptJdmzuxiFRUUWSaNrrb2XmMt4+4MgnnyE/aJH
CF5u7uuX+0qY29uEiwkwq39P0Rty9r1zOlJgq7LIxIYnTog3XcXGR+13r36y
oSdBmzZjzxO7YY+fbTR0VwT92J8R+RrZLg/0IswUcrfIROpRXID17vvbxeJ1
VgiOdzFe3YYv0T8IVyz3EuR9NibbYZdF39mxgghM17i7or08PNs/lZwi1/El
EUdPicGkVDNLc1czYQ1SgiVPdO9st4h5PFXtgV4oca9th5VKD+hxSKrhRINq
7Md2erLDRv6OaCKqMyreTXN1DgiSRMZiz6odY0R5TOaEvAtl0FSxXX5mSbSp
FpQo9Ggy9P9teNe60oltwqW50lPPNyh48upMugFqVJwxOiIhT2DNwy+BQVVk
6PeRpnerbG1WE70QrgYT6D88ECddN6hagAkujVdOKhu2/c9oH6ZtOI7mMCx/
aYzIMXCBcdozXEbZL9KInXFx0sSc8XM4fo8NQfa5hjRqq5P6mf9lfaa7x1Xt
GqxQzzGZ3B0FaM3h28en9uIA4oHjZhSk4jKfLyYoKazRBSnuqPVPyEarbpDb
+KafYcxKnIrlg0b01nQGE6wgt2f2aWbE8x0r6UMXdzUrObLxIh9LMbd2xE0T
Xu/EDX73MwjPN0hy8ZxMoX78/65l2g4cgtOP06XRSPhYW0S5TBZ81NxDtgPc
vsKH3EwWypFGTxygAQVRY12vMLsId0GGLg06RocywHRznYVflV4S18oFcXzT
HkL6SEmnEvZw/2QjqhmxtvWbREWACyl99V7Cz9u7YntoTeXslWmj71AOlqCD
pFQsgqYcHOSnR64dwHSqir7hJWkpU+1xmnEf9esZpcipFTy6u58NBLnjyWYW
u5WPrD2CsFj3vtLEF9mVUpFtXSYDg0MEzY96UY5jnAiYM9wmTAyfuUjSe+eW
hNHY2QLpUrp33GELpybPxrMIzqcBNllyLlNVe1GlCKJBWe4JZxpHlL+Ai5NH
x8oEMPCLsr8hvaIWeFbklH/yXOd876ODZssPADfezfCwHiudfXVqwtDsl8ua
TgYuE80lL8YuADaomU1ashsdhRhKeUgxQl6J5pNxdvifCjrpqZiPfLfsyswi
L1ZkMFLqNkgSVzb05L6ZzCyZIZGfLbyWZqqbDRWZhdC/K0c8sqi357UEnUgT
vjiqiV8l4G9U74acLI+j8jrh9DDi6Rr69m/2PZfVUlPDWSg742UoWCh2u5Jq
irdPdYSGeDpcqgmVmcH+HGg5FQu3PEW0ULy4Hcw8c6PUp2lhyf89CiG80HAu
hT0DKr/nxpmuLEXEEM7b4ZeT5ErtuSCPLer+Jkeod/DwYT7wfNQfVaDiCJeO
TG1pSH3yPj/YPkDxfp/tENfYGEDd9TC5Ws6Vmz2el0vU6+KAT1sRrxwoLIVu
niPiUQOujGsblh0PS7websJs5DrmAEfEnjAixQmU9KwhLcUB7sR5tP999y47
nxG/YlpSQboWcoQc/VshWytGBfQTQraabU7hFWC55eoSOwMPTS6Hr2jOj3id
OCSao2NLIzawqnuraBSBX+SyZcC/TvR/U58ojpLGabjQpWgt+XqB9llp/4Q2
xjTLbwxVjlR+iAqqOncvC+/9yEUqzRGQDY/hMPoqzS2A93Z3lTKBk8ICr9nB
tCTy8aup2qctwpSPA3Lp5KckM3vRvkKetq9GhvMm9PxvQKNRgVX6T1oVaM+9
2dfLzI+uH4uVRKbzUcsIw8lf0bc6qrShP5rknPQN+5cH11PTA2erNNR0h6Cv
B5b56VaLgaZtTpf8DSqtdmHAI/z4QZAkz3/1mwJXpelSAfVDtZovkjwAa6Y6
MzsJ4hcSrjA7vfEJTLkqd3Ob9Fih3Mht5sXqhbLfIx+mfievXoCQzM+vSHWB
syuYwXz+02cBK1SIz0Lk77vFbR8B28Fe6bjokLn90Vcu4nT5HppazAgQvsRk
yl+BeRGm9ZqHPM9KzAdtVoj2GPDvbp2HKNumo4NYW9i2tL8XdRaoAs2/3Iim
Wq/OyexEJvsFyUoJh6ANixFKD+vGHc/KiFGwrHx/g57vnAyxe1oBvSnvaiKD
Ud30wkBnsYNofptZ00hVAmQhxF8NT2V+G9Gbwi+yJNafcZCztZ3bl4rG0QXx
s5MmpNxH2xQ2URq4dFbsJzHfrirMkdUp1wzFsnv7klkYPv4xTf53CVnj6bAl
amQmKNvKGYmCSXHDDfanE9dXwmRJ6XgQedsY+mQkh/lkNZTzfEHTqqJnsMFr
Faq+eb0jYEfDy68nqMPh1a8qxyBx1YTO30un0owxidmU9QXwVlK52O+CjzP8
lu/4Tah2Trl5rznCHqq81Mlwad85z3TWw1L+1HSHuK4GQpeixpGil4pF1dRo
ofOf9xZZzwE8WJQm2Cf4iT1fgUhtAuOkfBUVUtUnmwT5eiOtiJAjT62QQUAR
Tqieooh1h4a0SdfvzJ05lj1bMxPpsR7NG31IpPs7LezXmKRTo4PgpFBeM5Bc
OFdKRCom8JyL5GpIFWBdOtFar9Zr3BlzctcU/86e8uANRKXEoq2g+s14R7Ub
mNoLCCqU6VUfjPUyqYS+jrpKsHFtgN0g66Fu701d8A921zUxplFzsFgHVCm/
qHqO3OH8gBT+N9A2etSS6rHhroviFNvzuFOkUoUPwaSb3JwTwVohfwgpigTB
rnDZbN+pgnwRxMpflX/WqV7ZL6Kq3Rpj941TtPEI/OkSaik1PX8hA9gxhm0i
s4yRfDYHuIcFRpVd2IFGdRwDvTSDx5HCNbDLutixC2eRa51gFVTGBHiCEF1C
ucFeh7UnEeazvmY6HEh1RQGFlaH3lRZjqZ/BnqiHfinb+ePllywDymQOVX87
7odCTsbKqCWNt/l/sx/eegUin+eNChnDRfRHA2F9SnsutFTFIXZUb7GflBGJ
gbUBWqE6NC/SH0cihZMDKEXZtHovXxAo0GS+gt8yLagA3mWS818m8y3StqN+
Qyzd12Y2l3tEpFkxp14VbIjMJRDZfEYQvf61/07qvFx2qHLdpIsRDq+ewQsN
88227Yv2LC/4wkAJWCK/h2tgzlv7VXyYLOv1wpxsDcgd/Y+PUxWkN05Fhk8L
qSpe1iOH4eF3P1+y0m3r3IBEtxLbjt2h3ryIuPKbHwRUuE3DANM7phHj2b61
lrPKFaAt5L5UPz+dsZKInrgX/RWzOpf2Thyuu1D3zcohVv9HljjFtjtJUi21
ZWfgEC2EBA15C/+ZKzOHtqx55wKAnfvRDBOtKDfUdOZRQPnZugqRJOKBNP3C
nPwsnPF/VVFyBWZTpSplBMsTvja4KaiM8aL9XLUPUIh4YtbvTBmkR2v60Rkm
PQwIKKtYfxpXtiy/YD3TF3LhCGfzbFJGId+A/4N1tg38WMuz/Az9GUtrJdNt
VnbCkRl3/p2L9pBovjAq7XfL5wj+tGV0EJkD+s9nTnfVPi2R0/pIMKKgWTnP
6wGpsD3iEMLmuHgt8Us9szFrsaJIQOcw/AJLaij0jTLelh3dT/7Jay4UOoPi
7jvyOBzlg6QVbvWlFFLUnCCo8lnPgzSwB+PB618R3l9DPJAYhHMnu60rjnyt
jNkH2NnCYqPJlenfzVBxWm7PWN61xBOpyIU5oc7AWAvcPKsx6yW1yrbrxQrj
sV2q8iNzC+/2pRPno7sS4J2ebu8vfFGlH0lKc827FZofRGuQiB/o3FqSs5/3
3QK/IXvo+6qsMwK8ghzq9K+37XqGehR1hc+70RhqLoPgzmART8ehtXgHIhzH
5tP9QJnrAJwcRSUmlxbLNHcOb3LC1NOtc879Ku6u87SfqnTpskGS48iXqTB6
jK/lCPPgSqTEtVsl4l2SNSLIMu9LFitsb0DNHLRmc54bDv3Q+OQ18PoORtO+
1hwtnUAdeYfhcWfr+G+ag2gSsYYza1FTMPIeW6j1Yo4YhAjdTJmGXEW8bnYD
Emh3IZwRWH6XtHpqo6SmuVg6h+aKolBfl6RaLvPjqb9sOtznoDvuhKJuHDdJ
Q00viyuc5pVMJmLNwUHVsxPB20bKgcunqjHEsjlW/R2HKDasmZ7tSwBDv++I
ZVTy9j6mlj4CaXCEOqFRbzpkLM9TmMnTJnv2Yewx0eH8NE2iDtM7Dk8qM/Bn
wF5lcvOmFv1CD4ewDdqzeia3WVmdc2KXV6shFey38lLvCqVO9TsDTCUyr66s
m5d2mAS9/5uUNchckmK6M0QK/Tqk5zMK+J2kHW0H73hwmWPPyiJPKTWHse+j
TGJdhXeIQICdlFS0BQkagnvIoQf+w8xFZyz0Xngr9gKksUdvGig/EjZ83d6T
FH7FaGjEd1K9NnbexQMiPVpCS0xYA/VmcK8cpwKHyk6wxWRGG9+t+QZvAD3f
HNNCMMpmXMPdDk65/IMcFCcCFOfcJ4jdblilvuIrXdii4f87eU6r7QVw2onE
Kc0R5qg8CgQYqd1FlSS7QF0Hh8e2QWjlL+HyTIxmRrMiPu3g4edzy03bKRp2
hkCa5+1ALGWtxnJnvEeHh1X/NWnDBiNwy95x6OKggDqzGZXBYyfWrXTqreIz
9j0jiA2mx5JVnMKduwQMtLPFkNjmOlG9dB2AENAOVjhNV85t7zy2VnoZDtBk
I0N+ThGq/VDoqYWfxrWz/PEB/DiAlsYgo27a0gznVPuflrIVXwputZdCVsPp
OebKofYVjk+M8Oeu5ZMCDQ8zjlPj7wI209Ykdxh+mWYkf0LvdHWSau7LZbE9
dxYDKM6kAVH6eL+Ooe7giFNgL1DwzWSrbJqSxGTaIwiTVEflZYlylCXHwd/U
eddu6dsq/cXotT/JBYHqKrWX7+GMBojHZw9fG2T+GPpab8Befqpo7YWwFkjd
Dy+tRf6TxhMzkYzEhhiJddLNA3DbGDis1XCIqQhgpIOokZxAO1RvH8JqDO4c
seLiibR/qZm1fHu4IW2zZ6QZOHX7d9HTGX1W0lcuqXSizj3CXB+ae1XJP4rT
NWAZiJxFk/Q/iQUj3rFFL+gtzAD0CCSzvDLbiShXozeXy/F68WvkrSU+hG4f
Ts7PZOOs40xTjC/t/wIamTgehsXHKDBf+ewek7O20EWvncHooJ/sSfv4KSg6
UxM4PRJP2o1Pg2YUNyqJp2elsJOn8vTWMHlXn316361L3x+GNER5FUAwsgX3
32BFwmmpJzl0I9Y3CACaSitYHmJdPFDjOQKUrEqX426SETqMnMI5+dnmxhUf
XBKm0uFjq0cCwXvS7fqiNM/KpgFFZbKYFdIRw+AvHFyTDJt8a805foWsecad
yMFrKwvMffOzvn6EHSAHMokMNIpaCdwldY8HL19vI+CMyBaQEuDH/l6tp1cO
KIsVHKzI7X4q4tBE3Jo08TC8fNE3+QTMSJ0V87H+CSc8e5MJQ8Bb/vc7yq9w
P98GoRig+mfho6rGGpEKdDaQ2drVMTgRUNy6qk8GliTGjdO9BbRHRY6/JGSG
dR631LmDn7noo6NtpO6B0ztcqzVWn1oGt4EguokJwJ44n51jHmm43sqspRaR
NNdw5W08QD5I90mhQtLdM48mIg93/AvKgvPLnvkLLADKxP+3EEIyf+gmyQcr
BtdAQc5E0+36n73ye9kPL1ECOI7Z3GcfT4chvYJMXGgdYs4ztUwF9d1QybEZ
4zp2pP/6AgdssVEQiO+pwHksdCIQqJKY3r7ZerKOuSFXybkUd7DhU/712N9M
AOQ6zetnPm4PsjDyl6ZQX2KjPetx8yoRSEJ3/IQeBJlRTL7xmrS+z6kezwIq
hn5zTgFXAoKGjk2nqEmHb7JlAFqIuL1JvkBwcj5XZxlj5Xz4dor1Sq+fgtdg
tDXgydlar9vyerOMoxKWXsQK8C2cP5rKZ+Mm5+ukRR2nxUKnsNmfp5WRO83b
+q4OpYG+P1+G6ER0oSitzub0Lbsh/wzbllszUq//kUhEfELNFCq0hW2F4ao7
Z4+sEsENCu80rRV8O9FzjsJHyTQCZwT527DQOpRa56Q6cZ/Ced87cL58jAo3
gZvdpl9P9O1Ygyvre21fEmu9B12zZMNrvoJ2FDhlLQQY7JvPZBIrDatUff08
LJlJEGVlLK3wuIw6lwOA9Rg4pcS3LfPu+ic4BrfU8fZYNMGHgchgx7YMMKuD
EJW40XFhxC6ZaSEYnqw6WvTbJZZKTRKUfh71XvQZBbiCsugOOHitR+fFW6tX
OlWvu0ij7cYymtJ2f00T5ZeBGIn8c2nQorYk8E3jTBlXOVNxL02QOIwss7pG
JJpN8LTxk9WqTitZhY9hRLkJQwiHV0F1yGvQzno3rSv/GhdRQDbDMZ0630Im
q8B2Wi+/oCg9LG7GgxGxCFkAAu8XNAojMhiKtX5EAuuhDmU9LyTBWBLBd245
n0CvSViGjgXW53fLoL30u42lHudoCzIHxRgk4nJBBgkjjoeeqpbIXE3yHDZm
YkY5F7DmYI0MGVG/es6z1/wWrVMsS6iTBLmWM5PcMfdbgBM/d52IXzQx2lDZ
uk6OYfVlalKs9+gSjl6xhc76OxvCa1e52Hkta97hfKQHFvzDosLpbbXbgfJc
IYzlJ3cGCjnQlHHZK5iRxRzCSdHLLb4xfV3biUMvBle5zmbth4ucWkr7epya
891BxjCAG4T5gKH+M2HvLO7KfGmPLj+EKEY0VSgQnnRlI7yeN+0vHKheEfty
aMIkGx/gcwLIIMG3gY/Q3RVOxAMJ3C0d5480H1l7ZC49AyyuKqiApG2pq5xb
sqJWGZm0yF7nQwmEe+++Jbi619dHJCo6ayjoQinFN8Rva8uvLvSuUTQkcTE4
LWKZ1AGY2CQXUKYVxWEf7Iddyx3utfCY2SJDHPJ5jTOK+IkrVasBxSoBESe+
O6hHkSSa711r/Uf4IMpTPAlNKmgpV3hEv7umfQ0qU41JVmoAysfk+D5YUsIk
ne4LOV31j3iN+jFTodsU9AGP1iCoSkraYdqLsP/BBaPOEWMqZW3VTJZbLcSK
wDj8tuhYjY9ttHK16dFMM8KZmZqSyiPT2AQHQFGZIepSmxoiFkJ2R7N9yLYR
MWezquHRhZwtqB1ikGKwT7Dq3BWlf4ZTXl8Q3RsDeXRO3bkleZ2yp9ggpo2i
JezbX773b5ZW+s/2k7rLoeafl69Y/Q7q1KWK5swif3Z0WsP9DoBFcShDwE1u
RBcpmlJNXNuN7wW9t8mt4kExSrmmOHCQ2WQE/mnUHoAS8+g6+Tc4H+JNyQ6y
ON4gULBGOtipV5t/7qo7VFPJlPvTFBWOw2rGqVtWAAiIhn1Mf+Dy4B14fbaV
hA72yiK5EwKVd3hjER/Wzuadc+JkLR+EvLNOostnJv/2xYPsR8cwp1nYoEjt
4QeG+UGqhzWDRzTl1TFekOG+IBq9l5Kbw9x16a46zhxbsXIsmFQ8Y9UF5LRU
oOF21fzbvjZjQJknOe483XF3rpFvg4wG8IYeuq8BM4szSvPYIGG5JJkk7aH0
9RKicf9s7YlFRFApqbFW1u2FXjWtQHk+o93OX5vLNDSjwRGcwbfmHYM+M9zE
+tkRoWmHB1nywfvSvpuLyMRlPUcs4lRFim89mypQRQ4IcQvgGeKfm+6opDVT
GhK9WccKSHtXuZnQaHgNQIRpZ6bpFAJUOqTM7njt0Pxqxnd+mUguA1a3U6XD
x7xUsJk4JvjLduTqzZhX1ZXiPoS/tsy45RwXyHv2EKGEMJ1aIQTFlwMHBuVc
izZS1rCUmButuW8st1oVTTwh/1i+EOq+Rgr8p7EPyfYPcIGVB4me7mO5AxdO
xTC5aFq03ZWmATE1KrzGzdZXHQ7W7xUpP6nYhuEcNVQa/uxcZOpvAoH1JKxU
bC7OAlrU4LQO601fTgTG5Ei8BOv825d6N5+6KNTK2h2J2bUGht85WenfNM3w
ZV3kZGQuldznKNW+MoggfTE7frR+SaYJaKLrfGGT6C4RYSSS8ddozaSyM5v0
tsWonmDdTiIowxi8lTAnUQOCkqVDgnQDF5dg4ZX3/ImdXXuv+LISjuG3DZTT
MpCzbYlNewbFyD8/XFO0AHKe3sT6Q6GomKkB9eNYDJdSUtkC3F6EOp4HIYhE
VdESqgtf8vGoSjm49K1H2HuuiP9QBlVYPYyI2csQOrhj6oqzxCM4KshKtqcv
SIplmMm/9TlCxvkc0zyVsV2h9YS+KKOeQdBx+KTxbP9Tx4Sn9TjdiFepcLMq
Voq3sI4E6ympgOzOb/VLxzFHegSDipXR8de0cF5+NScPGTSAefNnXrlomwjY
0ZQNyqIxqfN1Dh15YOhx+Gl0Ksi7lMedXHnjsNR15zlr1dx1ZpFFNjkr5huh
yvCI1zSwRwVuenKky9l8zIWmI8IZqNM91ACsq7svxIIQ8pEmi20krBpIksXC
naHAdKHK8RUROegivttAPFOZZz8O1fT6qzoE6d6eA1oVzcp5mW8FxdSnVZHW
BsBHdf6BmRLWNSFMxHgCvbf3b24hXkdXNyBIRWesAk1oEj7LnueV1uTYJPWc
wYgKPQ8BG5JAZhDy159lcBW+ENvC6mU/QGEvejm7UIcTWVCl91nhRd1XZoxU
BMLZQ2NXze+EOe2STRGsZRiUl5RBV6wg5dxqskbIubrI8t0ANe64zgaX4Zap
Oc0Zp3TUzdhpJS4YWnONkl/AlO+K/KAAVwFJ1dqSz+1eVmkOyZQbc0xtw0DI
FClkLdtO1vCQpaz4bnZKbn98TzLbmu3lIjHOwD/UQ/uF7p35DZQmDy/259C2
l2cgNsn/boTXoOjUhKe9hgLuqe2pqluOYJI82KkzVQ56NoU1Bmp3HgJ4TWaf
FhLCfxQcYNw2YMxOesYtTASe81/cWkdT3wKxIfs8j1CSgDJQK0+uKx2doFLG
eXCwjSWHDFasPfaQfcMuFLxBQnpOxcu879bPL8BdUpQtMAJD3yYkmeIkPfKS
ftR48uv0/x9iMv6uaCqsRUj+GtDCvqz56JdNd+rbz5WqwDqH6rCFN42Chub8
S5UJ2AqJgtuh2YvayqGz64JuJdxL1aBHHiUQg9AgnQBkfbObaPjoyxx+iMof
xF2z86xOyzgKmvKtdEFi9gOE5WWSnhT1QeyXV9v0/nWs+/oOmtxBfVvUShJI
eFfovnoab7rTBpaqlVab6ktWSwn9LAgwgf6Fv8aPHJgUo3tspPWtFcrHhYGy
0QCvEXXcCrGCORaFkYYwSoVAhAwIrhFDNlB9B+xFtBljUhmVZac9ll83+H1R
4/QrAk9LbMdxYvUdtRWEO1mdtdvxQxaJQJiAOD1nV1netxLDbNk578r7sDyX
y5VlqqKCKNMjZzq1L/U+OhW+7e3QG/L5SJNbU4LpwBAhW09wZWXTknD8sDM+
jG76enR3u/OWKYD/iOBfDeCRaI9Rt4cpcTNvnwm8OlXxbI0BBHRYjWAuKee2
/Mia9TFPegTJwAeQqq2oLfgLLXJcdrg+U6vrzlm6kjKHKpIQgeRuzE5tGE5G
JS80emzlgtO0Nj3E/I+mFaBhQ6uHD1izMM9DyXVEB6NIrOsY/zCvWT6Sbq8m
pGcq+dFS40h6vUA0A6sryiHrxGEy/n1OuYc2BpZtOdmMgFCSFitRngc5WtFN
UVhULtDdvwH4532ACiv84TCYhEcE6e8XjQKvlqACQTQ8dgeFawr9AyZX7ugh
V4zJvHU99GeeEFgS2Bk4ZI5knHaBVryaU2Nj1XESYatMGHxW94RCA1HqQjcz
+GhXobqSOURSVAEZ6jNjZb+5k9L+JvAA/T1NkyRUT59egsHpV4DlzC1dtKdh
687hSY/70g/dgVXDQ+cg9OdVPqQ5gB7zPeScq22nSbJTMzG54NmQgITMpOPb
KCLWXW+AHuBOKTYVxsVj3HcLNLXX4mchlEnAHuHF2w9ubPzEX6iOnOmMWqjK
sCH7r7+vkjm9e0F3ydgcW9FT/6q96V4tMKVhAIGFsao4pufZJI4GkOssZnBq
lrRFSLxni0KS11X/E43rFPiP5LwK3S6y8e+GBLsguBvaoBwC32a1VJszzvcd
jJCXqlWsM9bSY03BByoOzoORF8BcPJNyKHt8aZYBCkk+RpkS9vKBCtlDRie2
ODHm7+fIA9iOnYP7LnO4wUxpbwXiU0BFU8rKLA88VHbLHafc9rqZOsNlfx4s
zJ1fYbmCIc4R0mbwOS49KC1oEf745dxQ0W9j4rp5meJLz+5wMoU/z3vU30IM
5NJLctefVdYlYZmewq+O8q+UZ7EEzt7zdPgK9tjBFIV/8mm0cXi0QSbRiBgA
bFm1wDUp83A/qyExPjPmULbTQ7/raYjncQRiIYRe5JOp93UFijDzIokbb49h
SpIMHoHN8bkb4hrdPezlU44DQzV4ESh9LqBHsQhchJqiib2V0/BKx3CJPtPP
Vj/cGZ0eWvU9DM0gS70RsjYdkfpgZ4Kwhk5RAyA7HQtSiXChtul6Y8PowoLN
SXkEDoPCsqfDewPbNo3S9TC5pH3Do2QBh0r5ZMuk7GHixImTen+Qfi2PdhhN
HEEFbbTGJA91m/paIWoobXGbz99U5+q1+h2SX//IfC7d5Va8lMQQq1Yfz9Et
eRWywCUkuNfgJOkxf1wzpJUVvb7wq1sNx7gtCv8v8nuZ+IWpErb2x5cXcdqW
w38DsPBgY/zk4ChXzwm7W1nBMz+gFquPLVBNGDHy4t0unwwMDggUhsy5hsdN
YoyOznhAvIkA7IYWu0b7vIWfPbTYLBGEwRg78EQSXbYFcY99TUtp/PN6giEO
5nHxinNHFU1ofaOkjHKoFk1fYTAfQoBVwWnq5LR/eu9MHlqLoa/0rwvR1ifH
P0lxyizCBtETSxpZOE8fTDTdrzlwXtJUOxozEitCCdI+GRE2yLTX4FyPFgGo
A3/KJGOtNljAjXKI+qI+1HNJleMvYnWP247xAz7oN/4gAxWvv8zyMqzRBbrJ
sp+gBodCLoiwtuY/GTpRRE7JBLWoL+3suDEEzlQPearXeWq8vWfehfPTaVWf
Z15q8AuxBFiPKvpT11jwPpE8sAsZL/NLDgT4jO4unl3svj/rTXAT26pGQlM6
j3LnFo0TKCJ3TriABqALN7XPFhdut65wutcvB1vmyvdGcYXiRLmoAr2Yvuxl
k4TIDTmh+/an2pkse970JuplNzY7SRYveg7X0FAPs7RLIb28L2ecxeOUdUbz
tcBAXwCW4Lu29p+FOpSpfAqc+b941j/U9mjEcTLL1r8iH8dUjljOTosmITqB
FwW+DHZcb6HEtFiPyJuW3pctwnW8Cu8Y6R3GjLMCrwx7Kz4VWCDoqMmkhsmU
bPe/Z18emmwRN1aHWnv0g03lvnoIj6DL+jaF4W7mrLai2RlLdGiXL670nQl0
++cggVVKyybKMONilWD7h8qVr2sDvs6Oy4jCdgtprSNAATisCs+zW79BD/WG
Xn5o3WC8O4GXgHypOgBxUEnVF88CTEVvZPWZ0zUKBmCtWvfWXTbY25zbIb/U
JP6lhuolt9xQQ6XQR9Kv4DkXnxnZ0ec0gP/cMt2wVypnEv06s/kMpDDiELFc
nLFDWus5OQL19LRjIQ1TxlFmauIL+lJ+HK/C++pRBkCTBiA/8QwYir1GdKDN
n78HrfFYuGLopW6v+BTI5q2cQfUaZLUfN/ZhCpKb34+lMeuj3o6KKlmv9h6b
TwB+ny5hsAqUv746yCbFJbbKDsbNnxqIErc/7Z/zoErqCcfCYb2vEbhXrd/P
nO0HLTzNzlMUX330lsg5KtZMK02BLaoZJZI//7fJ0afJLADKsA4WVqbigbmh
qvMK8omhbT3ygPj/+T3DCopm8ZHPHtFKzDvDf6Y2Q2GfmNivw8MHNfi7hW8W
eY8sSL7o0PIMLFQKduSSC3gMssZevOzsGHCk2U/ZN98g7q3WhJTYvcP0FpwC
SOeBSkv3nCHnUCw/Pfq4KDoKFCw8/c554vMhtXE3ReOCFWzml+PPQS9ZxiPQ
C8Hfxhn/yM1cmB+nBhn7jMpMYV7HlzJDJPaHlIDt1h/mH8P+34p6V7t9Ltgx
rmEKElqKr2xYtDp3ix9ZrjnIZI0fIkNypI5rHyGbMj1jwDOtEOGUEMEU5D2q
96BSYaGF2FWKEUuJECVkK0+ULQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mCkktOQL8KaH25mWuPSletu6hHW1oA3dnmbj0QRoFJIOerTHM18Y8DaK3thIkS/C5xXfwbQj8f7cDUYT3BkCeGQc1qbNMGvAAMm8PJiW7Y1gzP0Yuu1z3n64lxSBO+G8EXzZKcjmYHnVhu7Kp+rjBtV8GHpW93eaaEOmTqQsOLg425m9GROv24BvBCiyGwlZKONjGUOgQTnItV5BFiYNAHsOT2YBCtVGwPYI62sVUZ4/xfB3mfvtvRhSA3EfFXiXEnWM2TFcFRvNrVscgZLb6c5sxac/cLMOuHn3chCG9OI9+gGPVfe3bunoMd9CIVDuz6l41Ym24mlNlT5zl0AlYM57Xg420XbHuvKKpTkon4j4zSMyf0a1yArMUZjF9+65rVCIGIEhzT1F2ob1hghwfS3X+7IzDWwrljRQ5JaMdTGHuMswVrRFRJQ7bZCzOCmB/L0tv8AcC0PSBd9//JRxcfe8SARXDW1f9gYfxddG1W8gBrWp9xaL6aPXGnaepx9wWCRJrQrvxGMz2zOt8tekaz91tFBRudLdujxHSV/GU7IIe7+2mW7Il5ioIwUXrVPBik579BkXZ7PuHZVLNNHBH6ic4+QHGT/OMHHHOTQ9Mw447xUNEcKg4edfWZEiNGImVx3wYXN7FdYCrCcUGtenS+W2Jk9euH0RPMpcwfmHwvGrl806xct8Z19En7kywuAmsQw4jbX02fE2HSE9ZPst8KodgRF8BsFlK/y/cCFWaJzYNEFXVPb5Ej/WmwSeUyvo8690L5a785wMUam7rGr7cH"
`endif