//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c9bkk4vgFphV5b+p7y0gK+u7ACLLxKqplwHKo4DPRsJNWTkfsay20z0Nvqbp
gnwogUsZOiwd+m8HIskysu0KBMjJtwBZNSMLFvw8HN+/hAQVIzvV1JUHjDVd
KTsgYGCpJDvaSXOwYPEKkCFCyP5zYG9yBZcqJT4luLg0w9Qfu8+4GQ/I/xiv
P8xZK+90vwEc7TKHTd/Ojw0aFXc6PY5LcqE4aUImz0DVvegw822F3Sg2nS1E
BM39Y4G3uYTNXilW3rgOj2A7uu10z5MQ6AELk6kqjTFdD8fOnURj2lpCe/RT
94yIT/qnGeDqHaLaYZN4fofe+pCZCjKnq42E7laJhQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S+HN2/I5TOjhZHr19iQKUQwCY8J6wxJKzLrdzVYiFPxLCnBUzfcN+JP9I4yC
EHAo497sRKctYgWtRm9YxYgLEX/AUP5lIbQxtIYnwK3kSv4XFHjY+MPi8vRe
gjbOKNsPOYtDsXQnc1vpd72KCnn+fRNqVCB2UDC8ueTTFIzQMrs6hKKIxF1l
PpPMtGTD5QXlq8lAsYYPQaSwI7R3/QGczRY9Cn+ar3dDr9c2yZlm8TMYrDfP
/8Jb9KeKrKSWgQMnV2hJX2ENmfQ3RpXQpU++39SBglIKl78+u2C7uI+8nl5B
bpMXERPP/GCNHwdUhqGq3GBJlGSnVBWxhigGDJ4y9Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
CE9qCUTn5dA6z/nNLEr7KmaJiiYN2ihQE2/wc+HJ3Nw208R1y2ib3SqW7SSw
MfHbMhQIwAtnKyWaFmgDpsp84/lYSaNuRlVnDyf7YQjwC9F+4Bkx9ZvA8yRD
JWR9/gKI7FSgJXALAF/nS9IiWxYo9ShKI4DoruhbXNuzauC/3u79TG99lWP7
QLAu9vkn/3izdJxec4VL4Zjv3strlpuER5D+B+MOkDWNAZygAtaQDT0ndF97
eXBD1hsls1p+8q7ne6Rh6NRWvcLoIF3HCEO5gOSR/MByGt7Cq+JIJcATe0oM
zdoblwJ6hoXtCHg4eyS6uWo5AFRoO7q3wpNX09EfoA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
R54tS7hZ3PcPJBexKz+Sqbo53Oyq6Nf0pTslKRmc6be2HWIiru0xqDFOeMV3
mYHlwGTqLNWhZbmwxCXNJ0FFJ6fg26tQF5hV5c5l7QZ6RENil0/x7kDbYLbv
kueLq1Xi78SPBjjlrKy8YwTF38Up3x2woeb+c2OcR8b9FsfkKpM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
dE3yQxIMaBoDGluE+FJntp03wviiqEzlocdvIi6u0+aEw1NWdHGW4Vi/hRcv
9V9rZXaNCdHD2LrHg36qtG154ZwDKHoV5/bavahrONvo3lzcEik7MFo8zkdm
8CNMnjx8Y73jzc0JLVjoW9cWGQX/8++65ZF+gXlsfLe/n/P6PmrRHCWy1wfI
1Wplej8Fpk+eIsC24urr6hMTu3Pw9fQewnqhiEVo4B8s/Ak2Krdl8P0vyBNd
5fglEZQSWdCCeZJ/OeIip5//73yCxEKG25HBW4rBeUs2jeijwWEs3n9+VupZ
Sqv3SaBJSkPcxa/6XnGUmzyCtf4uRC6PCFYyC+tQHNgn5T9KpVZoq6/WCpDR
9V0z1KhcnaoF4ANCjLfCgpZ3uuMRa7oDqUMoelhUva3X5UYV6A6uRUFldFqY
BFtwrwifXCmt1Y42fMqu7AlRUmJM0ORz40N1dzbZJbYGBblwbhBmeTbQpEVi
91jw+nBfHeJ9vpJhCT8KcuMlxhvgsZKo


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KxaPJ+wWJWTZwX4GWFTcZTnNWILOb6DYsjma0zjcKrK/ouskMnA20/CmLZ9j
DecVCRvuvQ9bzPIhpGRbuih26UXFw4WL86onyaEaHrFI9RV5N6IO1Kl52630
KSF+dcd40RctagtNyO1YkdFcpi+yf1DtoaTme4ULA4YFG3c3nWU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
E7hXFIZmoocuNm0VsEVnIXl3w0ledYzilkgSbt5SJf5xLHsbhiyeDE+V5CZ9
a/+ApdkVQFwqGlkfAIy0kAkIMoPkykEVl2Vb5McNsy8/l0CpuOND43o1Huxk
3ppVZgH1NdR8uCbz8wTGmGKLGLFRH5xOrPmXa2ybHGwugSw3DXI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2064)
`pragma protect data_block
eBepE2CnEwNP+vYFiu/pLU/KviXskcgL/7b5o9nExxZuFNup6bJSSpje+wxy
nlUjohoGAtlU9M1a/CnAVkMkwVKCrI6dyChT7dx3SJCAFlOQJgbYN/wv0G18
ofNfUiWJnF/NLZ1Qw+Tdf/av+qeMZEVI44ad78sWWW2bXbOxQ2H1LINcsNMf
RA0lb2One9xiqpNUAeHBdUbaBgsFVe1CstIUD+ig5Am/mSV9LWtNdZZ9HzPh
OiXNjNrOP5QV7hYIkUb8igYNf3g2dXgFE9oWJNgTl3R3ZzKpEH88R+vgKAbm
zU/HVadkbb5dFvbPG1USt2i7D3vNrxy7rAdJxSUTMnkdwCZlQcC4yhZnVBS1
UHuV/UFbc+5ZRZZdOiCGhS6z7abrCRP+l1HovAAtGZVyxzVPLAF2U9gP9sxE
4cKgiBKqP3ZGYlTPfHokjKkJUaco4Npo8zAeUsY1fpN202QVnt6Vuj6B5eM2
fraafhXc9RAEXlNqmd89eQf0Cl9sD6XDJucreZuYaREb1LjA00CcYeY6zipy
OQIPwCa2EPEYF64HH+cLfl17ozdJ3SGa/nj9eSpoFA/pBDW4NDzQgZ2HsTlX
i1CUF3SBQPEmRO6nMN/LFO9+u4vB292ssL8Hrs7HQdtX553Qwkl5q86+FyWT
Mw5/FXEdjkhZbDIGJT+qrJiH+kLR0XD9K/A0w2WE6NjtddknqnAKXBFQW1Nv
DOnbzNSB/6KZjlcXnCPDMxXZh3C0ETfxpBTyVGKaijWki7nN02Lcp4Hq41qg
tu8lr6/prcn/yB1kur722uj1DIcsOOU+1t91UEcei+OcK3JJcMIywKLx8Cl7
d3Y6FTLOgSl8K+B03/fymPbnwMwX+vUjSGZyN/fd2uDJUIxPlMOawU9eSQ7x
3z1qPVJM96KcmU+xvoAcTsfP/cYHnq+vMFMKdLQy/y6onwf5EdFmlVRVlkeK
0tjPAbAnvjHAYy/rGtHY3KpFQwVP54zBUoYgl7oPV8nPDb+0jAKewkcKKxPB
Y57B3ACcgjlkdbhDkNw3eFKGJKF/FMyi9f33883x5dVbPO9ktIdktzXb5Npq
EyvRIvJBpx+iUWR7bb4OQZ1/18MUHJh81YXIL2bYQmG2+3RZK1UfssPKQg2f
HQh3CtNyQO10CxVj/vWKodrDiWO1HkfZ0NC7lP4t6KXHZm1Jqfd6uQvEWgIj
cjZpN+DiaYqI4LocynFhjy5g4xTWPeQYZd6yFwNN8fzSRoN9AAz5zvIrOT++
YtG9t87W1vJqyGWl1KH2Hct/tO/JmXNZoi21gE813PaXh043Ddc2z4aa4R0l
Uqi5NttaykU9+LbiCRqgY++2gyaEA4pujbNdC9c6XX472iXZEsu13oMAOGjc
t18lzUmmESRct+bBqklMpyTbDUNybqnlSnaxTD9hO97YZD/fHHsSNNQRvGVb
+drOFqA1OJ3eGwQe+Squ1U7xn2JHTUzShvw2o1c7xo7yGPs8QPCYsA6DVzmt
R0QS1DMVVTDZpzKfmww5a+elSoUPIS0uDx1M9UUSQGEL6kaIkR37F6dNl+ZD
/3H880dJgZAzqPc177AJvZPWA9zOEuc3NcEVtBYdxXrB8wQ35I5uzzevhxTu
RajWCp5M5pPMGfb9YEA5ytelCwFU/OCGbg+jmra+ozceL56jAD1V9dlzVZEX
FDJcphCmcq66yCD8Qs+VwRXL80czUzIOsNSnY3ej9M/JQ3UVD2lIe6HuVgS4
y3dQ9GmO22B23VHmW/kculBfs/O4EDoo1jsz31TAPP1EE2n2Ii4fqxMFk6pI
RI9NlUrv9sVMJ7imFsU6OwB2lmTdpdXTcKQT9aZFdqtkCK8L5xckz91bFzt/
50xEY/QI+lBKBL9wjxFzPVCqnbt63ePHdbSpdXVmOeOi1Jq9sSZGb+aF6DdL
1kwZo9ODd9ahOry8OwlsO9zKbyQY5euoOxMq+N33czG90W9it1uVABOCD+/K
lHq0nVR1lkrGCFugB8/bS0ofJPEW7uCE1FjRMkI3za3MYMK8SBdqrCRLvQEa
fml+g9HWMyVhkCfE92SzzOz2k60m8dXms7FgFUwHqzkg+OLsAqHwmE7SDe2e
rWgCNuuKNRx6YvT19fLA5rAzhFQ8JW/flGtnPvWqlZ6AtIGoK15NHGujwBHr
tCy7RyGkXHQwR7SHzi2xhFQFr/vrepqo9PQVMR8gR26WKQpKVFbBK2kI4JEc
pVWL7a0Zo/oLOj0/AgnH2TFfT4onIx32tvqKklfyT1eCnCzFS/XObGLjyhhw
ak7MK3nW2lARZwjDB53T9fU4A7uwHyyyk3TfxUdraYrW0DCMzUdQs6hA5GQz
VE+uoCaeS/rslyMCb6ul90v3LBdpulDceIfdmF1ts9lUpmsRTg3oc3Z3lmu8
rm5q0iSbOjl566SpeEHihWrMhC89bs/ZE1fWR0tDhudYS3NKqwoxwP6ng9eg
UYn18BhuWJ5ra8HEzhayWDxtL50FzXsIntmdmNAMIURlKYlv2Qcf0uosNaos
0n9oA8dQtUSHt47AkZAo3R5GxDRVSdnZXKL8RXspYyd7xkZoUDhHuWfnxNsC
cPfgw8mTxEQtVgO/+vPwzHer7TZx0w9IE2MlIuB38R0XF7HY985yJzokqfLY
nONEY2dufciDJ6D7Y/drlhqq6oovzeHXvoyCsbpBFpvSurjIFxAaEAro2VlT
lAcMM1q5s3UgD+vit7hKdd1k69KmtCgBI6p5dCtYi6jbZ1huGG8J

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mP3l1ONJNNX9Kwkqnje4yeoH5UU3JPkd+PKwjNTaL1cgjZPVW3Z4qx9CGAzVrX+RPQ0SLjOmbOlA+XDpIk+zhJ5jedtPoqYe41+r5stjaIANE9qsYKPML4qtvc+2ya1BcyKHL8FODP5FuGeutBIruXvqevpBujkHLTWrwGS855e6IDsuSBocUVFQhAjZoQWrJfFBFJTYraR9EgrLXkZZE+blqzZR1+ew2n0PkIV/mEdQ7+n98ILqs+/3PfRZlo2o8ySqBeyMvSvKLFiQdFmCOabA6XZDgcMmihplZ2YBDcJsvLZM7CkmVGZuyRtqFCFZkIVq475tegwXLRMutD5kMQMevK1/u6wXuIfmHHI7fkz3Yz1gQcrBXKuZvKPD3n5EvbeP8t5cpSF6TCIP8reo9HQBPVJU4YIKkGmfFyHu/rOvhDdodTGuwHotxHwzYeOyKbtNiOtrWgQvKxDSCCDXEkEIizwnAbki579aNHKAOzSFWP0RP3R5HpykolO+dkph6hd+eeA1ZtwbAjB955lv320NXn38PJD9LDWUB4cw3/yKGIxDru6ZbGNZV2o2B8ccSgErFGPTuHVRzr0hepDzVWV4iBkEsxpzcV5oGg1KbzERVfrT8t1UTyyiSkoFsz3Uxz4CzokTBladJRVe2VtNqgncPXycVnwqCDzBCfu3e83SGAbL9hH5WC5WW0OfIe+j59wp7opX5SFoqT2HAnsvdAnIocn/VRvlvjpDAk3CQKJSFr0pB4kDXMDDeGUEKYMmRLt8xCp+ACD1QMOwljiqAJ"
`endif