// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JWWwSVtr9oTarFRJ2Q5YH46zIQh2Y5Po8RGoF/dT7iv+pdbsPvkZfzLXcJ/k
maycBNRUdGuQxhzsmH+woXgy0KnBbavP838m1XyDylmcKDHEYXX1MzkzF5Th
5hDoxdGDg0o3p37gkEiVUkvZ6mL61L8yQyTvKgvEiV7lPtq33BVmk91q2px2
h5ztqoLUPcJoS7hcZq4SQAf0uIGSkvtGldeTVNgKtY/SFIcjubBxhBOtarMI
K2eGXi3wWFXQ0xAvIafeCkcAMXa/1V4LGJqYL72pBdtqnY/mDLlFPSeH06jy
ZWOjKsttZ1JnTU5dijvy5i25lImyc1s+LPNDAdV4MA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Crr1ZwQespz7yG+pRfGFME6W3K/S1xhG0sPNqrbhkwkIRaLj0JOxVCxTYr6x
eZhIvW+cdRBxAkDlDb/ENsYLDwOb3ZwmATkkGZ3B67mDVProi6SfdSoTliLw
XdaJus2z5wgTVAYcG55ILBrvqeow/W4ZsIhgv/jc/eH3pme4y5FhsmeqL+cr
QdH0aEqSzO+Y2aBYQTCeHMElWf2uf1lK3++kvaGRQ7jkhhEB725VztwFqSaL
cS96rrl8pBuYSiLdRzmfS6MkNAsUh/YigyGN/KW8XqOLD0X/M2cmqFLHLr4B
FgfCEYuCDtbTZHbYF6AfyrP7uvUQh1upfc7LMkJUgg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ZZMnH//vIPKhjMh40wkfPAfkQtfx4hu7o3ay456/Bgcev+/7G4gMlvp4U6Sp
v7QkcxuEEj6ktogMs+CzYIxfM8y7iCGQwg2nMznsg9jEThBV9e/GvRfwBKPV
spMscp3fmAhHeSPsUBhMmBs7okCrvi9EYrviholuerc+fHYnF9BfFCdiv1f1
8Yjzv6nL6d9apt3rLZLHICiUxpFP1m8Rkf0vPy1227CtcM7Go2iGGYtoeT/2
NMqO6WD+yr67AFF4FaqmHEUZ9BPbDOw8rRN8/shznjukI7f5sxXgNO7iUP3u
IrucPIH+I62VZ9sxUfHsB11rp13zyzsHHTjyC02/sw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VJIc6zA+9LeJuAo85/cyH5i99LucNTgrOxGdVyAH/Y8M0JZVnClP5qikXRFe
J4wf4a5Bho0U2H356OaxBODgfecjDHms7z2gV+oL9taAsL/bEQdeoeBcsTV9
PfkyOUdBnR+an+PcEmZPkyGVmFPnb4pUVT8xXp+vfnMK8qkeq5g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UlXIArwxN+aVkKvOUnYMcZodGvqe2vgp2byySsBGjUGE4WemXex8Ub6QdAna
pIV3sxwtGnfB1WT70nQHVgcXRnOGvGmb5am8zsdGRnb5awSiGU7YdggiKe3/
49mAc+PfJO3fAEWALLfgwtmTm2edy7snQn0RTZBoPxvO7grYCWjIeFVFTFXq
Jfcyh45Y6tULmCCnP2adnZVoBuQyegSb//egfrAzfJS/HtzSN0KO3wUxMObU
dBQQjFTJhJoUmx1I2kSk6Rvf09C2cN/mF4IFottfx3cYJe1qpxaeDHao10s/
khf6LCUkfszE4NjtfoJlT9hkJYkp295rNJsYJQJRiDB3DVusrKberdjyvJIh
L+Rt0M3GhOoBoBVlBdv+kedzdBs8Zu0UDv9q+Z65gJPXc6OW9WfZDyAH/4xc
gVomwdegLQuU3kCtM+y1wTZmjnnCbBQ4volEZgIxYEJctV4rKJ2GyD/avlcq
PIBRPN9FiMUpy82EQqY174X9Cx7WhqbJ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lX4c9zzxBctOrJyXD6ILU6B9bbbDaDZlY7GsLvEGAwVfgHQ/+1Pv3Ntlsqfa
YxiHrq0k8i+oGGqjtykhu1vom7mgd22TyS7iI4Y0bZJGwODUxEaGcGcldQBx
EfbWr73fTdYRKxmDvECtgUx2F+01RQP6vDYxm7rnaFpyo6T+xtM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
h2Ocsd4AAaW9G5W3zmHqj+zjhO2IpNzGt8bc7GI977RvPPM0t9XJa/A4l8es
R4q19E0Csj3SG4Uhp7pcQgglrdzIfT8dGK9l60MSaSi4TcRMV+SATcXa1+gd
02sF/WUeoP5D9wr5YQEPYNVFmjoGtWeD77FeKjCNa/U5rXHoZVc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 10288)
`pragma protect data_block
n1LIXb8ZfoebDMNixb5I7jTj82xGtw98kYly99mGSRWy5tfWRFGX3Bx9Dktr
mcka8/C3G4/jIQgBgqVdd+723rBF408x7Lzg/TJeVQpS5dR2+OYeblZkM7hJ
xc2h/i2n2jQ2Y0Lpqa/n1TQgyYGryw20dj7M6Unh9MF6qxUmacj6WFPM4XPk
C4pgjjB9Pclm2OmhUPBRle6Dmos1ALd9XuWroUTP8d8Vb9zwcYkmjXuzOJBN
aJeKlr9fXL6Vk5T9+C4WaefYBCaqYyah/a/viuhGPw8WtoGVke9sKA/2OOUS
Dz24Y56+cZ+TkvAFXdI+2NkKM1h3mITaYbhNpLb0Q7GsVyVwpEnm17L3K8Ld
EGmJE0cgNliIce/sQq+1Rjlv55oc7pYI7YSUdQJgY6qYBJnNa9o/sV4q4nlO
Zb9+VIogHK+bU5e39IxpnteKWuyAT+hWhR8HoArOIAutAh7i/js9Q/1T6JG6
i/HhDRUAlnKnfr8KCAKCzBux4AXqGp9WDw9EvXr7N+opWO5WO6td5Ez8svyN
/ck9tqNzviA3ivVRTumDBZYFlVCWEGV7TxCuzPnQ/7HLoemlOIn2Yf6sprt5
2Lay/rAFxEHpAmbDWmBeEs39lzj21dq3Y4HR4mh8fS5jH9KFRnMBEYFta7Qi
V8FgqSJsHL1ogob0ODES1Xo1ly8x54rE4bF7yTY3STjTQ2DL5PC6MzJxqnJr
vLwzBzKz3w2h99/Jlz65F9WteulDz3nOC0bHarsROm8hIlEzQXZ0EdXn2/Un
5kM0GXOX4ptkEVzdUSHVDhvHHUcjnW8UIg1rI4SI9AwaFSJuwOX8xOvbsmMg
M6fl9HBtJXejIEjWQGDSGPB5jFE4rgFfHaaB/fon1cDWYabrpDsMo+qFErfo
LUxN/BNtlJS4IA4SrQNhm7m/UjHsn49PEWscG10UaXuQBfJTMad1Pmvfyi8G
iI2C0i3Nkj4rQDuL+zBXgBVdAs8IZfnouYzClVHqx7KpglIkBJ+BbMmsim1S
ls6Iv8xNqT5DA8nQppK3/LmQ4n8kYHUkaI4waC/6Jf6FNsIbQwVtucaGny/K
+ubIuNP0hAEf2hfyDJdVe2RHC/c+hXcd6PS0niY4a97Ay7PWVvHID+lb3g4z
t+pQPv5ooSQWQjZgguQEHe+Nu1f3hzuPOG0bYcwKNuF04EfXNpRyXgZ0eVVu
AHhhLNqm0HQy1Xol/DRcJXswyJf4Aj2SdpxwdXL/+XWQE//X46EB4dbkBY5A
cCB0Vdm+0mZFm+sjGZHPEi5gWBoWxQcR++D/42Rl2jHit/b3l7QslrU65kky
ZBSeO/lJhPZCWDYsP4lWMrOewvu2PdNcPbw23S7RFSWTkgui0NY6BYfOFJDy
t/UmS08Sf6id2t3BiFRzqP5Mf901edpjurIOye557F1Eeu4DZE8BWzMAmLJQ
r6SyGFb7InK5fTI7Ia7qFPFHq+b6WvH07N60mlEzJzp6OJ4J87Gp1GHtKH1h
OkoWuchEe33LvEEDwgd/36UcJvi3ot8p1bHgV3HsicKRRESF5nrK+uZeXQnw
z6rx36rUjN42tR2B5DJRy7Rxy+zZOXb1h/USHpEdTQ10VNWJYC09X1ZtrgCb
LFJNL+BPDXlnFU9Dq4sSqaWToIY2v1aVLSsD23ZPCyQPgNVH2GNcvi1OU1pP
KjkGgGk62pkZ3Uf0heGr7t0ui1i/q7zhyhmnD+a+f8Fh8MI+bGnJf1JGpe20
5Tudjmr3/7QGg1N02TXnzkqpnQQmUx3RDzV3Q+AQpmpHFJ90txZg/oh+QoM1
ZHd6PfLip+qsSn39Ar7ujrKMDeE9UBZ7NZL+8eEKmwWO94kOYrpwYHU2nd2s
+PKAU2STWUg4ZlXPUE3UdMUbbTEcVTDNXqSuv1JdgkZGhI9xbqby85038iBz
kqVfF7pEK3AUsVe25aOYwqUTkecsZ+Z6bxHcZYYRI/QHg5GSI9p5Pjgfhdid
6OwPj993jdztswO7uuk7oQOZJGhBVI0hjHxCJNbbUq37zz2T/eHpmqW8B1hs
yiuJ4ZrhUq/Sin3vROdufw0ZHZW9KdDNQ5+oPX7Zrz5l5Ea3EEKKBS9EyYIa
/8yFEpw1zH/8xLopH9jPteWML0BubrfU1bJ2ArseeMZ70zYTH/kE683P8C4v
TTljP4MBnd6t9SJMZJasJaxmCleERL0luo4K/o0Gb85lWuoknXXH/UpQPsd7
Emg4uox10CBydHvFrUUF6JpDYY1xErgllmC4wAm5V7TqQA5z1RajRbaKJI85
PuG3MHx+u3TK8sd1tD2bwoCBv63oT1wXhzy+kAs5zgjfF6R80Gia2ZHr7LzX
YKtlT7B5UdYPaYukWx/eBU6/5frhRJalRebYP0Zm7GFCyBiaaI9MlhQD+X8l
Pjw6o+/FutZ6fo5UK7s1Sw2GJ0GsKOO59umIwI3AZjLyPR4gWUdN/DmzOeqC
lShqmAKC44iIXALqOXs4MW4ZEDDNYLCci2P/x/F+9KrkSetBAFB0GqYmTQ8e
MocDsASm6hrBU0OplJyPMUQQYdQMfg1VSUGq9cs8K1WXeAHlWYylTuIleeXw
Hz1+76OXxWzBKgyX57tm4LkBNYuW4qPEI0aZZii+6fQMVX2KZloXQO8MbzS6
RyTyND+RHHczw359njr+jdOckfiPfr3GcwhGH2adRpjfcsUdehyCvvrV7TVX
D9l/RtMX44jf4Mqd+HWF5oQyWpei3RN/TG7yod6l6GgYQZhcjIq/FldxIdcQ
5XEg9KGPmytaI+0lrx3GIM833Fo+08HRq7n2p4vgMEG1wAALrKDd43P5PNoB
mojqUZW4c+5VqvI1PB2gasxAiSdqJz9cWDJjndLtLyNiPug8QZiLJ+JNlHNn
qIL2tF5aJAyyqN8c3WSMtLKzFbjNA5Qc8Uy/7F8HlOND2W5HvI4sWhFyPfwE
XfR2ZV7Czy1zTsomOENVLprDl08IycQY4ofwEb+25oZ1vhOq5S7NeTa3woLt
2fo6qX7SaGEIjvDGPVthwFIjIO6LqipuekgGNblQV7gbsd2bFT91zxxoSX4v
JmL0be/WIZizW1yfH/Tu9ih9p/hHLLeXv0sfR/NjUhTGDoHuHoflmBTPShGA
Mga7ejo50375Ezj9R1E3O78H4i5Q6uFubpesORVEeaJOZ6XoDm4xFz2DyBfz
06kHUme0Yorat9OrbWsSinrAef6smhC23cxvc5XcBfGAyNM6noxFGRJtJE3d
IDXFcgYwMFpdhtQ5jTHzDgNqOGULcISilbgYWwLyOqYIxqUVKgsFKKt+yNfv
9j9r6LYdr7TfrnV7G3oE5rszzhNgO0AonrB7hr+S7BI/s9U4+sSf+Rojfpn0
LfEHBvxFjPyOWef6EN7RK45Up6Tg+nQ20zFW72naPTJ8nO12iAWANAWRtEXT
/YmTMKZq9p6wtAlDgx+apb4OvtKbJQ22DJMR3KHBbJ/+EhOInGw821zq6wQ3
qLsYRymTmH+qbjVTVbM36P2IjMILJsTEWGYelGTPaW4EWkF2zpzBPT2cuaYw
IQzRCo8hYJL0f5Ti46ixWoRNs/G62V+g0ZC/ffTGN5cgZ+I/tygZ7D6tyAun
HcOiXoP3pFMHqxuzTPSkmY2djiwYFtTzIRnBBG76Jvz6shP4bWXH909RS7L9
LYm54igwCzpx6agn1MJG3XkK/BLFNUmmGUvJ0Ab+zCq1m8Izw4iqQLBZRA6C
t+ij+hVjO0dSgEacsNDGFSkqXuRm3texyZdHK0ajp1R12jRNWDL2q3q7XBXt
6KgQLWsmfh8ruIUiMWhdC/ti8s86nN2VBZlqwoZfkSgQs8/SS3yoggzI7PDu
RyF+C2lVuhRhY1Z5cHL4MaKDbWsvBg+7EoZprtCWMJWEXmMf7xiKoQLqCotO
sEJPpb4mAOKsKPJnOGgKFInIvZ9HpbnFLqiQkBqLf/OnFINOIHTfCveTevd1
KQVaUaLeF4vNf2q39xqR2n0/x1fJNN3JEDOQuLPNCbjGEDnGiD9nDmBbKxHN
dTD4En/t/dpvLd1R1BNDyaL7BmCheIDzmPiV6P9805q0+LvpuRSZy6YVQ7d9
Hefv9YOQzB3Ijma5HxG+SbWPNozhdVEtg2GpxYm1oHmyXSayYx5emeZAhnTr
BjpwfYAcgu2d7SlICQBT2ukE0iVWZN0OglgAptfpIEpcPFapQ/OWFgg75faU
0yHFHIy3Z2H7uSUQdxpUPFVwtYtZUI5Vum2Lg4W7TOf15qm02OG+GFDvLCRE
WDcajgWy+qjJGcMnXzZ+Be2zdAHVj2Ragz2hnwCtV8Qg5t18XL0ZK8HoH4W4
S0eZ6W/9caK+rJAPsDJpFoaYW45FVKI0t+HMuUiZLaYr9/+PZU0pnv5Wz3aB
tBDr0Sjph5abK2X4TBfGCy7XGczhV+N10GMj9B6VCB8PHU3iROwZQUTN2w4i
RoOTGzu9l8PQV2P4tkgy/pHe0AwukqPFjKMlZH6Oeokyxnihq+BNQtaO4e1N
csRVllbC4LHjxe4Y4gB7woMSQtNKXKO0TbZ/96daIA6C+o+EBttHT3w0rOkN
vrltuGtcQjn9Dynmc0iQ7ardWDFse6BTc9z6Ue76rP29DTixHTsddVllzcd8
OJ3HKbDACUZdm3Bd5inhZr+6TmM5WPBwTCqJgzPVcbDxIjaOfC4EoHJBeoZ8
0WX6DJjZC3aB6DTvsQXCQ0Rcsp5hjP6p66nBExwA/ocdA8SmiVYekwrK5mS9
4k/0hNalvr9YY/iBCHIzK7/urk0+CenXGnWfAKTkqG44/jLmDEd7yxavuiSa
2lVvnZXOIRszElVaR0vKzczN+QPkTWOL+GWBPLJRqv6cmVCX7KL0ftyjSmdx
wbq+VFqyInr2/8H9ademPAVY+gLFI8lzFBVCHIpbjYaBWP73RodU77ebTLyZ
ZHLg53iNA0OP8i66TWgV2OlkPxL0AnJk4CBlL8ThCMe62wMpetX11x5gO8RD
TpIUC4ybxEquJ0l+vkG9Vws4UiVFyl0TI8m7baPktfV2UWxBBKtYrRR2tC1h
dgNwREzP0bkSvtsPtx32s2CKZjCnGvW3FbX+yOfMAMy7blKsxEftPRg0+Ve1
pKbDPGjZgMB4Du5yJ+mDvMzg8r/tglWm60C/OD317sesZmu0zTPprv8JE0m1
GtsoMRr8d2sOD8Z/Szs45TEha0u99MCevdDDrV6bOhhvR5g1alv4aLXqoBx2
Afr1KddNuaD3hajjbPu4GydwWRMziiDEJOTJGqT2xittoZt4Khx8wrCk9uaU
C5Wb4lj2JopJCEHHKLwpLRIwmo2vFLOfCA0nKt1liyGZDTiwzF3v11JOyW4Z
deGbM4L5ZmIacXP4zZT38De4cphUpGUFz4xhtun/e3omExzsUwCeesvPTGz1
c0UeJVnEJJvQoc7llXYOVcJUR5h2G7cPbRXc3zxazRs0Q7TmreCSLxdqWcXB
GziqMgipOHrSXQB132jnwDXDpuFIJXGROlY8ynDi8nNtIoU3jc0hdpfY9GZ7
ulJqdvjjHggpwqsePsf4kf9/X5ATk+CP7GgCRATOaA0o2QhpwM4f2oaugAYZ
wmJS5iEVosodhB5IwoOLVgmmhAJBraw0MH9UhjwOmm2Wybr1Wczh5Tsvwd2n
6mFNUWG5xaKDblxrsqaZ2jVm3SZPDyL/dOn1ukDn/+N+M9L4gkNtWrSFjqZj
G2BBaMfk+M4eFtK7Hi//WJ+j5comzAU+7auzaNobCeyBWQUOivu2hDS6ObmW
vpZmfEHXEqB/4JX0NM+ZOH4x+vX3w1pGVsfzNFNjpwfYZWtY0WK9FP9mkCjX
pSN9fo5DuqRLqfuaSsOPllX/uvdN7fnN4CyFq3Ru0fZmgY0MflcPBc5gu1Gx
UG5iteSGwheBo6anBXxm7RPLHZHbvAITb+YLRhgxcflBFdJxEWu3/LKNfJPP
t+DpkvaW9FGJKghxD5kgSQpgwpZ+OEjzf7oU3LY6+BwPZFueEejKKqOus03k
EdYKrLInjjDmf6mZQItSW+Q+9FaZ3xtwzYOCLPGqgYIamCyA5Il2xKZuTs4a
WJG4MHhdMp20H1pv0PoCqI7u6G4TGILIlo1wrmaSpnGZ0lakIpwAxMhQ9e07
0ABoLJzY6G8q2CAKbZemucCJ9/tRQHCzFofIEr044I76Io4aD/DfEyt9bk9T
yI+5GiQ8zMCCz6NIoNLYdTn6ixiqNfiwl+ARoaZupvCqiDlbIUj6jahH11XQ
ABE9X5jsHc5cX9Ic7kIwWAqbid+dSKUe1510GnsugBGBMIEq5VwCDhuvhDpM
QxiOwWidF3HQIDAfxqPdawzo9+7nquqh1ONwRAwc8Yw6gQxJZSZNwbw8tsId
DluCwNx5Z9RKjpV2KeUHdwyRC2lWr0fWFd46WLIqgl/U4xHYfhuMq5ZJNde5
PmX35qRjxTrcvjzsbvHDU25uvEcR0xiwdofLI7CrYzqGO+EMq0bId1bfatla
36W0DixKGNXbGMn1TdzWdnKuGa+xJ5vsp/dNpQt8foT3v/g7FGtpZVmi8qJr
sKL+CHBMoOX1D2+zYBRNvPQHGmMsgqvLWGANZLFKDbSEdCTLwywkanT20TgW
zfs7O+a993LZFlI/XGHrZE/jiCgBOxrM45BUK47etF42oMNHVsoSOo8Gk+ln
zcJRx0VSqApkimFEaQQvN3ksqInT9zikrq+Wf3Hs75PJO3Tqcs2BtEYcVPQt
bXu1eVm78flIkZ0CVh7bxkEe89XO/Eb0V6hSxiOYre8AbxeSsUl6Zb4kd0l1
bY77All7Zf2MtISwlg1bZ6el/n/FANO2FMTryhsEOzUc8k91v8IU0CVzchI3
6x7nVKBOlManu40ilczUCwLGgjs+NpoP79mFDRKNdanmtn6ZZY54bqGAc6j0
e8wfuPTjhvef+2IF3fSfCIzM8fJ1dCEFkwqOpPPcNHO2vN2ZG5XEK/lCkPR5
vvvdymsEtb4vPO8HVuHQkQBZMmR1j6OVyni04/Z8Qv9NNIta8mJ6IjioszcV
yzXtQnwCoOq1ZYb62WbgYhQfqcg3Bh4Jq8ab2l9RRWv6Z3zYMN6z8SApZwIK
eSnjwJYQEGxEoVUyD10UbNuDGLYIXwfbpYR1buBFon3kekJuuDUG2kbBAzl2
+5KsLMDcFzpsLmhIeK7FKUbpOIlnyWYTj0bYOA1PTt6GV43ky7CkIUMdhJY9
pSyP+lrJGpRIwxdpLLkkCDdB10vyXcLbS6QEsC4FL7fu8YUXm/WKX2ANw7Iy
kg3uoWWPQvyIcRPIf2349ub0ck4K0AdAMjQupsj6f1g1ojoAME6Sx9TNylBI
YVWtN3wWQV99wOsP756Clvzv8OR99efUl07QS0dk9XGplG59JTy+bDxAhVcK
YcMMnW8B6J/pp2Uv/CfJ4E0j2uFNXZ9T5+pqycdr90AAGGFOprQOQDh/Eo+X
8olRjXd/ZTl7cTv4cMfFxC/WIw1CCkPnwB7Fl9HcytcCn7iOFkpQJPxa4IwO
KdKpN25VL0XNnx5PeCQoxhjnZJOMAF+qxni2nPiaQ2Zxnu/c6Z4HDFfQ9ZrH
7LjljHBFradPqTeLegzz5KfWdJcj0tpRMMl4Ma5iBlAZOEGfNHCVM2IMVGGW
h8rjI520/AbBXsNYlDI6z+ljfYa8VOBHQafnZ0/otC/rJF2U3XQc7idR+ap8
/5JdDy9nGRpy25F2qVwbE7/ABDzqvuDx+szrBMcmVLB5ttO0IOJQskYLmvsL
uygW1pjeYi1rZ2JPPPCbBCN/qa2kCYgvIgCqU0D2D12Zj3luE1gWjw1sUHpY
RK6vmv2OEmz4iFov7epm4LYGFMxT0QsOxS/QfEJEqo0Gg3cIIxtnWqA3nM5W
oH1RYFRhffjn3Y15gPy7Rl/apjRXJf8k77KDL0GRBb/rdVK+tD3Z/IIzVTv7
JCpRn0WV93oR7WRoKuEjEHlRFoAe80I653RvfVBobO/bF6LoVkeF1l6DgVfW
CHZXHjEiloCkSKbrb46Cx0aVVAp8FjKImBBiEtRqDYdZsRdbW4NmJEAgeA3w
fG1pnni7w7MCb6rxj77rUXTiBboaD1h04FPbQZCndpbrZf7pY8buFhfblc1t
l/KkotRQZ33DPCfzXNVzJ7PHXiBI8hJEOjfXa1yj2KTJaI2mwUN3XpA11uWE
LEgE9VzPaNq75F94iK4pzetAyeeHtwlKdjdVfh3czEIKpqpB/a5J9frrYSEW
OxgGd7SWZjEgQenpGK3eTWB4W1EyaJCLdqeAphjVGl77ZKLEpHssRh1fEZok
g37xBcAWvsS1UeYVomBjOuRe2Si3xQNqH7U3EvWID1IPS/4oaoRjU8QvUEt1
Rko6+L4PK7NiJjqBSgkml87EdC/Ai1WNvidrBgaelSYsTKMQNb2TkCsawZ1g
i2MMaRDT8RFv51YYzYSsivHl+cjnHQLBS1ld+DU1b/0IpqoSlEcoSAiglnbH
u2OfEa5mL67Z0jWJNd8I2Vlj/D9Y9BeN3bB4y2knuaDGY8fv35BGF+Og4p9Y
WZV03Fh4JiFa7q8TdxJN6i96Gp/sGuHJF32Cc9GKbG0t9l4ccKSh7LHz/Lv6
0Yf3+W3onyQ42JaxxaByr3wVYiL+b4XUDKNd0gbC3YUID6pL0z45VaHt58jf
eW1gXoHkNznKqZgi3xTKzwSBh0Ot4wMhG0M2LMHIRfrdOzI1/pss5fzbNW/I
pvIOfWSEM1nOGQPvjfLL9yEaktvQHOITDCQwua52fDKeKEEpOieOvsoUJOOA
BYs4r9oe7jkHlpunhYRaNwFmqEXEOwMS+vGaYfVnlN+Uk3NS4UAX5EHnJEnD
pNVOmQFR5dH5PZOmqWH6ZewYOQwtJ5rAaejDb4KZ/8TPAwUoHFixS95+MmGZ
C+IvSp4aFTFe2Lyw6hYZj5Q3vS69xVYJ5h8V6PdQpbRVa6U0SiW8w7iK3IW9
QzZja9LPMxA7Zj9E8Y+nUqXhZ+pISYsIOqD328jJqSx9NSLi5D5Eicz+Ql85
zvc/mYBTwk1+Lz7six5fWNKNpU9DgXqkKlmzV4EQZKOpkxoHDoNAOMdLwrlK
TJAYTdQxfA5k/wUJ/63B/H8rceEpE655wtSmxfLJlUwyaMLo/Q39pe1Vb3b1
Z5RKsg51UvopuKBdJDGQN0RLqCg0Kn5Ju+iHTqOIDoL1kmEjkJWTImaMrQBe
PpMxWt+h7yuRej6NvlJxGXe9DwqhTn3QH7O0HsUnVcGSUfYrUfeZXw6KytKn
mU5uwiwqJy3FEzY2masdXuVI+28nZ+2PhdhBXZ4hjv05IPbrk6S5/zoiwv2l
x5PZ0SpTGM7AOjRwFlkOViR98c8tSZhwziZgdQ/fIFvj7u2xdoXxRmc+DXgp
OOBxh0khMrHxdjpcriwXpN4cK5s3LDOc+l7IX0pFTJEmWaOF2z0LzytF5ysc
xtiiDpo41Xkca+zas0AMktpgLK3Roj3QT2wmn4jRFV6HNNXJI3tYkmzgdT9z
ZKbXNMPx/7xSLAN4z3BLOeGmesa0bMzK2HmCqk+dZtgwz3BEv4Jx8uvS3acS
wrHKRrslaUbtgDYweiFAtdQjXy3h8G83s0a6702T1tPEVnfV+EAaWmOwPkrF
Sk8DY3UXAIWxjZiw+UaUJLr4qyXDiXAgXgCR6MTAjEluV+6PO3XQejJSZgIM
baqz8MObONha7TdSBqt0WWIJKKZ6qLxVy5bD63irmciB0BgRGPnDspwJpHp5
zlvmC6emVpRXRL9Q4eVr8clj2GXU4YKhJigafevExUgENxhWq1VNYEl7Q7Ul
LZiWBv74DeF5dKXs8yWUirmxBVyu9hBlB3tah93XBnHFdeUNOScdhnXa1Bpv
S0KD+r34+7cOrQVxuai7hPd50S6cX4QUcx8/YQrfK3cY6wlfTg3sSyjAqs98
aTfRItGNvcT0DLQL9rVnZumWt4XT7CEBFkjIEVrwLMbvCQ81VHlHrFamtiIM
m+CgKPuHMaSyCx+7R4VLEHXZpHZong+klI3IRfDOfTFk3szeOGHkD+iwA/0m
KMBdX/J7Yqbun/bmTm68OJVUOIZmZYILB5HvfCvu9wNgDBtV5fqftcypvzgJ
KKjlST2IO7nF5NTsh4Z09UP/QIaSzI6VlnaIkIaB2b9rwpDS00Tpjkhm/fnu
pwju5Ng3k860DoeqGofWELhjGqjB5fPBH/o7hr+KXUa7HOiABohhnBYiN1wC
ZNOLp0AJjeukBleU4NUrwQKT2W2hlAjZGrrTOk8haI7268pQTV3E0N0SsIEb
xsirklHhsANqDQLYORFpMhcPXO1Ydrcw36jcRP5aStpYIjWIVaIBYeEhg/w4
Pmk1XJW+VrF8Bzz0QA6cYAv7GBm8NhfgydV8f1cJe2cYXRJvDw0sjR7OfKVH
6rUvH4Os8R9WyTjthmRZwkF6szcZvyCHPDux3/NXTXudWyC3nz6Bx3OZkxvR
7CEQzzaqux6K2RDd2PSw9zjtLL2f0Aeo8ReaVEimBAFQTXa9ohgk7MO7BScR
JfW5Uw8jQbUsV/jpO/lIHWmMHaKjXYdOTqQusjLSz1JpDzsV3PL+SmeSO8Ue
cxtiXzjdjj5qepNyKV/klHhkzHdITBzN6lm6D7cY3wVSHG6pECAFwRolpXkM
WNLk2icvURk+zAhYgiIojDG14WdrmH5suqUTAZls9OTshsrInC24ubgYWL+8
eRFKmexqwni2jCAzQ/p3kNM+YVzp4tBOR8VS/u94WwSMfP+TTIOTwFLEXbF9
/OISLstRuCz0dlOaQQUXzw4BJy0/H6xmLFjRkRk0F6CUogDgMFG+05sM0Rje
83mkAcI7iqND5A+jjEEMEv8LP1WdnvrzvfOF2FdxR4Vmm9FtbIXxVe1AdmEJ
tqWrNlEVEotDc+m64TpxQe5WLV+/KI3dE707pHhRiEOyglnt/3t5bUXpNwoa
6v/XLrRG8+cQ7FT5NijUTIul08SQSYMwvqWjPiU0nhh2lCm8HYYGqmc+C7ww
CdqH7EGrpWTO9QSoZk9sKpcH6VQdpG3crYzYFe2qGbvjrrXjwlYtzdjmOPQM
m5ky8x/tSRqiV/BE8StQBL6eXhzU2Qi2ia9OuYeIynOV7UvsrN3DzhB2tTzL
3Y1lbMAPCMcUYlQkinTCIpnXXvyR8RfAAlXyT0SFeTShn4v6gGxbPfTvmLlq
JHGdtQV/S05Gh3zdNB8PCnpvKaAuvMbz5qxW1IG3G3BpzdzC38CeWA+ylpD1
chIqrYpsxElQ5XH1nqdWYEndgq0EG0yDNlW2r2Ea3PzuZ5p14+1N3QIRnUMR
pn5PrqEVAAiro4a9lmkJuYIr+0XX4JmbuYq2pKPbWAf3kdTXJ4/CxGUvet4E
MraSl50U3chi6xrwno7wubuw6aa425SyISGcmHiHsOBqZkqc6TCWFq3qo339
1vH4JSWc1HdtSndFTNUAVeRl2pv84N9QGoLmTnZbmVqk99+tqDpWAXkL/uFI
1DWgZMBrz8YAwkYnmXNoPPhDevHnCsFXmNi0uBN8FwvY4BWlQH2uzsRjfVRl
9Pu6da/Qkg1arJUxPUPOM4tm/p0HsmeweeeJGvZxqWVW55S0Diz9wkczV59h
Tc73Wk8QzSHPp+zUEjTDiKHIR8zCQyPn7upcuH4MQdQ//DVH5zhsrttaMQU4
19dDNvXQ82j6PxLHsKn94NCXzWARIVqu+Haj0TGth7YB1xF7towMaD3fFvbP
Ej3HZuo8I/k1K46zNCuhwnuj4wfUfAB+Nd4gHa73mi5Wp4KsR4F7mbbJ/fSc
Fk5mU0C7/5X8ls4NmVNdJMQNQlMTZXKtmjVeyRkAIs4mX31l0gpTUDdZKyRc
xqI24hD8xzwkX8NoDYFZmuI0Va0h2cu3ZZquAHCa0rifCeSv4PI5wht5BtDn
+A3nLswavT0WyQl5VU4AMVLhNtPuRJlWG5JtZAWqCJyeL1/syhNV0qM1yV7k
uEMUVu1OCXA4wANUPAzi3CAA6F4WEA0Odwt/Y89clu4icnGU8JK5e5F3Ee0O
lx5BytZkBTlU6DdhgfC/me+Ku8btbDOrzo6qFGfSj+CH7NBgFmgRTuRssPLf
1INDL9Con22DHK7rQt4VEPNVnkCFp0Y1CGHlI6ypyqoCyfHj+txf3wDSXJ1X
jY6v5lx6SR7VP+UbZbI3liNt5svAWJfGTJzW3i4Uqq9TcK7AtVHK4VoC2Ctw
c3jgJ7w+cJXLhqs2RMEec4cvSWyN5JtIqgrNImDREeJlTUZex+QvtMd1yPqf
Uyf/j8RHVcv6mgUNz8J3lRPvDcSEyvrCIA41iDA9GLbjBf3BveLHXAq1lZKy
4BLwPwfTQ29i3brdtCVGBpv7IR04sUcGpUvo8Zk/MvcuwTdDWWovzoJbY4dY
zg9MF19/dCjm8oT3NQua4Z+2TsnNos++P9Nx8qabLbnHH9uJbgvcbxtsKQ2n
Hunp8//dZRXV171U/eGxkupHJxqCGE3xLFhcJVKlU1BnNbytnMm104r/54pi
X9nTZaXGBbShoGsAqp3ZGnHdNNncIqEalCxJa1gBhkYaCzhLgIrzuj5j3dh2
10yS6uJHsNXhndnkztoYi2vbAiCMqLq44mgjx/kykHrxWuph/vI3G8ilUjqK
ATxvIY89NiUatEcrpxB1jUrRiO8DHm4WmUICOsSnQEZ9d36wEhpuzMIhO02W
5q38HV+jqLM9f0wvML20pyr53K3HKXxvkGyf5vCLgukmbu74FQSfhcsRGVga
cvp0scm6qJzEdXxQBvqOn++2D04NNr1bWMbTbHqtmqUe9hg3hHoamy7UuLnv
rGtN9SpcNMaLSQPi0iQ1zkQTWAtVhjkVDI1kTBh583O5c7mIvGqqpivQx3Zx
fxYgtsmlCqaRPh1ELfCbqLJzS6jS7Gql7cu2LF2YnzAzD7SZI89MdYDWPz1T
cGlGcC6VhpFUZKXerjx87X8edI9WsoeOm2dM03DMvx4pVy0gD5xPFr5zY2PK
bOr1GLZkZgPA3Xm3YEi6dUV3TiHEsjPViHXpomh1cpu51dGX0zi2cVfIW7AH
r0PeOr5SIF0NivZlFCdfkDI5Vd/ANW26QS/jAfa1KwXxa5spQMd+z08bdGo7
JIH9E8EN+H9/sGrjrxXWqQMABGv0hakpE3rURzVI9TlMpA3SNPrAVvJ+H5vE
P6LHxUgVUMXifPhhXc4n2QMW7cn6sR7uq2IDvPlfRxr7SuVYASSZSXwHh3cX
giNF2Yf2ICPW8AwvOuCE5Gs8gh8z4vhcIkaSG97V4sKdBkFrnI7jPxI3D87x
1UFcoxPgE+eF0erZ4N4fvi1FsoKt/HHy4RJPjuHivqvKuOcLxPjYts7lsjYN
P8btWCpUv9yZCCtyp1pwO9EzbCEFUr97NOMpDULhInrhoZws55MzU0p02UH4
YXY4cRZ56HKhSeiwtsXtnwfhFqwwYMdAF/rqpXytZfyQP4ZaPd9qujNDdDeS
Jnrf6ZfqykHOW00SBYJOAPUKO3K6SBdX52RzZ/e8iXc+RiPDVU3g7/E/iBmm
bNdHrUhxACs4h3+lIVWPEVWmcFdd3QGnTtsWTWHKYX/5XRfmgGajN9UCnWav
U3sCTJL5TBq+jcWHRJJ/ASsZvtxGZKOOsfav8+ZPjkLiluwvGGAsB1vXCIsl
D/WSdbMCW0u3hMtsck3RLhP6LK9WUV2+OfuGr8LozjI/Dod3VbGnCWPaxQQJ
DlUSk2ppFEtNaMuTwcQqiPB9IQei7dsmhwtqWw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfRwPvq5q5I4excIMzUJYlPsFaaJP9I8DOLWeGQSexbSH5dj86qKFhWYvlwa/ewFzTnuNt6nVCHBCAaeRdBxOUG4C9lvPIrX6M2CPjgndRKvhyNNU66QHiMW8m+pNOUQ3skRp8Gqa6OqYTmI65CPQ3BpFDTAQQnmXy99hbrg2rGBfoPj4BsTK+nk74qIXuYJevAFsMd0SvELt+7Zd5g7T9cy39rFy2l8neIToG1evnxMzYAoQgRaPJBR7mOLf5hlJ95a8RxzTKpUQ+jzjW1C0SCdh22HXOvbgQsac4+DYMWpxwGyGZjo9MUSz4iPv1OTSUciltwVWtiWLHc5kv/IQlDCM1jV4pU+6vEDCyEmdH9AAYs9uzrqA7wgWr6pSWrSweSkY6vKy7N+eRX0wX5DSTvE2V5N3+PJ0ZUvbJ+kylWoOTwIOqUahF0uiFHKqvnC8hkYnKe1KPo1qUqm3/R8cgmL5PdbSrXGzoxYt3U05/6+pro2cTiHCOUMvLJNUiUh/leauFCNRL/CYggZ6AqFzJzQ1uR0VKORb7oYPukz/QljOWSXDmjI+uYjiJKKOGHzrscxjpo/ZOZlgUrKMKTvKGO8odY5GymqG/2qbrYu4vlgfIKwTosYLUq4WEDcvSarJ242rqJcvjeMOcFknN/fqytd7GwUbzbTxUcNdVCswMASmMV1lqZLHZh2L5PMasfdd9FdIWaPaXRGlqgZwRhkP6VOqfAZmrnixrRTtXBoTYnSKx9RKLmb+FuBJ4j4IbCizhOt9tnav8luB0LFQv0UuJuh"
`endif