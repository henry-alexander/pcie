// system_iopll_0.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_iopll_0 (
		input  wire  refclk,   //  refclk.clk
		output wire  locked,   //  locked.export
		input  wire  rst,      //   reset.reset
		output wire  outclk_0, // outclk0.clk
		output wire  outclk_1  // outclk1.clk
	);

	system_iopll_0_altera_iopll_1931_naboooq iopll_0 (
		.refclk   (refclk),   //   input,  width = 1,  refclk.clk
		.locked   (locked),   //  output,  width = 1,  locked.export
		.rst      (rst),      //   input,  width = 1,   reset.reset
		.outclk_0 (outclk_0), //  output,  width = 1, outclk0.clk
		.outclk_1 (outclk_1)  //  output,  width = 1, outclk1.clk
	);

endmodule
