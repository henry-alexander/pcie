// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
z74ElOORx1uDcIo/4p6tnqhhXxYGLK8TrjfB3i4mzWHRPVLoee7zcEVsvtmZ
BfJz8HBIQy88Dyi5A92hIoVwEUgWPeCv+LbQLI6RTqomkhnyfHH3cWUTJ0W/
4GXkpQ47nC8QCMkgFzcgS/eqPdIRt/+vxeEAAhLdHf5P2nR3juWdC4eHWDTZ
ISFz2f1KlNGj+Yif5gcsEE+3y9wrB+OvaYqugDfOU3U2a/XTceued1aUH8dx
PdYmotTxQtdDM6Be6LcXAynsA0zySqIRmNuqsvXhd5bfVsrHl9flONtVdl1w
4k/5qTPnKl0T4yt+s2B01HCcxW/DJiNFYhdjIwa8iA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hFR/W6Mbuvu+hvDvLIpzh7wVbCUY0dGiowASHYGM+EHGR8lMGeb6F8g4ZiiF
8j4BFznl3LZ8IYQ34O+m/WpznFtI/XSjSb1h0SEVXFkP4iF8Cf08cmJa0h76
mHiznMoqVK/mzeKId1vyDXJq+5PKW/H0b2PGr8wsI8iOF5y9SRau5vr+xLPw
WniBLC6NBQRXAHz4PPKNpP1612jtum5oIREwfgosrnw+EAOT16S0PHvrjETP
pgtC3W5foiDNO2AEO1D9DaJmSQTDtXsgRALbJWaJ6iPZ2pjr4XGIWsLkGbKe
ZZgK+N6JQRBoO4KJgWKBXISCE6nosEAVO6Pk+ZfZhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D3ZTeIB3Qej6o/nqqF7MirReAGcHGNMRYlTXlWKJY/ZsZeTxD9AkWdhpO7xJ
K/WNWkgGclQLIws/fMBKhLeTkH3vU7PGQLAfff7/TE4u75LuOMEylUSgJNst
0iN2Qz2MjdypvHEG/6BEYZohrhFpA0ifmtV8W7HKitB4QfB/p3/eHDv2htG3
BdRGVqWhBP0HeXZB5ekvZ3AUTlD0F6wU8RiAGDRrd//9s6mAr7aBmJcvy37l
lkNShpdRZOv4oOpM/jTwPu5vW5W1LiL2PrpJJdfZXycX4HBFlt9Hd98J+akD
4XBMvcZIYjcZjDscBgZvAyto1A6hJBHLjjDJuSKRlw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
d1HUgOMeHbjOqdDO/R+0vXDLolSfOmkK2nf4QPXBFWDTBUZw25OvPnEPY649
Tf/1CnjEmXofyw98MX0v02y2LD2vJ1x/alrGY0fCS3cUFBAxf0pr67F035ZA
aK6ZAnLJ6MDLHvib4NMikhM2+YZcBJiExTOX0dtw4arVk+Fm4H8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eQOhUpBRnqZB5Qu6OZwWXcEhPzSebFPAdYPMG6iUB6rZMSsYvWwibFegSzW8
9PTwl5Rkp0m70aE279c6nvbKDIYWm11ima/iJWCMr4m/ZHYlClYWtAvgLcyW
F5nR8HI8EM5Z9TrTQ9K5360w/dV/tZ6K0i6b9axo6tgbyy7C/7bkE3VLt8Oj
stLqiyGsi410LGCYuYgmSvDC2xjEWjPrmS2hqr4LulVZRWDM5ChVAftX8LI+
ykcl6maie+fmnOd9wzaQYvAPZohKAo6AePKq0HzJ0IUYvArf4VzRadnimxuC
SVDsdahf3I2viiiegTUV9+fwZuo9mKEICzFe92ud2gloCQLy2JcVlYdIV0Md
8+cwQRIMnUt2Q6qy940x/8kCVQRIqbA6aWtd7jGg9iVehg8HmY/QgxrCk2Ss
gBAsNJvFSJuE+Rd0tyTqSeYse9OSlw5uAna/+JPCTAc9JjJF2XI+U3gdAIDU
h17CkxG/mQqmUPNjYEcwX8Kh3EFVtIjy


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IQIJbdgDnI4zs7ENuZGn0Cp30GsHvDmvc/etmJU8ah5meE+k+H8VNAIdFdod
ssLT19ZdaXXBPAsbbnvVrFI91obWKkI35VwtxXusLkO/ApK8fHDJcvWFP4XG
IblFAxneH1mDYgTkgISzXUkiR7howkA1KtxkjtJWOrCq8Ns1dBI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ps39m2Jqq/tOfA6oSNG6nvu/PrlIc7hpYZBSiytECo6Ex/DCI0lYK0ESs+df
sNwP8tPtNSHkx0XJXxlyONNz/EM6dmqdYENeH+ioplcwwJ7pTZhfhMLSq1Fu
l95PVV9n/XnY6WowhyHubTXstQdlu1KxIL043zk7GHoqNVo7tPQ=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 17456)
`pragma protect data_block
2MExausNi+MEqjWD9cyIi3+QeVxRKifXl3yx9Dfs4gm94ryVhxq28L5jZX4P
4PmXp4OH38igqRfdjfFxNsOVLM9Ioki6ejhrx89i7nV5LIutAdBJUlWfAz7X
GX0Xw5gYgQ87W6PIo2B2oaVS8GaW+mgTPPD4sc9Mzebeq5dOZ7/WM/uexuTO
ttSTd3bQjGDx7nmE5iCSZciwbJpofZmYhI4uzmxl7jlDjhjXC9O57izyPstM
4KxhA5M6Rlc4tBVHEQMCn51+sPkSiOFESHrp8gFAVoALZMy0vyXo/mJUizxQ
f9lWuyhSearGyyPANfVd/bfAcJPzuBv4PkSIfBh6RQQ1F6jhlFJ0Z7Z3r0nq
JYs96oJkPC1sK+1iBxHvlk33LsXp/GQ6zjLHOQXKvXwxf/RMTHkyfqY409BF
F2HckcIIFFn3jaCUbsRIz+oq2cZYWBfYxZ3sgC5CTKpiA1Ut5Zd4aoUmSDN0
Jd8wuxrvncBT6DMkeNb60zxLaRDo5gvXYffsOubl5oeMzsDaAZ4DLVnRtEkQ
P8QbMsbh0VbhsoLy89GREw8BYvKofbUOhnInwAtwnyYtqq8sNsf6meGxT7vG
Z6ozm3XNxEoQiuCpUktvuQJCjNdyIKQSgTOIcxKEm/ckeddFHdn8LyzqQ3O4
53KZqcXg6PesHx4YHdVvAejBGSYP+K0BvQ/QntvcOofbm2EiJz+LhVjjo2xz
Rda+g3Jq0wPX06gnhoo26w0M2h+K1QYABRfMioGm/qOdiRT+jVWsPel975h3
fofhYau7cMtHpQ1Gy1fxST2KOk31UzdGD89pzwEMLJ5+CbRNeTOxaev+z8vD
F83W1uLfY/Hb1GH3CyF4OgZMVXp/ZavQ9NZfh2Z1vL41fnQmRky/V7Ur+wKq
UOOf7sxsKYEWH5YIQW6bLcOXJ98egex1i4g3toxdMiV9pYCUuMDPUjougIlU
fw3qEBdXjoNmn+JLPFJxAAbLfW/8LmiSe4RQME2PcL23sejaQUl8p8w8ThsW
dDu6+yhsrn+2jYIn5RYAorFOV5+rWwkcJ8E6OYg2DJW9TEDqm5nl6SAU02mK
3mSwPGyFnWYp/TIp//4BDKJMy5Dh53jjePCgoh4+DNM+Zl7NLcpi50Egdq5P
zFOTxjQjHLX7Fa7Z89sJXRkB24QdAuVWCcgKLcgCt+Wg4pML1BW4J4FsTHYm
x7tL0WCyVCuhoEQuCjrpLuyrb2qmsKQlaoGcrfJZx+HcUGv9Dwbj/ZQ8Rnwd
zzauQeQ55oEu90mzgDTdzMvN2Rukhz+wzUAAAc4DTdlttXpULyisLX2mYjWc
90O44hj1DZsB3PePGAm88EhFuKsCA0iTJqqAXgFqkOxG/zKwOBSWrktXLH48
89Sr8ZHbxBNqyvUSlMkOKRgtSCNJ+5OEq03Nq38HWRdr/97phYh1xu2PLZEE
ffsYVIrHRVRvsIkWtILO03x8x6W+hjxvqYRJpSZ3LcjnYpJ3w/0XjpYIYR9E
GBnPVSBo5xFP76DzAIbRpuOnu2llcdCZJ0ek3S7JlaJ1Pxo7NJ/y5a03mZo6
Kqgm/yvWOGWYdUt8gmz1xYZt7Vfu0w+GhzOH3TT2xVhRQF0VQk0ALtE1S7ub
MFeQscRKizUsUBXZPMRyBkcZVRgyTlznG0SahrNlqkCmHGtxOWm7i0O+E8KO
QMPvoHn1wfaE70/mcXLL5IH8T0zTNzkFYYJsyA6hr5I4kAO0Wr/hsGlSbd7t
Pp2O6rhlUH1ekL7zUWzt/XZpl4NXdIKKDgyT0vZFIcKouKympd1p3qekMqNp
ZCBIGu3qaimW/4FF/Qe3JHtze4VtwCT9zUmIUmP4Uhw80791F+gcwgsIbOxE
Kti9PnK6TiWhljarMQ3vRZdyF/lP8SYfwSm0RdjvOsfbQ3XdG/p2qMNvZ05I
s93A5Xo6nZ2fprvnr6r9FTkk8nsFh4MNtljjOLCQnNR+Q+64rFpdoISCFv3+
lkzDfS3D2bdL2TSiw+YKTt0xYCc3fdY4Fkp7Lcb4RMmHQisQgXhMuWLzSl1X
uzTvWbn2J3B4rjvnLVzS3NGmM3ipPZ7olFCfswimsY4aL2vNKvx5uC6dqL9d
c3UIymBFATDRSSfz0Ym8gFuCYhsM8Di76lI2u/zqwBq6adxZdPOUg6/fuH1m
IrV7rlv/2Wghnekq8aAKP1VwxVzT2/quWlxRkxYbk97yQa+C4F+bO98wLapW
QOXDtJ1vLoAB9ib8NwMzw4NRrAQtAOEXGNIOUSQtklRsxsH6MV8uRZCDIchQ
Tof8dTyW87JuMCI+GGUDgsZYgVPMx6Liq5AxUO8Okpo7mQJx52LTTWd/sGlY
3lDdE198YibIHmEPjDvEEqged1C+o3XUJ0qQKe2kGvKcaKvMvtYfP2Halffn
gHvFuqQVZEBkqyDGcCfB4ZJzF1vlguKt7nFz5QXb/2A2f+G4thdxQnFO49v/
XJPPBDCP96tV4cgRcdRHMpkG1sYFGKsyGBJAX8ubU2hoSV3tRo1GFSrac1Ig
wlOawANYqMeYjg4efaSJq+u4KzNAg3ksyYQv3IWRQKh0LkD35K2QGMGYA2nI
n6GWoiNwNM09D1x2bz9QtYKSc5QNeALfhvPlNNvkZdVrz6tcoGtavOoNJQfO
N65333IVkwivA32MLxy7951boVnyAMSr8uLrjmMaAxIleGTQWNmlY8DD4EWH
VYlhkIqqJEDFhIK7/oBlnsUfWoehI8zj/54gdRg/cg5HFdt6Ck7t6knRk5JO
cEFGOxHSa+DMkmCAxBgld6newVbPWuPoekFz1XS/mqnLwpDV9r6tP7aQxN93
X1Yu90/8fwP/8RACxK3ecH47ZXPL+FSppZpAKQDI9fQA9Xurqfl884QrBlhk
70B30cadDhLW1LwAMIF3MlVv7GDTJkN3tInSvUHeZI/cd/kkQIjRVr/PMOYb
fC+l+yjdcHpGmfzTSGiKON/pjKPgCytryBcqKOGeSc3+Xnll0sFic6vBYR+4
ZS4rNkYKq+egAloANPKyThxvLYY3XqqGf90AR1bslxkAH7aP9Bc7ERFpwBCf
G4WIMWHvLx+lhD6z4PLPyqlLX88PBSEAu5lPsO/csfmP4Nv/76tUyRcbedcp
IULpcWOUMzpZoi8uT1AjfdD/vmR9/GFOAb4eBiP8JRU0nTIZE6Xk3dTpS+TN
W0AvccaHWzYeTS2t3ik28GOTBTMZq8Asf5aHAlvaYz1UhTp3cMenY+C1hBsT
MzRh/VCVL/7fhs2DzUDRcELDDy99146mL0p4Ma/Hly4euZx7uB1c2CRDUZ3w
GrHiQ9iM6AwZ3+k8q8iwVop8oHpl8Sk0VAG0DIRSK9/dwvDNqbcuddLssJCb
+9ZPAsQG2C1B2ILeipf5baXexGclgQsbUpQ0zGacD2tH0vqYIrohmv3aYFyg
AcK9XvNvwjz38AKEaNS0Ajf1e6XQAiaWefLqERDzJg1aa6WmL+jqxhZdIMMT
bsVIXwtOgha8AAhB8S+fnz2/+BENKVK/ocbv548DcOLt+YHduv1A6+Nr+luS
NqMnjtXMRH7Ns0fY8suRosgPq6+6MW212eL3xh75O/J3GDi/8wHIarozuIbu
+lsMR7LS7AF8usnrPY/9ENouY20ZJskHP2a+K5SKSJDNvVugdqfMHZ7MVOj+
aWE+GQsD4zhndmRSoU+pYSMSENHvAX76gQwy7UAOYT9yELDn7i66MkIY6xe3
5t36O2NrJS5ltOTMy4QCyG+RRstaVbBhQh6hRn2tJdGQTgtsd+R8ZBK5SjJp
16w5KweO5Ho4735JLpnqIv4ykbA+baLcntV+x0MHxzHaHaB31gzDCe1PjTzM
Wr7V5Ez3ViE/aVGIw3/eASLB8UxXSji6f0poVqnuQjI/PLvRkfiGU5On6AuK
RA7Ldp3MNeWv1/YoD4kq12lB0vhxBzmzJ4QM4g1/c+hzz/NW3S4x9JWXSQve
6kDjt1QByCPg3y3KiFA1wGpj/6jvgtP8SCT1vnY5NPkf0st7z24uLn0UHliw
4b+VrYn5OIMN/yjPwWTx4O9UbTxFtjlVoEL4ezglH+u5qRa0vg5Aai18Mh8r
yEPGG4tq8L9kPBmYjudl8NfWlFT4iJTJUFUJC/khrE/a6zvu1XQlUw7Aa1iw
Wgn+Kh9lPnKjD3WJiC3UhAqXY+7UQBM6hxczJnkdniNjuy2A693jqBRom0vT
iYO+KTko4CHL2GCvDeTUQddobp02uewOjUGtusPP6jR9nQEENJrqFHb6FHIo
v+ivYzSfmpvGG/IWsinnLGXGoZodYBlnL7H2SDiYUts+XMLMwVnJamez0E+v
1KFUw8oiMfkRPzXNCE+mrpG+GvlPXEhRY3GicbaVlwFOSb6o6JzhtrP2+8aQ
mYelv7TQzr/ZhipIGaCws9eoSrJ3pVJoArDtVzTNZb6fvhNIblkPfgTMKPbB
rsvSEyb2C1AJmzm8NF9H9/Ahq4rHneSUUIt5kzYt/P0TJvvgAe3F/FOHCZ+e
1gQfHUbdx43iXWTqN/N5cloICOLVHo/RzA0fkAziLjW+rKh48+cgI5Hc0wv0
lyf3q+WNrE84nZ2YgrvJ35rTCsZlVIT2+WqsQSjDlHcFkk12rIH6Vgq1C5YN
XgyzxBq9UolCO1BtwJNzTObQCzD9AIjhg3Vgg3hbQb/5nNasqhKu8Jri7aLY
7OAbU+QBG++87zQqPBVpgd0PBacjg9+MiDWpUWOdAdLaAkK24Nm8Riw0wD+D
tKKWGTZk4CLMe52E1WO+YJjeb/LkF2ZgoD0xG/a7ECKGplK+aRO61TzIWbRJ
ZaZPL8yqpMg3fdHNwrpRGmiV7QqNrZ9SUbbfJLGzSlXeqqsDhW/aQlMVA9C4
ULtqg+DROKrwKl/hKRdSIblnU3ikqHPxtLlHCFwmobrryrZ9S9iquDv7452o
i1XLp13XE5kPp4D9oKmE97MvUofGNWN+sXJfabuHCJ6Zmblrasn3hDQXjOKw
o1LZCnQ3xDUU9kArN+SKiKMQudbcg4vUfNbKxe7uDggm57iVfZ/R0iA/+8Gn
AggIMRa1M1g+SoteSO0K4n8Sitn1NQy/+jXxGMmXgb5/lD4RWZajzx278sa3
7dBacUNcIRJ4bX9NBhKeSW1nBTaZ+CAQMh9hxYx6lt4JE5hwzfvmbN1TnfxH
Z+S2aOLWWvNjVearcqxE4MpSaPNhv7o8rRiA7+ajmeFqPiuTHxXIiB4/5az7
tbYQSiae3bIzyLCh6EGYXHQD5cVDz5mFAxqj53/+9ygQ6Xhb8VV3/0M0MNGC
m+IYYPC0ruueQunAy5g6B4hNbwsf02HiucMfkrYqj8Mz1SrN9seoHQvkfThW
JzHR9O+h/PXcKw7Ect+X5X0Bud2rYBwUmch7ya96J8sm1cpjJD2lX4BVE2D3
Aph9ISoL5nGFB9RP1SitcqUjrKSaszQFC1x03cRJ8kPtZWwiEKvK+/9pUoYz
J7CvCHJ6fNic3dqFwASDui70NDpejD3GTc9BAtQMXVNd0M+eu4g9bWG6BmCB
0fZ/eiTX0Zm/dwWBhrn5meZTUp7Sc+NG8lwBtGxa65ezssoCEx2t2kuBBYcw
Bk1CSyciSiB1WENNwYYVmXsWXWfH3UBQjacGi5UANnmQuO/4L5xRYEzE7gLg
vxf2ypnIM6nUf7iL3AwfpLVO+isx8jK/HmGDXPHM/tH2r4glhHRfaeSEw1sI
out0GSFrm6DrT6hZFdrO9/kDvw9xVOjONdjNLu7Po4TMRB/ElGt8CwTWe2Ho
hfVnfujeqYUZemj08aPhaVgzRfZGr8mZz+/A3pwYkCS9qBcmdActU+Ohe+e9
GqWGA9YmbhqGP4Unqm4/POhXTPu1h6d7vz/o4BO8JK4o2W/18A7DGzjxh4Bb
ld5VXVwU5Yyp00k6GfXs7QTWwGa5m1fJTG7LDPj0wQaXA8wyq2XFMYem8B1+
gytX2wWWUx7iis9FfEXNoAlJL6ku3wirZ8y/kN+sb0oWiCXtPY7mnjRIwQ2d
WJAkU0xkcj9wrTDCY0P0MsDMAMTpNxFxsNQaueWE7be7bgoQlpPOvnz7jaAo
bnvMrh34lD/Ezwjw1/R+4zSooqZNAty484ePV3+VlhNi8MJO/0mw6tRVvnAV
JeJRDy4sW0otybAWGd4hVqYAfFs2Qa1xPCTtvOOgnrpScEPW+JxLW/zAUm6U
B5NGANSGYoUac5hITV7217+IYnZZFnXRFYbAE6pGAb7UqYhmyoe0aq/tdQON
GVMFciFgkNt2dpH0tg//JJfVVoTCcIO+0DRKdBB306BN50Z0LqGHEQoXhAQg
8RqgPfINqgA4MhUgNl+871wdd+hJIJD4TAtv0eh/Ps/UiplvHEF4oi+Tsn4y
sKN+l/elCDkKx3EQUEKU59zIEE0u6XIvfEbEzvaaXwJxUwT5H7S/yYL9RFAT
LM4lFt3VB29biixn8Gvznj3p15tQBnYvW6iPMUZifaYoRsz4O32WEWiR/YNL
0fXVPhKkRP+eFb1s1wmoPUHyik+BKStw4qmHNjru6jjZ66yz++QKqKpvJPt2
9Bug7E69/blODPNDiccLHTgHyg1RwzxNd2hkfoNGgc8cvBjBqLuomzhAMt2t
z9OzsRXtVfw/xs39kFBSqi39WlbGQicaVojHspJz9fgH69fwuK8WH9iMSjPN
DD166Onm46S8F1FQvEd9gqWx8I8EqPq9Qqy6wHEzv2MfvXKOBqrere+LJ4If
EpV7DFjGRy0YjNE0Bjr+C2HoUCxv/Q0saRrEtLIaQMBSafZFKAxDjgyyUTBL
LgpOjnPpOdFQOBoA/N8xjDbJ31MtsTnFYKKju7hIdvIyvzC3/5kCLlyAbcDx
ty0aEQ/lyweeOB7BtEaiftNdQVIyDkpgf7BPnwfGsPu80aR8sVe0n1F1dqKQ
UcjXaCMj8rMHN9pNxTroTm9uTT5ziEAG8jBEHRZM7Bcnb6C4ZULtqSuZ5LgW
QqFmx6E+K/DRJv7zrzNtPni7w1d8l00i/t5LkiOvQEaGTnr7TnIBhL5c0DDS
ZPr6dN/d/elQf4Ci+fPTGyFIA2q192R9lhD5JsK/O91HtwanfxhWv7INN/t0
sjURP3LEsZbxe0/Rn5qoTce/s0IBUmdge2ABKMhk6+K11RokMuQVyBkXZrmE
eQpp8SU0JgAgTv7B9PudhJGJu8woA/icCPBaqDbF/vFqfKx7P6aJtjINvi/Q
mXmKfyeAMcdXgIqngaQODZj1U9+2AKgOg5oeJ98Tkluenl9FIbVylpLt8XkK
5xD7mlGOaX3HxZOALHRcSfGlvCLkoSVjjT5Iftv4nH1yW77rcHhW7eu9we3b
+t8+yvroQutP0JvIOy59xIzyPiVjI09nLHameY4U2vFMgYyRdVCNKN6sRMSc
iTc6a8KlUxKu9ZdZNbCwLqOETlpxAeIhVxpiMCD8G//0OZ2Ijg7qQeDKodVQ
uM1Yb4tV9XX20GrnjfZHS4BtAFdKn7CvFla9oLyRx4iU2nu04uYfSCRLzJW2
n6Dj6+KzX6DzaatKy6v7Mt3fg/VBFKE2dwYf38xVh3yJtL6kDbaSvj+lF+3r
dZNl1Ecw232XmaIyHDrQvpGUjBvM/yYakRLHg3hMPTxcqxosih/J68CobxGs
m5SIBsPRXJHFTPnMc5Y5q03oe6TCxHFmwpA0DkhT0TlIdkz+RXEqSg2AOVVZ
UsYumq0ltu+m6bY56YnZBbJt2sCpzaKsAFGl9nNEhKrRrPfYteDusNV25AdQ
qqz8W7ikyAPlC+Qypszj6Rbwcs7Q8f2qzRNy/AH1JTQC5pQjJfOyHcZdhnJw
Kc/PNKNYJw/aBSrUgmF+FWozZRj8tXEMBG2ov+vbFO3UDTjNzFxOn76RRyOg
GvIPFtlVqdAmoeNnLRKiMxuGuSIK3zEHvLjQnmGNcEQMrpmhz8jiwdKXXY2T
Kx/1z4RII0PEFBeS2cv845WGlrIncwd1S07TIYUscUAJVbga45kaIjLhNrKf
lesj8F9cKaMfHiYvw9xwl6ozuVWjhiM+drkjroJ1ac513ry3AhLDHHVebAak
34bZM6x/zlV1LrQUpm4JN9sr17IQ29hFjU4nRUurCxeWQUhl9s1QN1RoWx/A
pxnndZwXZx6Ml2IxQplLfKOQrtDZBlCClY2k3pthHg943M64KFZIybPYCN03
STHqAB3lWZn6U2CF9jvZgLy7CYH8N/7jAXPfFVynOMOHlOHUaWUhwLE/wnCU
j9qdCKdZNeR12wk+9IPHCZpMYM+f6SwAi5lmtdIR6SCl2MSN3oBlsIi2PyOq
y4BlNJ7wjMtC0PKtkUyUpRc2wcM0xg+25Dp2SLHisF8sTGxrUJSmewRUuQZl
0bY6Zlad8F9avAKOJsEbFGMT0OXXlgIOVfuWrPTCVJu51xvtfzYs5cP39HAQ
olZG4hEwDB193Puvn3XtWxS9l6IMcbPTV5XseA3/5Dvf04UXDPYgC7umwCye
2CJZum4VZjeVZM9kDXfq3GAsSJrcAf8Zx1Fv4atgTw40AR0XPKAwHibxkf+u
sxLIZ/5gOp0ipFN9y0zhATumjDgUagUYYKpvKXhragV5uuyhJi5d8EyY8DuY
HJXMdJj0LvE3cZSFfVGNl+knpz5ebB1X90j34Zg3Xb982Vi/knf573bfTJez
SCUo37zWofyWzppCEQkz7oSEsLxAwUVe2tGll4hmk/97uiWgnSO9CS8EsZJ1
f+3T28MMEuu9IEiFx3PRiNPnxC1pEhh1kJTgCILT6bdcBhBFY3oN3XAHTfD1
r+aXREGH5SF+mV0+8jOgTrWd7j3o2Ql8z0sDacarh1dMCEM/Gh2edBBBdzhD
gUQVyI6cl+EoXc8NBYB2s7mahRs56giMlBR36Z2Pj4UM4cBYh2gbRCkh/53b
btAil8R/5yuC6GE9Jz2T/OUWJ+880qp1ktmQjwljizfFHqDDN8tB5Ms6A8QV
PE4f5U/dta2okUOpSgK3xRi08JCb/UbwTJnt9Gr/YCScL0Rh1gO55e75/qmq
PduR+R9bB9vVHWN1nElvtu7xUWpXQSM/ptP6qWGxdhS+7UsTolkAK354y+Mv
AckOTa7Hsb3qKqQz00sSJdVJ4YXx0mkoX4cgKKoN6bPubmfoDCwJJG/dHpoc
UlCD/s1s4k+r4sLSDhzNWs4LjorBYE58Dz9geou7/p7PM2qA2pXXnSs8x+Ft
EyV0sl9n6FbueBiJRaexijfRvc+Mp1FIvsfmqsYjoZD2yvC7p1wkW8STGVLj
QJg6yDRsEINM7r8QIozCjwwDbQKfsw0pYg3I8f0edrhQzm2X/4S6A1z4EVQh
oAYWmiWDpJlZFKfDbwNa9sYpj+aoytE0AEtxQFSGjR6D7877fTHjIzQNUKZp
5doPDrpZ4plM9+R1KtkRCB6pG8cGAajkC3m9sdRvcWTEIBPiaJeYN4rxqDrh
ivqPtHUXYKIOrsJPD9O5ifzJ0ldFsizMNmApzty62NdGoZNRcfJ/jueBz9pZ
1QcthgZeeav6cQdKDvaTXFEql65EZVjt0jD9U/93KfwRJSw+hNEq9VkWJr3i
nPh0bgnlyc3uROkPZ5YKIFv98anZhaetR//tPpef7IaOzn1r74+SQ3EBOmUO
ZabvNeL4LtysYiSO+tsh/rX3GOLPzGATv5s8/pvbq2I4sdZWNgozXO/9G7Ai
ffNe1un6QLWHwaB4sttVNz6i52V2oSpKZkSqyZgvqrtJyOa5EzJWICaunuVV
mdwrVSrd72Ylc5JrXn5LYDgkYG4F8mqPcXVPZ5QNizJ9gcmnLoYZKnxKOrUq
YdJxD6knOzqI/2/jgdHtgiZgg06GbSrJcyCU0pb89/wK38+H3hgVFmkE7CP2
LFw7O+RorYLAS87OrZFN4aVGkdJIgI5plml2NMMdAD043GoouaixhN4X3mQd
QTEOsUBcidwIwN5rn817N2WasVZyRAyqfTEcI+c47of75vVTpZ2Vb3mF2NVx
z0lEZR4uEpEoEpLwEwIQ6nEANjptDQJEWslE2UoQ384myIMHP9S4EsXebSRK
x0rhb9KIkGqEAIWtPOHI2acp3O7iyEsca59Wia4nNjVjIvgK8Vg3fmdi5Ec5
IEOgaiCPQghYrSE5KkvaDUU4fp51mo5XEYgZfazhuHGMobuv980sMdtwpG0u
5f4LdzM3bGzp+0bUVuw9QLyn408cbIsZZWRHhKP+q4nKGZYA8pPcSGxYMzkn
ryeUMy8tD+X99JL7xSa4pyOJOv+qmrKSlMYJQwC3EDWkHx8S6ZXpMea44051
UjDD+Yc1WEiy9WGqNepL/be1oWekot+bBEhIfmiUnn82dTISOP52HPhfPvDu
HGS7gKuysQ75p1nH2nzyTUtJSybPIuRrEjNNCc0OqUbM+85aVRwE5UfJn0FB
NK9QcKE5UeUbOfgjxnNQaie/mO4bA462mfjF49klkm04O80FihpyLK6pfZCj
o0p6hU6D3R11+UjBHPCF/PhhaB6e9cShjzMP/N19d/s3xMVG85lD/B9IP5lV
8u78bMhCQDFh4hqWPPaVvpgBZFlC+jmWMzXjBwBJ0KrzWYI+q5cksIfXdesC
BZ5LDVSk6908siZrHAGjHfh7GUM30HwEHhhjvDO4MeAJes96DCZ6uVWzxXso
aCK6RnQmv5TNMV0TrvBN/D1yq21z2o35c4zJZeAW6IMAqxW5GeJrrU4UdgL4
e8rImW8ubDmVg+B0lmt6TaZu1j1gsJIQr6oLnV3JA2KNH2AG4DlZnJRYd1/V
fEVtluMMW4cGPmWAYVlEJgHCjj6YqrzJ3sHTmkb8bYp4XQG3XgJVLM8wZsSx
aZJF3tXu8vf4wpYj+ZEF+fB9hNLflon1bV9/Y/rDafXeEEFDSPjfNzMTQmeJ
rBsDnr44aNFqbnakbxY7PcncbOCvL5NPGzoctXRzGYLcAMhsMzIybQGiJZFc
rBCMdRgjILr8wvy1cl4/5r+8801XTxHVgNi+IsnXJTLtN69GIfBt2hqVF8+r
WHDwRw8xXTpMUDnu7iGqxsG34ukqysGBpxQC5mWiXQUAs9sNqFrBGSRThY9J
ZcnY/X/lByQBig5XOxJXDtor7RGPvnCaZwMaXYh9JCIWhi7Fgrsg6PJlIPxP
DHhUbL/9zdY0LKe0fV1BLGuCG+clE7HcGPupkwpSAki6z/KxZfJ7ZVwd5RDQ
h4jh1ugxVLMqkz4HD6se1HpmeaIgm/H6sqtZQ7PuC8yJme4lb/Q9cUGDo+Iy
kfw7SssZOwbzB0P5ZPEJJLkE/SueOwyyWGFk3QDT3LkvSDYgPjuEi7PCmpgV
mAeTtfh+MmDxXwI1sY/6e44vUBTMfywtGiMjTL/bVrQbHtIWCojrLVmb5EU6
su1t21LDatsZYkE52VVxGzU896IAbTogAPQNqDqwzRb2HhEQarqd2dJLIzYE
wut/Iryprg7LcrL9Am2jTLPNSZFvFbX//HH+MvUm92zK69gQOepQh3Y+2wC1
Yimv8XFEbf3KKKYXBtKnT5OCnrmiEMSmRsro/fYyt1+OVL5MicckBONNSKgQ
GBBGTdfVaRBE8KJDcaNZCKaqnMKRo9Bm981B/zwhh6HM+D9ivZB4SUNgJagk
u0YFidLLfiAHTiIrdTxr1fXwVdWwZu1sQbakX99hVPFNjKZPZMDIKPT5UfzF
iMg3/5ztD967UyAY6jy++JO1liZWAxDUhLodFUsoOy9mnG6rOeDESQGrkexw
NM0GhnYrX2gKIJquL0xpU4MFPUTM0OsWew2CXGX9WX4N6K5C//IhplLInCQr
MNIbQo674ucmMBSmiyQ3zNDmwuWE5fwl0pqKxv5nn8WDlN65zc/kbgFLrCSe
BVFs8KHa/pRmtT2dJyeBFnLLN4BQY2gUwB7rGnHwmjxRI1LN1vuDCWE9t6QG
OD5qDvZIRr2U+gu1AKwtAdAPOxO7D4DN9NNIBl1aqjtJatm4Qc/mGU9anJsq
x5bmWncVhkVbCP5jHXy7h+KKhMgH5c7H/3bmKIr+UjLyOQ18a1a2Yd7Ua1+A
/OJLyf8BGBYhyxNHuQwILJEP9t1Cs4/nt4eFsLsDj31ULYGQwAdSutnj3RZ+
/nCXVtmB9hsgfLtxOkarLbzQKuJIHm2+/3AAd8T2KrEDRh+CFc72icNMD9Aj
MAcAOPA7taHC1HeygueKYA+gzIv4TXep5M5ouT0Nw/6e4ROynrohDP8mDqBg
fAo9poXx9ihMflxfjKIwVAS55quCAQHf8VzK9eaLlDSZV74rNFpW76U5Eqxh
NAGciQE8OcTrwbUem+l9fdVJXud1uQA0+kFuzhxFkpi1/4KtsZW4EraY8zE8
B4Va4IMIWjsIqtSIaudA3IeR8hrtOnpAvjBI73fIiJuRRc4V/R28n3k/hP6l
6ozxEjM4iKw7D8Vc1e4hkiCLL8+JvPZ2rtFZJ6VN00DX8lN8gKEArF0ZYvZk
2dO2MM433fV8BJFDh5M2nwIi+wlPSFGqXPuWSSiKLoQQK6Z/8lpAdujB4qQs
a7VQCvd9eGkDSquB/VTmVSci9wLB9S9JJAOYcTXVuovR21Y7n9sHUblM2S+Z
Iv3/Eg3FdvmfwEXxI+EL75RNIuOONLWHK0tiAtJO+SXlKjxhoz/4ePbYfFKC
YuBK8mXT12fhoHrbNImIF/P5PK5Bg/qOsU7YV1cL6KehjLm5V+Vusfujs/Mc
Yw9XNiFZKLRh38Yzf2U+9WFlFTJfzEmLI6yVuCBfRvH2B8WlKlCd5IEC1Xge
xZigqxESekeeaGM9pXhn2KxRFvM8mZB7r7JOVlTL610s4ZkzgjY4EASkwF6D
RmgdQbpM2K/mW2R1UdGlARYIdte7eA0N1ps0IL3xfxybBoSj74TcZ0DUpCgn
RewGipoJ7QMV6Spr67XaSJy5XkgAsKxQuNntfnhWFutPlitxx3dZWTEx8SAP
1YS7F0t3mUJVeyGvYyU5v5rZero8XwqkY0WPwaObWsbnaEmoN/B4+MGyM1aZ
DcVdhHE0Xw6NBwHzObP+DhgPSUCY7Iq5ZvnmNdQG2XUsKWsMli43I1Cdq/TA
PvIscvabbWD/NiZOyTr50yradQL5d/cuOzhllkQ7dHlkGRQdCV/ON2Ktqz18
+Hk7qS4IFnWGnLYfaPWyo3PeDTXTnG1Dh8zpayFvS5DkefM1xiZvB9NGWlHA
SBKxOJsTtjE0HFszUqCx3WFYFN9E1rpCPe/iZwqajNyCZVHzobGTxYsdYx3w
6Y2bc9hFx0z68B1u4hRkGa9HBIabVsHhmpJOXeOa+TlRzbXPHfr9RLqh29s/
JgG72XtXf2RUqr51ZGaUgMyVsFLlYUx61OQ/I4VJOCHq0rTwzMcLrlgqHYLc
VMxfmWPG3BdCKYZCw7RDIYr7NIs/EazYscd/3lNo9VOLhIEbWPXO0s9nX0nO
2rlWOWzgi7TQVGRHUb31XS0PRi39GQLpVM3A/h1FdBVzjPqRh8ErST+pNZcg
r2XSL/JpiVeaaqyXBOJGk84KXHpo+fBdpRVEwRRTLNkXG/4Jz/Apw8sGM7mM
wGWc3lrBn6wLDB8HQgPqrHNjQwfJBkqE4mql+iW8N54dwTNZ7Bizb2eWTt4Z
wblsqds+S7UW/iLoP//tKnu+7NxU0zQyawi/vleNBHXedRURZRqp8HI6Ycil
7Su9My3dQibxOa8Is8kDgi/KIAaqvGqWawLUWaAXTpnPHWsOsluMCAhF/vyD
zWKJ6GICEMM5YJ3xjXR2Pi1rl96gBcaemxVFIbeogNp36k53Y9Ucvoj4icO2
L6Q5hjGbXIxsPhdRmLww7F2iNNNmb+HoOJCKEK+8segmr70kHMqOkCsLtkEj
Ld4n940ePvPu4QAFha+44Anc0Lz8/e1YTOrfnYUMrGXXUFd7JVuVNYiYiG3g
lJjqrnd0pP57mqo3Ghq6l9xUMrdftYzNWJkgDJfZD6+pYu4vyarTFiVXRoy+
dr/GR3isqE4yhfUbmoUs9P7UQ5cMPs/muIeTH6PNeJK7bwkOCOVE1N4a0uKE
2XeFKt/gN8jCybPl0mi5Jn70li9FmyzI8nxWSTkUddcaKNLvhT+UmZJ3qGdb
Psj6bguR046gXF9+fpkNmbQe62/plsP2FoBACBocVlfYL/jzjR7T3HR0Wq4O
C/U2GFP7JgjKUu4yzXHjeQAUyzUFq29ZwQgFiqdhmQ3/0/Lvc0E1SVnUbE3K
4apNIbDTWXEV8jrGGNKFxkHmB8MU3MS/YsM4HmBUzwQv2/VXOV+4hRK496kf
1tV/AZjIvZXSBbyzGtirXSnaMum69SvCujfSIHW8gGfpKNqP1eqzmsvRGU5X
yppeCGAHGOHQ/vIyioYAcO8OuwEonnPlUCyGWMxy2B8xz/UIfo0jsg+AdIVI
a3hskN155Shgng3oDSR5jHSI0q2eRYxDjdMvjiLb7BUDZ1yub+V58BlvkcGy
5vnunG4XJWMNdgT5B4OaJtP7nTe+TRmN7/4G160T6tkDShTvRMBzRHYO2SeK
gaJrep78x3RbtmyftP167YXRveGoyHtd/C8DQCGOkkZN/w49tLs9CTJSiy6O
LyFSUM5DJBRyPwKNhsffJ97AEhDnSyW4hEHaBNMx4Eq01dmpvoZ/+/fT1k4G
y0lDew+c+px48vEgcuoqpyePUESqQdPP7PrnxtmJgTsyi739jZRGGmeBXeza
94RcmsJSdT/ywM0Ow+93MAFrEIXOrFLnFBmsFVfLhwu+n8+LGBBNxAgR73D7
+8G5XWgm/RnQPlqtT2+eP+a+IblQKkIq8kkpG6KnCgv01WMiubU0bHYLM1/o
AQCWbI87qnl22O0OAzMDEaTaAEH9hlMxNBS36jIhIf+XeTssGrnDSjn7mW1g
9hLToLLk7c4SGPHGFpDRwYYmtcxcOwgNLkIw7BqwN3EzUJXjSjQBGQ+aKVpO
4Qp3uArLhO9fAq4aUGRS+ycoyI96kpngwDpGOu54E9IOuP+WdE2QWiM0gQs+
FzVbM5fNqND86lolepnqXcG/fS3MGJxMPis4RlL7OqDOXMbB/AbX8/mtBLmO
uQfcOKQPbzdgp0Lwa5ZYRIwDhBlu97mnjgyjwfFssOO/rURF6Kbg2Ooh6bwj
KqCNYM/zsJ6reYpYAMu1o/yPQz5eM7xkqtyRAsl2Df5u15imVNMWVhrtsqzZ
DFF9dPoft2ijFcVW3gwngc9MVDse+ekpHnPVRJHYOi9TnfMlCDyV5GD/ONro
+2eoYG3sVZ+I2zgyRPM8TAy+3bpFR3kJXHHR4RUzjW4f/OOGPRgrHKWFRQ30
OWhMNSjtbagbsJj2Fzw7ExbXFNZLl75iaF/2xTE/TFFXrgXAl+F3u66mf348
N/XjUEM8nwQFqixujUWm8vfGNWxKVAIap3NKKb/pJMfF8XnfUCooF3eSgF/d
nYxn4cCiF/UOi/MEbEgqzg2rwrSiX5MUcuN+EgGC/NE5W3Ah9tbdWcDIIpRs
5RQobtiQP/rR2k1YxGGlUqLhfe/cc6f/2LNnsX/8kxl4DfhaOSuZUAdjG+wz
5YH89LyzNEX6BalnSARmfF98dAhTys35FKrtQ6JEYDmju2FZ3L7uTVmnI5KA
90c87RkpuUw11S09HDsfHfZEahs6jfD2ss0ga1KFMO/w4UeD898nmixtHDVx
LUkaRXhFLB6WZtaseVd5EjeA2RyYpTdaVH1NB98KLCQpnjnk2VMbNa2+wK0v
L0/X9mKaOKANOZO/dwz78Vygc0C0KxUF7lMs4+/ssl/bBxqy/s3goxr9SWxn
GgH7LS5dOJQVeoW0+WJQezDjJYJhTy0EYXuCU2ZNJGIf5xGSO0fA0DHcC8Mx
YWBbeWphcZ+Od46p36/nSdl4ydIgXnGKBlO0DlERfM68DRhGwrn+d0cDnKP4
RlSgYezLx9WZdHM/VOHWpn1hFSoDMBlDB/nxuIuHgPh8xywvbw/IYAMGDbJY
2J+8zq5FkvV2TIJ+C+OuONN1uQFsPmlfGUwhkTdJG9J6HED04qnZMYFd2T7+
D1nPlvAroErRudIic2xfRtNh0736tg0BzuWR9czUmIDZt8qT8fT2hp810rO8
kXJN8Z362lLMgH0w6YY3ciF3TzwvedEo3wF6A/ZqdRDJnspuhJdmcuNcwjKY
C9h15JT/IDphErHvykBO5o4qx1QoTXTPulvZ1vDfryHfkMNL6pHctmYIcgr2
P471/KRi29AbYIpKyJCRcz90VeqKY+8yUl46+lhefea6Wrjeqg+GkcZeYPPb
Oxd8aGxi9OcuCNrkflkGoMcugZRWdN5pz/QbYxcEFtY+clK/WrQBZOCsTDdd
0gTnvQXB7gWKlRFFGYp/7uGQPyR+l9+FTE3rrR605vA4JHGCDxkjoV57nJid
Y8FZ9frAJ0uOYA8ZIfRARSfz51RsVv6n5yABMwG+6dK/ZOS5ebVfKoW2dhqw
iaFkheGrBGppaUyyS9ZBLx7fER17o6GTRJZ3MQZse4+qjx/D/MmK1VHC3Gj8
udafz1klGIWr9w1qcetZpLeO9fnKpnQ5eMWWk0Yrbjw+vTqVdbbRzbqXjjJO
hl/rC2bXwwXv57cPZZVZ5M3Y/+N+/2CirGIWHZenodQnIqOJNmFZfII7r4Lb
NIgbTmEXde03b6765Bl28pvGusT5nxOc2DdbCUnwDHW3Sh6gCMy7hguH22o2
GnHTguGpOEH27Nj8RHm5QKBV/avGun4KD+h+lBcvtFaPp2hIbeDZOK6iRl91
OCNy2oCwEHuZr1nj3YRjL77gmJLZ1y18ShbzG6VL6N7sDDs2rE3mDToSP4fD
PptAf5PTMUExuOZqUFC6RlZCj/4DvLX79yW0XPG9Y7snP/K6ezKXyXh0OgCa
P8JYlCHc6mUbiUpTGzuYbHXtV5P1MSCdx1NNa7XXbEMlYza4pzItWqQkk/9m
TlBeZzIetKJmWUpRyXiQtVAR1BOvzIYMKCy4ea04vzLNjWDVvrW2W3G8Iyey
b/GUKmtWI4OIx9S9kVJbgdc7TYhFueuVlZKEQZVnHi6oH4+BXvBINMi0uEXB
lhMZANfj5kiEYbgL+K3//In7BYsVj3L1WNxE5fw24DpPEpZyee4gkxAIbYe1
jemF8MY6QRtS53gOVrvInAFXQYOJQjPxdNeLhus9jqI4TVuUfPz7+O54kgSa
30WtSX7Y+8Dy52nmHU7rfl71W1pbc7dYlY8QKzylag6HF+r1d5i9xM0zkBE9
oIoJ629JfZO1FODKY8pO7//EO4cszFoNfS745JeRnAGB5gy5r/xB1qXaSqLM
Gr8oulL5K15UHKEH5lvIckjvempVWnk90/Kpc9EhOQh3fS8N/aSpoiMsIbwZ
2Zg4qebdKFd4rR/ZQEad+P2oIFnJ5KmhkAamYMo1rCXI9WgfZZKIUbWTFshK
diAMXriURPxu1OV6m9cmhULAECwni6fiFgCBi/HOh+nvVgT5k9ixvvabEp0H
t3WTiEwC3zhaU5FBEH+nf+5Zxl88w7BKNmJKixL/jJOrxAc25U1k/h+MAgOY
vyrfhC/ORuVXaKGzz0PUYVLDnWvGQROxBmw1CMGB5IE9qzD5AU9UKINhU8M8
2u0D5M/7Vc99rdIGd31tfIvcCl+NPUFqvsnurSDb85PjJakdfIjIg0yUHD9m
KNtlx7cBE9sl94tmDt5DS23D6RcF5EpegRrd07qxjU/j2GkvfiOg6QV8YTCH
Qq9vKBx3UUrX2OQVckoXcSNe0iGNfo+WLfjAJwNTcaM787tRC1p162lI6j5z
wTdVMPZENDMMsu3QMvDfpZrCxwWZ2+197INnxD2E+WkZUH+Bx8dTIkCYYnX5
XOdbZ1UP5jx6SqkhNBKsYRMxOb6KhRrrEVwP659c8hUvnpG90Z2dGBBGXzLH
PMl6IPAcj+5BLqC8ElRkRYfyl59EO1kL5BmoLfG2iZxLKZyQGcG7Dus+IqTb
D4TkjjqDFDbndachOnXmEBqdoG6jawOV++lhw+rdpl0QIIxUlafX6E0M6SIB
ErnI7waP8bTJg1jE1hWzytMd12hDCaXPhWoAg+j+Mi/HZltWfaoEYzc9F9f0
+hJUtJUlg84c1DVvOAMvDPFca2PMYTJ7xx6W/tw2Jz6LKAD6ljKUnSyQthCt
FIjSbzbIVZs48slXBGnQpgrnXskxf1Y1aE/NrTMqKDQR3PQa8a7G8MW65LjM
UdzwyTnlqDkDUzzfQczQ7wy0Ottqa9kjNgePLzc4YTECqs1zSCdGdmV7GaYj
Fhk/fJKK0BQvfQ0Qk1Vrh5J4SGQ1KLUar9Saq0Xy38nemdoqYn8StOG0PvBA
OhnCOGc9Rji0iL/yQNlq4dHsHG3VW75Odc5ohlazxUQjwPfIICDGG8T+jCoi
p0jiu++Lcxwk6K4fSNEmoArxOJi+o+GGR9/8hrkGFwoF5wMo2BzbyuoqpyAI
qK/S4oTo5oB5oetOvf/f6cVD1pjLzaalqYAfvuQmyPwUpX8BNnOGQeaIWOl7
kF+ML0p28XzfEXdBGixKpG4XZ7tnLGBhvzdC1sYV9LXhFB2LTKXYCx8ZfnFM
OI1rSKT5gHXyAAjzpSREdmKTMdIAmqqEKrnOXJ7y/jOM6glILEQyfwkQlUfB
TOBeL1KwuLBKCeDHCMqYxnF+Sex9l+EGyHq4rCV26bzvvqM4TV4Tb9ovkhk2
ykaSEf1PeH46V3n+zGZOEi2Wm7QzkhtC61LD4VQUO/Iw+1VqiXoKZASwAIv6
jEewnF3EO4vX4pgb8gnavegokzqgRzi/oGUha0csGOW1d8brExl46SVfhQGu
vMxztkkOgKWptLkPF5W2mfCB51DzrHNVEiK3vraT5wHTR9a6yMhCJA/2AhRL
52sB23+Y9m52vsAzqrs6zXud75T9uhu/BUf1TGjdd7Kc97TNLTWlZbgQzdmo
iaMY+WVCzqa77mdQ37J6kgOMIijfMHrjpXQkLPF9/u1md4YafvK5ztfDmVFD
iaVfiAMBRyzeT1VtoDSOVFG4kL10NTGhBUWZf4UksPF0hqsS4recuesuR48X
4gs7F25k4PZLZ3VENx/XVSaRGJGkuvCO6Z3gNauz5KgeGpDEZLlqGS6fbQSQ
I0RWY2bk4/X0L/Z+TwIc4lhCd3pZCoKUv1ANuyeKeCE69XtE5zEtXoLKR6bE
UU41EUmYGnXpEADHqcQmnyK3LhGzJO5x4RvqP+5l510+/nuddkQYDOOpVYsQ
TquWhNGNPWghfcoxnYZ2RJ557wX+/nx9bGZdrhaPyoG8YoopgRcg3qvGWhwY
+1EInDDE+32Jx+GetJ59eRJUlw0ivqbaJ95R/Rcqc8bqydiDAF+39W6k5EyM
nVScKu/lb+zOwmy2ELtJbxyvLiJuBPOUjsZEx+7Arb1f4LCW+6Uu6t7xWAHI
VnMGrnerNu+Q5WGq21Boa7ZhPkLtRG9MzqqI5ArUOPbWzCWY1ge4TTECQSdJ
cWC62GR+vAee9DkxJDODFIvBfXfTbit/4J/UWs+w7mbSuWEyCqe3SUZimh0I
zSFu1x74n7VTT5AVI3WWteaq2BXFE9l7MFNSnjwfg18liEpGmeNJDzpgz9Na
dG7BiAE2YrImeQ/jP+DR3ttzitot0dQMALhg17gMPmoXnaaWi21u4WWJab4V
SjWGFAGq4IcOrz9QmQqxVG2oBTNEobj90ChTBGLEiRSg7WenIQ8KV8J07dyu
mVf+znQuGosJmdZcYEEEC4dd5XhAk+mr2q3n/ml6zpogaf2qBuhJfUXcX7NP
9eWs/zKWZRlpkmmNSHrVCkTIJp4OH2FYpl5yM6HlcBJnutxNOsQHQXmr53YY
3gUaWRotP5SOd+LlabobKxZPQKNiyfKVtn4GMRHyaofKeQMV4Yt5EJklp/cm
YtYvVV2DNGfRiZ9UYyRkx+T1rgAWvCh1t1vd48rcgR+2sy8hCga9e3s5yEv2
sdolzQtjHW+FBjGww3R1/rsaUG2NQp7RIsq+HsR7NOeota7fvp91GV7FV227
93ePWEVQMR8FBpXY5W4BBgKj2SHUQDNZk9HA67z6npOQHEdlcNx9Oj9gkemp
lct11VMi6oD11Zuy535H4N6lFIX2tIe6KRAeydYF7iItDffIUss4iOamCTW0
pE05JZkTJ1rei6yMFtn2sWjNQ6JxCxC/67xuWqfkgd68UcCpNqMnjZZ6L8OW
Qqz2WrnWFg+2deEEsdp78M+M0DjD21rbb55TOTF52yFKNsnVgN8uGVd0awBF
WC3NtPPl5CzK/IOZoCTB15xfcJPhV7P1mUcqkp3nTETZsReILE2gejKUV/3V
vEzxMZ4+RkjL4KdXoNQ3eCfpfAjIfXwiogT4N5gZLR/ixlW6ua5JObqd9jG+
JSsll/N4dktRTTzM64QzUEi3FboGi3Rv7dEjNlsGJrvOo9pV035q3W6/Rrht
Z2Xz6XwFNROYjk4QIZH0mtgnAAdoohqVvXZUGxvrKIiEkZ0RMKulXl/ufjrz
fBXUkwc7bvN/OMxhjrYFbi34otm4d8muoIdYbZns/dTEtsaedoYrkmPGhKSc
2XWwbE8sl8f60PFIIAq19h8wPfIbDNTjbcS6SfYqQEqzOJ/XOUJhh00om+Ui
eTJwwIBJcNZuamYX8oElZy0uQVWgxlxNeiEIdJTFeQljafk2Qu/APnkJ/XZl
NwhmCDXDDKwdh8+SCm8d7bmBjudI7RTv7f57vSEJZfUdTFcBiNtDdTFjhe0s
E9972nrAxhWvpipORqKmyESqMp/15OHr7e1HVZ411PoxAZWdXnOWXzcXegW4
XsNWHpfD1UllYhAoucprDqoHWa8KovtJs+Gmi45jZZRmAuvEYD4lXa4bdpRz
jFjMB4i0zBmMri6TQnnyiZ+vboFpM2Ts9dHPfRGWsEZDDqWuV6ato3YhFmtP
BwgmQVfUFxJ4pf3IrscZJIoTofbS6gXl5UTDtHAuN8mvqRKMnEqdbzoN4Wen
65CJB0rT+hrKAPsdtzo+rKhimHK1cKbpOlb2y+QxVhfof+U4Fvmx67KFZC9Z
592wiqYQ8ipDaak1hhLDT0y1D52F6XvmphX5K53/MvvMLADmCdjan+eLaZia
0UKeJrv8RrrBc6QV+WDaALNSemQGAMGhubpUv19p1s5DODzopsDnuf+KR4WU
iaAD+FTwIaOoDLkjDSau1DzcJOD7hUL5mHQPa8eBkFEak5l4pcH9UJWD0RFx
LvknltIgjr+ZPH5oGkTtrajnSFwCF/G1bGK983tbHiDBt/fNAcOyLAKqxM9I
fakqgX4GeFtlGaCpThjn5Q3pgbWXcnM7nj49K4BJqSaSugk0+LKT0eSqDDuu
gsTjwx6+tIE0trc3VoPEerdMHGjcq8Ub76PdhP0JCeNIdyRDOvZzs+OxHHdz
444ZhgIDxo2MShMDwQ4aVAAorsn/DMhP1j6q+InygqrduW58qRdgasD5IipB
kMmEgkZz8EPAJgbinA3h7g/31di2YDvI0KubuB1AXnJTvgju1ZcEh5CMzwVT
Jk2TaldgpsMRZYZbEE/+MWwWolD4LaIPz8dghn1f+qO4SScDgwESrk2KjyMZ
XIyB7WQ74anN/2St3APw1DVyh08EkrRol1sr/hTGDLBwci8r89M+QdUG5SPc
I89+85wSwqrPhL/GA+esFbvrCGYM+ONbgn8nO2WFV3sIUGA7gwO3eqdx9mju
I9TeB5FkDSuBP7kd+/9O29ADnTHnV1iPb25Pe1O6P/w+Xm/Mfq2wl2en9fdb
2wtuYcA8/EYR10swDiUIhfvjoYpx06pTN+XuQURYM04JzuiAIEFkR+PvlyRQ
IDE2hrrbpkjmASRxIQOuK2YxmzekkDek5eUM61ne2gTeuCKMJYlmZ/Nqr/++
DvjbNGLmFHqoPfY1HPtXACAXeHIVojAyNuSr66VG9QhpFAPg/KH/Vt78qLqI
eQVdKreETWT333+8V9UYk+FyrafuPbLoOnx7/7Y/6UxtBiWQjV+JzVcQiIA3
XvivonPxEzp8nHHfi2g+OsUPgwD7JPhqGFdkgawxXcCl2QXm23wi5skEzGAk
SIckfdtE2wfrBG/HBB4x67FYLCnJzVhCWyH0SUe0kLKjVKrUwJfGVhf6K3p2
D7O0hFkurybi9PKd3MnNBqyVoQZJ5DEZUbrqmMl8CuZ6dDPX0Mda/TiSPYUJ
NgNzVaPHxVt0ijxZ43YWk5sgFM8phW/YMd7n/u55rLpvgVUSjVqrXzvDf9f9
uiXimUT3w/cCZpmwGq8JRpwVLaF3ukMu6VCM9dhMhqEsRBgZtXOtEoeKvS59
cFgZoOEhuCTVFbdGw+NvmytZbERIxNjngZEnf4hB4kVFF/Tb6hMFvNFSmZWK
o3SlQlV3MKe/OUW7qZn9ryaob396vuKw5AWLyWHT17Vhd0YCvN07muZRyVHX
J8Vt0uQhhl8ljB4GMC+yRdPGOTuIUrse7mW4tdrL121UXhPQU6K4p8C3OLDE
zn9R9HztgziMZtckw0yIRMZCNmcpo/IRWDCS70wcjCZUuNXn7430c5tQPEGJ
es6lWcHx59e8rpyZAxfHfeLqWk1LshUTCZxRwnbhOC9ev7YZn24VIJOR7Zde
EbNpK5La84NLiSE1KJeAYurWOo76PmEBxCPtf5zC4VxG4W09wza377mqSLwj
4wBcMS23q7lXC+zt/UJVvuP3aP8yfW9wXqdStuK4mwg/Qn1peDHHUR6ZiEOp
bnrwt//fGEpq5Subl2q2b0r7bKl592PqV89clWhE9iRLJYxwLhOhdEmkFa2Z
rWOGOS5f21nM6AbB9Q2AGYCHyA9NTZ0UYoR/KBgeXJ/dkv9oKs0kGEzQPRAW
sQufIEwo3JtmeGYO8V3+k0mq/EW2peXodPR8Mh/SaKbFnQHw0RriHVzahbh9
fcEcbs9VzHeiEy7MDFnosXB1f5876SHHNVMNo9iwsp3RZ7Ndkc4BwYHLsdrc
tVjbAucgfUB5dcrOmoJEtSLhvgGeP6YgquFWnoAQnpuoKwCE5zOBRXM/8yLu
VNhSriYCetod5rngv3EJRd6j15OyUlC5Ln6S5A+cDuXhnn0dvq+pu3YVWfCX
GS228Y0GJLsMgvqDT69u/ieUXzGXq5sawnl4lJ2nzQ6uOamoKRh6baOmVu8e
skpI6VKjxJOmu/RrMjvfO8XZemi3DA7OP1fW/nEyH9c7Dbl83lvq53kM+9l4
E8hwh2GeO/WijhaMsWz1B6+pZ8b8YELz00dydhl4XUxL9Zp7/rAIela99T4q
EdJJrdNq7AtjFlHbmtG/saNNuLrnNhz4DJMpQFMOHMprXU1rM8DOgLBDtXBC
hx4aPLj6I1zgmY8j3u1f8nOqI9zKrksDp+lvawdFmlHz38UFcxpJYM4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfTb1bmKPAEo/g7v+wnuuAY5PaqYKx41LVMgucrMKeY7uN6EO1EdkAvOZiI7OzSi0w2Im7KRNKeuQluf2T4LN3lUZVwzuKVD5cOEGbOb6wTSx+td/4J9JMFlmtXjY7g3+evu0FIqOsSF9T+Q7b/WhMxE39hIfK+/mgqR+PydKsSlHbKTVElyLMN/YRK68gRWfqbzAOEpNiOTUYmkyTShno8JQc8w7FunM4KIZDitOkeHMIIFShP/GNORzfkT4BccbmTOJL1jp5PAtXO4yVysrkSeA//DS0LRwlPQbqr5soFRyKy9IlUaqOODfV0x8MyVrm/vk8HuT68FRoEXbOj53yEM4I6dnOtew778Q4svqk9Qk90ljhvfAtVggUq2sK3PugYNo1SXIpS6T3dFwB0LKtK+rEmlS8N4l20Dvg6zQhF7VMuztATYwTxvk/8bcCBH4dgkz7lgqKoDBHpe5CVm36J4uJ/LPUH59DIIaXrflqFYdUCGMHKL9BCVDk2ri6gviNMdAm3wwn34L9f5uCuvdgPVLh027QAXhb2HRQbYRhFUvZu3jT/YVnDcUwSR6LypeeCcckkGllt2gxZ2jZKFt0KR/7iglaNHwPrjMdNWgP88mAKkA+tVc/VBLdit4IImwzAd6rR8vZH8xZ80+PEYghnTj5AqVoFUmbGXhYDAAc74EliVkor8p1IImCLwnkdgWoBP78xqeRqjmXnNrXTJA3u6fZ4MepAKUTpoQf6oMWhNbjvgrxm6489M5Erg0WHdEZt0z8l0u8Xb8qw2a4cgkfLi"
`endif