// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
GXXAGptmHf/WLZfYSKCgbGNS91j7CR5YQp/goEaLxmd+eKd9JCZ8pTUenu9P
vMMWxhU+f0WH4Pk/p47M8EIhyZ3spgfZQDmv6GnKZ2x4EAfxMoKaf6Pa4CdU
unf3jziSlSUH6yLqZD6sFdm1safnwcqBYovicQe2AyMwI/uLLGp335QfYaqK
oSZpsO9TWLBH2Z7YdQrQFwbFPA0K8BTr7BUXejVLJrpI0A4b/toLqLAck7xY
T29WCVWZYUO6w4MqStbBoSVY8+EvGDEn1MqQBE6qPglISCEuRlUY1xXUUEyZ
j1uYxvHMBAaaGRLD+hWZIddeW5N/CaduodNpeHMFpA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IHORoarbHMBQFFg2NSPVTlARVqiib0ewL8vRlBsfIMlgL2lDuuJaTnhYoHXE
qeqATveXRnE8FfwNf49swfXE/F3bePMdXZPzAlaZ/CqBk7pfvUz+m337bAue
FfxzyEHnqTD/X6bXebLWyE940IgXKXYBcZA741Cc6lOixLriQdhtCEsscpJ9
kmiQ9k6OYMtPUmfgZE1xGtwoZgT+Hd5EvDKyfJ1wHxqpgTLqGRj0zPx/MhOq
harpB8OYt09oGB2VtTUtCGH5rQnBchEiyFZOk5YgBuRsq9M5CREu5ap51Xb1
xAzU7n2IHxn8usoY3lQJodAKM5oqIRMq2ESsQRi0TA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ggW98XdxGB00dscz//fCcugYFuX1I9O3k5uoxLRg5d5MRJD/g5GFykuh8E4W
tJb+3JgYU42C+jKkkCMsvqC+tnToskP6tUKUCaMvPprdxQud7MPHVqTogRB5
29yDATrfnfIAwzwe4Ih57r8LmAgPXxDMoIoFUHzt2s6Thwl8Bpwk7j9sIkw5
GolaDA83ztOt63ZbAkiLagEJFyibk9G/AgnaY9Hk7ViIJY5pkaoX4TLGQ6ac
RVy3TvbCvx1vGxre8zsCuKwFOmkAaMyIaceBs918by7QFm4iq5YGOTo613Lw
uo8/fG4/s4Ec0rXkozX7empWYsxzmW0aMQ0S0jGwhQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KltQMgB4Trf52G+PoYlYNDDm/emWrxijeWGKNDakMzNkXJ3A/VIO+OqZRVeK
m0v4Ob4E2K2mAjr7OCdYbJT9+C9HZaD/WqNc0ll+ziZ5CDTzttlTlYSz1OLS
4q/XN2+KsAg6o8RdKZG+cKw/K9ls9ABQgwPpX3BlK/EOvYbeFTw=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
yEcDFnBF0SWFnBlbwlECPvrc1ftM1FCAAVvQW6cLJ3K43Jynw/U8w+RfoyGD
03U5/28edidBBqDERiDRJLPyNrEJZVkx7FLgb1tquokAgbVfyHI09yY5nYT/
XLpPcHoYUFweZLc7o4OA6Ve+sH9QrDFSY3lPkvrchck0e50BM9vRNFUDs5ap
kST0V5I+kiMS2Rd2stwaUxu/fAshHnTsntlzD1LLLsP1V+Vud24laFWuXUV9
0qA5k6icjCpoEK/ZoE2+daxYqVqroucuXpQekSAf+1S+RR5ABiGVZp2HKg4V
LhOi/XE9jxOpyp2Xw9F9Y+HQDcDNA+w3ZYQQma6rIYZGmwYpemyGijRiAe2a
A3C/71N4VSAyFGyNdgBaFl6u2hyACfysop928aHY9QgRnWW3WJ2ZE1YRbefH
RD8UBA+Yft4Uo4hZGJEnEtF6IJBgZkHSY5FBph6IqAlJVu2gYadZdepKEJtq
tuIn7IOMpwKU0ZehoKZujglQ6xjAzIby


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Rv3DVWy2ZE6YrsUg1tVHl9l14cN660DicAchLD8btGyVmggq2FevhBVPA9Xr
uO/K4+6M4chv77PlhwTyrvfwcuSFoUsqU1HkcrcaGi1tlxOSSCEAwc/iQ/Is
dlhdacg77xtsDBX2EeG0Ixy0njkoQi4U62eYr/CPIq6UioqhXPs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kHd7JsvZNrXtHS8Y//wkrAVX6GFTOcT0hjCkQ6QAlRwMMQYDMbwVeFYE76QW
lseTsy3Xfw+ghSNKGdfCTOjxiR660dQT3gnP8aMRD7m19xOuvEn+fa+lBa+y
wf8X0s6pX/rk0OrKIKwdoBxVL8DzApu+Jy7JF7ZUoRHLMbZoyu4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 32352)
`pragma protect data_block
R8jks6J7cn+5xbkIdUyn/2rtMVOIQD/yDyg0NmrB4/nA6so3v+OpMzPmXR/0
HvCu5yXPVtK+noccikLmLyXFwj6DF/OcAU4Y0OhxD0s20ryOAR/5rQm3Wdef
K6n/S3sDQoYF3dMwZEIUr/ppxdWkVRal2RwYd1wt7rZxstB3O0uA6e3NngGN
cnkLLlVT4HDF/Thi6/S+S3+lELzhiozFhI1vzRzpHQ+WJU37EQUsytNA1vKH
Fm3aALPbrG5NuNhFXfyMPWU5jMCeNcb0ST+oZSlcm3s8hLQGB9XvweM5YYzx
MgpUNIyrFk5sQQh3MP1JYhy3dVqQJzDqzNfN8XMbRMkhyAYjqeXJrw2tR/xX
GEg9cFMQfnK5a3Tx9ilN+sqgYewfe4D+Qgof6wXaTZUuMmqSC34hUvQM1Py9
qtvAamSX17nxifpw0rq0WfKdwU5DzV9AUoo+o4Gwk3GAXbm8hiIF/v4sBmbm
FXBRM5PJ+DMlBuzz/v2GE84ZZ9MdHuHOMUK02I3s2o3wVOzn6Ew++43BFXk9
Sx714eJYltHpbHXmwBf9az0xmU2q94u5jYUtE58pAr80Yv05Q6nLd+Yj6yV0
c+5bNAjwpcfST8uBclP/CifF1Phr0C4yTKlKkNf7cso0zQ4Hj1+DYj8x6mru
CEX2gZdCKCfsuj/zEHJckSSYejfAtF3vw+pustxGqzN4yZFloDyZoYpHrqZm
mTQOAkd2D7VmXkCDxxlQoq/sMQK1Vwdthny9fSOuYZgJLsHb2goFPikUL4JQ
zdTFxIjDctMKNDxrWygKIlfict2W52TN/0C29KeYeRcv8Cpkd+61CwUWw1FN
ouCaEYGipru/NukhkvrEJ1WDlSeajzaa6u3oRBBqlY8emAzjmdKZyn+HP1fR
Jag5OM6QkMP52rm1p+brD6HyUJleVTF38czsl5+P7ajNjoQxXz/KO73Y3EmR
OdH5YP9rHXxUrwYlMPq2iWCbMNxEeL//MAVksB+vfpyXxShZxJaOIRWw8xRn
NGhjG/q435FRSJWdsG5Vo9IHNbtTY2b4TyP/Auklo9mx7dZCb6wG1kbqBCtp
nitcjlurIrP2RnD6RC0XCr3wBN7f2D1euHxNsyViQYw3LqoUrYZfQM6jcXlK
ovfkkpfA9jbxqts3TZHR/8lzCve8afkA+OjeYS953ioQ+YPyu4CcSUzmFPrg
pWXLKfumx1+hG08O821JGZyVVPGA0CWqZk0n4g7refLl/gcXZ9RTmDCTBR7P
Zv6IvZ1gcVo53QRRkCK5vOd2apKJCfRnJMFlxw2GEwt+CewMFrU3F/4RvSBI
0nB6BiBZnwqY7/aNfqEKrU5LBRWTdU0707WZFo+aDoPWpeQQNS+A58vDiJSk
vOChrZvgjs1M/mHGzR9xEpawDa6CuuDT7hvlpoEp86cVWEzf37nqc6zKJ6uI
3r2oHfcTm18eUURR6PS+GHLFbBzp2w0Zh/OHuHXbx1PlsVXawV8EHvmC/NYn
1dHAyn26TcHOF9sxaQVzOrc8PocI4m1bZ3Aw3QqBb+m5DANY8LbieAJk1Nl9
XcQ2IbM6hztoIj25JJaLGz5tNn25heKIk0zvtcikdbNy/EG46GU1OMzfkn9L
YhBQ2LvQiHN8ee/h0H+oF+PMsGR/RO/GAQK5txObWNFs1U3ZfAtORp9NZrjn
re2qJLIEGpNmD8+C+fGQ2YkD09CCwbD6Cty75QOgm/av3xKwMeTG977PKbVp
LE6CfdstjIRKZlPiafpoSvNNojcVGkIVv2J84Qm1UZP/GM5Xql4i5xrVw4qL
kPW5LoeKi/BZbnhK0ckd26nocpEvqdPsKP1blJ1FvqAEJy5zliuKCWx2ukzv
7Xzuj5e2h7e81+hiFiJMqoGuoI3lvX1PdMoIZhygYrTwnUr+Nzbv9oIDfuJt
cVQVplbIm+kKVrhI+a6dBI/QWAUvKY5yZNPK8KcW52xl4ctVWVbyRBK/Zghl
LUP6z+U7LnGLUsMxA4qAjgIARAEfSUr/9JwAXa4a+RAXtyyzyjYP0Yg04Jvq
ySM4z9PNMu0suHu/VJ9phzitnV90eMGkzSCCyMqvzSfstMHF1nWf+WjbOr9S
aBDkyYUxSNVN2m6znLph5bbaz5KpAb6ewZ9vuY1vsa2RebV5+vAycLi+ZdqG
BjwJECoOaVYfYK6hGqmYYa+PZzhpPhtlt5OrugENNlVtsCKGabhyFL/5fJfN
G3aWls2h7P7SGNSX7wrn1VNXSvC+XdfYVmNoeEBR2rrEqz1BHDsHzS+zbZb0
Z/W6xTdmjHrX08bUolLzhZBKn9FLPvJxh3cZdAbOrpUi6Xqe6gwiq9wvz+i1
Vi26TJIO9efOYFvfD8i3lxtX/wNGKo+wPGhp0QEjcj560/aMsq+uVpXkaT8i
ZFyupCxR1MzXKvk5r4evwJSsPyLlIjz7Z4Gmt5EHOCSvS94rWdAQghhIuqUS
jEUVVoI4s/14+oOWxnHoDl6i0D7SVjo6IPlsDASuBmhg9fTLd6GO76OwiD4D
6ci/D1p9qU45eajIvH8MMxhGua0epqP+MIiublbMOVtDGLMMLzgzDoKNJuBG
YKOkZMGCK7jeGl3YUOPbv0T9PFiOvLhcsuan0drqwUKpuxHIrtxdujl69rBr
sBzEm6Us5fChweCtzRqY2dp61aTu/PTOmYSeaJFDF2ui9qNcFi7qphxFlRfe
j8oIAYKrpCqAcaKlu6HKsOHGvyl+5LK8U4kJTjSMWoWyhd/89aE+ziM8rV8j
rbnTzwELS19VzLvhyPjKSFnMlf+HR4U95275EEh8xiRroWmcbjnTXoBpVNKG
iedsBwjk2yDpRUooOv/LSAD4laHMmLe6dMjDvetLEjwNwvrqdeF0H09MCCl8
CXD9U3Faqkbb0roWwee9wJd0uK1XR9OFCLw4N9GHzEAtrCPopTTqj7FkLx7O
TY4CVBlPaxkmV8C0zvFWOln+OxaapDB1zDtd5KCxlVV9KVnCINasxYnKCLzw
c7F68sKu9tpb/YcKWd2DM54Fiqhj+gCMKTjlQVufQqBCxvYydMGKBq1Qkefi
ZpFJWQo5sb7VjKHYrhmBJ3UN2JfDpIcZS2JwoXyvZItLmBDHT+sgXN3CIKgf
YcBMiahuIx+fAmjt6JQnFlWMCe6A1lXQr1qJXpSoxSHT2pENIrZxXb1e936K
TPNpkp1r4sYRrYpYSZMPCqBB+veKOvxf1I4g9d8gAgjzyVPVuQ6NuyuDBsor
oH3T0uPBpUmn4gC8yIuxfefxIX7s18UYrDo2Z9jgikNCYxgW4e3Jyup4Qrpk
9WnMie5WodLXujoVx6Nq/F/R5pNMaZifbTDfYYw0m1jF+H4J22NBlnJVM4Kz
luZnogJlvoDOjK0wQjFa3ycVWeq7i/pMZBLj9QJ77hMEC3M6VpqPHALeqQxC
4G9xOQXhW8+9Ep17LiPXufEMxs20a1b+6yzfJDomsv41VRqWELoTFEANw8ea
iNE+DKA3hxFQSRAC2nAJJVX1l3sqmzu4OP5M82MLnyTXD9IavL3l+J5rp4EJ
3h/DCnc1D6+rh30rJTleb8FowgI2sXdnkladNDKMIZGVf2wOvublCnsBwgJ+
9r3VZ01oKJkp74zAUp/1b4UWqE4bd9MKdEfB+zgkQBrbUcYUWbm62xJtYmEe
NUzM+ISuUKNrS4VUu7JarXFI0tclj6qkxPTe2NLZZokV+0ubRUqygi4T6JhZ
5NrNSQnM5RHCUHT94Rz6xi3SLnWmIfyzrlPdr/ZaHVWFMhpJN/Gi0teLWTbr
HSS7sWkihrWI7aRM6tyiDDVtGJtPOfuF5Be4DT1QngTLSPIgeIlsgAzNL+B2
TtfcAS86C4SjhQ4b9VCwCTXFUqyswYuoeIOPOil6EuC7/mZnMj+kmQ41OaqE
XIR8vsCSpkUQfJDIpdl/zqiHowjMVmlf/2Ie/nLxQyI5Jn+Pp01lfmJpLq7G
Ao48N41BHL05b1rn5m/8JEOFibyeECVNND5z5r77jSx97SZQQVvzE9RrdRBB
Cel+c4gyJq/nzENSjjOfOWaELHs0cpvcplBYJK8hxzXyHTEkv6jn1TxQIb5H
mxwoYaAwWGfy3ijA5s8atwKBFeoLSHsNsnRku6QaZzIpZbKnUBfnp/bQl634
uZHeX5wq0Dbt5CVENo2mokgsAVw5u2QTOolIvaKyPpGzZzFso0TQ9kG2pA3H
eUy7fzgnd0cJnaGtfv1DOYO1MPylGH8BsxK9EfX87Ae/DGhweBld3ezflD9I
5U7J10ngNdwKU7YSiwALr6Pl1cbeADRMvWxeja8LQFm+f/rtGvmc8qApKGDD
WNzlkJ7Eb+nrPMwNDfwrqRGN3jkFWu4QxmMDPp2WVtlzDDsjX7FvMgcAy2Ue
1d6JiMO7J0uIIITeh+2uc8y8eMJN63+HZ3oduEVLzGpcEqGbTiegIhv1azrb
fVuT3KsTKnWKM5DDXNAQudGGohszEGbPNHj0QihaXsfuMi5oZFx8pob2WPmX
WUiZqvAmznSEueOYplWrIf8HV8Qi91SIU8H2HDzuUMEsrRYf0MBoH7Led3dV
nl3WjP0RVUSCzRJI8kr4Luabp/2GtobpOTisDbXVcdur6tRLzdCj3OZlmxi0
0iomDUWRKoZ0wbkh+ArfdvKmMOr9ZtU1yRRpI4jtPO6VzpnUqQY7I0tF4JK/
yz/JN3wTVrjh8kFukSsq+3WgpJtFCLhyE76VXYrFWT5xCnFMyJAXQOQB9zTI
scLlSFrs81cu3FBaF06hQ8/NrEqPr8plzInUg187FaHIUUgLDi2MM8w0FpEG
O86m1TSPCyqJXhuuGCLhc/9A/LCLGjgywRMec/RNXdESKxZ9kMkMCtWclLo6
NYg+rxGBI6baVsM4DweB54hyWSWjoqd6pFldZKCHWY6MAr6J86Z3iYngBOIK
apukU8db1prEG+dqEOk8kh+p3p5xIoGmu2YkvHSEVlFEARCmwB+mdas5effk
uoZscrzsPf5b50Z2GYCQMFcbREWKFHY+5fWiXMHNgks4v6LjAnjoDAjXSacx
nBZ1XhATEO3nm6bUFT4d+eWjKD5B+n8n5PMkylBbj1hPrdMyQ1sacHfZFdnP
6ghvByTPvMa3cw5f1arsc9OIWTscyM95bnkVUBpoK1ApbnEZHsG0h2zFUyrW
f5DwZqEZ98H26/JHgL35QkYJ9ablkAwHfH/1cYpbz7DYEINTmf/F9xIvorxe
a4wnYX+NU76cpERB3vVHCwf2UOSw2y5T0x6c80iFubh+6RMJeVkuMk44fs9Z
O1Ksy3OBfJhhc4aPWvHDsq/UI+4KmDMyz6wpX97R1NPo8WjKyBWFi0CYwSd/
ZOmzreNxTDGoYThBI3awazP93eHZBDqwC7SVBd+qiPsfYl4nUJSPYJkbHx3S
AcVvSNKFPA1VxUjeuWqDexKePEDRlx7xOx7XGf6ds/auwLq7REYO+qe+LWdU
TzP0Gu6hmgZjxQH5xayXlCltlZIFuNfnhll81BiylCWCPzHsB8E9PLZSmIPM
f0xA6IXmPLGcluo88Rfg461mvMqrA/iIA6pkiqui7fmWHSyk2dn5UsU8vz9k
d7jQhmEFK1oyDmR5IOhMxzpBh55HYtcUMtYO5h3uldIxgsZSdz4wgqoFVW2v
DOQGTSgIiNq+y5MdasTdnRb6VfCXlY5b50lj1LCLLsvFLhaI3oziUpECuODV
F5VC7idWMo6AfiaBWPNR3q/jlsZROn5vjTPr6ns8dMZFPHuPhwZ76GQfJSfI
0upHb6Ko7w9gPtbaPEoxTOPU0fl+vYa7nXlNbJW6qrFOA33ZQgXr9z1N7qU7
/zvtXFWDG2HlEx5cMNNPwqzEdKtCmM/N9kirBoiOVJPxHA43fpRCIN23N9Pz
YywH43amHgNVp+MFuWMPfOk3ZbLddTD2cq/sE3kE+9qlE0Lv7kCNVvspFQiK
82GF5kD89djHAeXhMXuaL8WNEPxYpwY+MQT6o4g9nFSlw27kH/dXndWdMGH2
3dNX8tbt9uQT4a8n9ejSil58SZk1gfLqRrBnKxiA+t1z+EEbS3ll5oS5jZT9
IIRxDnJMkiriZqR8PKDosvcWmfiRfTjLq49gjK0N1jIC0O13+IQTVx+Hv/wn
jxgGep/nfQGQM70FV6cJqc7AZ8m32h3YKOpoiKxT5N5RUybpE00G1gF4zXt2
Mb5+xFWFWv+AorDqKa8oW93FaKxaHK3Bgj0JsURLFk3UYfi1CfBv9o7UJspG
ElZFm59bz01v/QevVXYrkCmDmnODiqSeK1iV2dybZ9omMID5yvY+ZFOTUaa6
11AsIk47IzPpW1tBSCU1wZKQhKUlYbxzdaMxkL8p6AyXw35c/IXNrkubi5sa
LI9uGj+xXF4Z2xf+LV3+zdnwk9hm5OVwn16ICNM5BJMqnRrxvqsgthZKd3BW
Z9MABVcjKsUCumwnbr/5j+/b2babQyy3sOewSsd4kK3HowB3CG0nohWV9PPr
iRJl1nF06iNrkv0k6rQ5WcGOMjx+QdWKHQOmjb+QqJRVuYgxm7K2cJV8s7q0
XUVv2Zyx1yWvfKr1qtMZEQFLOSYwWvJBBWv49n/01mNCKOIWTNiX3T0BvWtt
YueSdEbt+qnfynipDuglLrd+yBvNrBmbXlNlJgVLO+IXC3sKIImw7BwNTMS+
5Fvdd9qCApKw92syg7ZvgXiSgH1DR1OyEc4g2/70AvtUGxguE5mLcqoIC0ex
3giJtAfXUgohS6d+DPIlD43BuZqFvBiZDWFgnjhknT5yhuO2XgwyMZYP1FEk
uSgkmx+uEX3jJApgSl4kRIkhGd7SqYENIqP88F7PSZJs6iGul4QMGywDuQJZ
WWFscws9A3r8IXzIu1kZH+cWAMfKib1diK5vLyxWBr/ciux8LM2nQyQZpxlT
W/WnFRQ3KncfuDssMNY9e+lQkfMYl33IhP3T0syk6EbBRHwcv53LBRhGP0b/
C9dis1kj7IwuK6L/q0IfhUQHJBvWTHa8peRTQRSqOsbNR/3IkNHs2FjcgVL4
/x7XTiROQHQLFHrtS2NQpd9tAkLPizGEkLdYw72/uXJpswGYWl++oTCRdEer
5JU+3vH9cg2j6c1l9NWo+H8r3fLHCwj/mSDjYvT2DzQlkqFx9I4+JCh+0GFh
KqcxPtPx/8BftIJTrHgbrEBs91eOw5zFYtvXa1l/gfKZUKBkRm0xxjkKw0sX
DPH805xiYxN8e0oDmEHhb3swAbtItlb6QVC7UtMRihyj3kkpLF+hhdpnYYuz
3XfpukUmpXDgA8uU9ixCYeDR4FI1exbMLnD2NfbF6uf5yia+09n6Ptvwp6Ik
wmAZ++mQbb+s9EishfmhCUjTeG1Slj2NJjyi4l8uFxsBw0/grhdd8L54xFuB
QLoSXaY5tgVp9WnNrGuHNVfQdFvmO4d9pDcj72NWXjEbn8DzU6eIR0gW1JZ1
3wxZRbPlMC04kj183imop3QBGGokoqeg/yQF1nPZUWDiKzNL5hXSsF4b36fF
J7P5WUmqLOuGmLDoK4yOKnqO3AvqlT/wt55gyJBIKpGvjldvSEZMQtJ9xUEO
+jnHXYEI5FDSkbshB34uOG/ETEQ4C56eUacBUMop0U7cY/TZhwuT0m0WN8uI
oqPSf6dtdKyqX8Rno+SCqm2RrPsQ8STdu9HsogdcL5Y0gtCJl9WBOc2lh17o
gWEhCXdhe30Uj8suh+jdt1olUteAfMopOyJRH7rGZA1AIOOUoMZKC1MQ+07+
xhSnS+9zUpFVxc24mHxuFSR1NCRSw2WaJxOmT7hOsZExG3DD7rPMikj4MKg+
ywIa6xTX+4K4EPI/95C6A/KffpjnczJVg1c6Ei8+YXh1z+esZcsPCBBUMema
2npnvV+xOAybBcHRjgW0Zp8qBYZDktoMAVU7IIZU5pMttctyw16W4vxMdDQI
lF4ptplP9Ay0lj+f2NrEGTvOSxfcwNjfx0R80Vd/oqC/wkkJtEscIyZv8VKc
8U9UEI4GJu15JARzFZXQwgoRqBB1m64cbRI6jxXrjm4Rmufb06DLiUaAcEy8
IOW/vcA74soql5qFoy1K+9VgclwgOi5EwWSBN2QC9b/2VTbNmX+pMf4dqu7G
Pl0S0GtrVEct80a1Oy5die9Mxt7GCBHBeF9OS7Tce3/H3eTFYB+Rvo0y+KUv
/SCCMsM/O1Z/yCbHdrf1yL//zLmNALxWrz06e1K+l37k/JDdKQz4FGas3xAg
wMTa0OUtwTT5Oeq6Y+3RMU4kzN8mq5Hzcb+d8Fa8wQ71KGH/Z6KPJtJ9Q2Fa
jyF/G45pU3s7EZJ345FIDn3InIOV/M7fHyU8S3ef687+wHPuCT2kkaAU6Hy5
mHN3bXCzKuL0AJUTJuYkj9ejkntAF4MRQh40IPMlG0TqTNVgbo5ZckzvWcox
1W5ib1AKgK/RgCiSYbXMibvdxpPvAXbbx5ftH4xLIaC+2zn5qKklYLpUQs1F
/MtY6MPiskQttBym6gl0ZIcGGm942zUPk1nRBNQKjPJKpVUHM6qgzoxZww0d
Afp6/YdGDP85GpGZu6zb10X31Mf0ZYXkPaGITQ9BrF3UuZNUqZbYgFkkofWv
WP81+EIDoxbdQMDZ9Dd4kfl8eGGQv+1gmspfopoR7iu5blb7F754L9OmYpp7
xB9uhxZGCWENrJ81vUz71nFTiEvZHobCuk7cUmpWDm5O0n3uqkvllE3MpGbA
jOuZ4uYKpSPbVK/S7SUm4gpUTLsUszL2O/XvUynraBodIWWQ4zX3Ggydjfsj
qfldVgCjcT1PP2qWiUNJynk4kSrOxK2cGuFSUe5xapXqifNwxTcEiBd0tHLX
a/XxWgukHasr6vLk9K6k2BebtfUlfTwZVWg7FwQJIjcKupw5GfdUqjKyLrD/
xQQlljhEbTdSr3MHr6rykQ1163F9fvB7Kjxc8N6NEAIGpUVRWrXhcmjrO4yH
7nyqdwtfYE791hymTLtzyHETScFbC3Ya13xvk0p9I/b+4hOWLCAZw7vDUEvW
I5RnJRC21eqjmN7HVWfQ4Ed4/kqHIIfv2ayX1RW64tW/VLh+EKQeey1o/q6j
XL5ULXtngB24CqzsnI4d7vv5r7d1T8Uzs0b6UBowHePLJClzUg7J2KUtPSF4
8jYmI2ZAMzLAhucAmuVmwnE8P5P9ymG5plpctVCIt2uoHpJ5vcTwr/R8PyuV
nXrCcK2qKSFPmBN+SWfEU+VzKMG6vwuVREWql/WfM3q+uDmy//LoBU3H/AGE
MR/88gF6d1zNX7FqCNrRUmmKzdih2ZgfwBQ6Cti3yHaDXSk/sp6mHQBioOBc
PBjK1q0yKT+lblb13y7BqPcyyXSKojIBUVdmTQOAZznHPKLkFkjtoPpDhF1G
lZ6KX9lA4gxGdGjDqGaH/Kdd+yRYbezxMVAkP1JnyWgzofkiwvAq6qh7GAW8
HsrP4QnM/PvLDxbbJbzQMpsvFOaaCKXcrHA1f3KjP42fRed0hj7192yM43w0
ygLEomKT98r1nb5znL+ENE/5y5KOhKx+syLOZSdKDt8tVHpICzMAJznF+CFN
DpOc1Iw9L6stP+cWwF+9ymh/DeyddTKwyimXE2EFPPTzJxx5tABEwqbNpXDU
qGTfqUgDDIcLUrDcEejXcHAsTuwt+osNNUAGjLoqOxcyZkITzWHI3+WY+SpI
GVD62LcIz5jSC0TtM1xucwd3LazPACMDS53sY94EzBky3VGzrM7jVrFNVbAI
j1bcSE155oe/vGT1LdFLGD6QQ/KzBgj4AWN2eYjWm5kTlQVqfxv9vtj0G3KL
V/pr/CWnxnNAAotlmHuh9bdtaLgLku4Dp1k0Rrgb9VVnQ+gWIknfUKzSZ3/A
hRYu6V6UKc7jImUbybRZzS8UwE7LLgtB9362LnkZ3X3dJ3dPOJdTDqLgn4ly
iEMuVmoKFg4d31HsLDnhlv6Wa+Ypjeg+Dm5wBtlcXNeUa8dtT3RY7dCtslAV
+1SzjQeAP3zoXShR4NeynsSfxeIE0PtUV9RW8iTuH76in0oCK5eD/d0AWnpX
CV6ZiQpoqhKl+qlfw8sPbdGo0PMQ7N9FxmbmDZq4KoIq+EKFvgBxI7lNKPiK
fVUqFH8DePm7AKD/yzlPLkpig645Qyo2epTGwDIEFQcHKtXl1SJ1CjPmRZO/
ZFqz47/RXtCWOVjcG26yF4UgJ2VV/aGs4gNMNnJClnckoGRTw+DXjNLgmD3z
enV4sI0RPX1FlJRSj+MBwcV8eaxwl9ifKvSphQ+2mu2UlwhBg7GEdgQVErLZ
5rT0HKEjijPn3SEEbnngy4cOIDDmE4j5Tl44rfdRTVsObzGIzeLvz9goRK5Q
z+JGD8Es8quuzTcb7RV7SQr79fHIrOUqRW6wGmjyDyzDy5q+6vY3s60jG6rP
VnafIMxedU/WAzBAD2wbiUzFkbo8vp+EVkJc8qIr24PV3ohxRqEw+Vx4xaAi
AeKnaDlJ4XZwKz82c5xHV8nxgN8/HDZHkRHE3umAX27xfhYpywktugh19sIO
/O1jpBt2vzUrszp2xbjQUurIfXvu1lK0u3Gn8C0mo6Kwa9kVcN8hnrXCwAGW
ITXZwBg6mrBPgeB392Rnjw44shtHYh9VDQGUAAP8Eb26NiLbnYC1Wpnu2x5I
PpjJHnJrMebABMc/Bz8MIpxK9cq02Jp9EGtwYCQ8qc8tdvkgmqeze6nYLW48
/LX6SqgRGDW7G3mIBiJO2cII/ANg0YKySaFuvSFF2DQdaH62dVe++E3A2idE
ku315v1Sjzexc5Mjj81NMgCEAA2nzl5XejZ53SaKGunJH7ZEKdTCmc8AXHY+
pJd/243G1MC2cgGRlAuHfhmVoOOp39eVsiIvoxJfo3/APE3uehf2rwMGXo5z
AWt9Jy9DwzIzmci4f3nQQ8GYyRSqbfqXiVg//KZ3b2sjx0CvkITsh/sdBkPn
IWDkmrkl0EOObNPXlWLn+9fxcu53LPtYIqWqfKd0Dob5EaYDuDQUjy+Beznu
FY25dKrIYxwGjc3yNi7WE2vjPtenUidDVF/9O9LtsAuo2D0m5tCKIuLEZyEJ
2Vj56B/fQ0FNgjT3AkiZxCJzkYVIFM/BPVa1KP1f/sGtADYmcNuZRC2pKWUr
e8M0S6z/p6HNdkMgwUB9an81tmWTG1xAsItKGeW9vPZLY38PEHSPxZ9671Z4
rfKjrZ+sjJFgIB7PcnLTyGL/3CnpdgBgK6lcYkl3bf2/flYJ9hvmV0DpaiCy
TC2dMSnGzBUq45FFUtAF/pF/vhhoyOQwSCObnSGQpmVQvE9YYWimMhgBEu6v
FJO4UKDFzMNMKPgRBBl0qEi85+Zlk0ZIHqM7R+zSqFtQpL3kju1qjXyZwIek
AEpDCE+GH6kT+lqG2LfSe5HkqxqkGcCszgBqxnbk+3deLtTWeieHRTI7he+O
muVtFOv3/7Cgz+WBVC8m0B7bl+M2UMbWGOH4YUkjJYy6uR5Wi0O5cE355CNl
PmJCZrWVpXPyQ9ChRWI3+InSLpABNYXeIBwqSh7Q98gHWbwEq45DiNpFaTD/
PgbJLPDSiM78hi+zSVCTEKtVmIpMwKCHv8DkSZpDSgTCorrMysXlfJOL0t9K
EffETvGQz8knR+wxW2vnXY8j0XCVllH/pb/qAFdNe76HIIXUhJNDFmXbKcCV
zZdEFg5Aa/fg84gnuq7Mk8QP/ieZwnVzRO9l+4ee2vQQik6m3CeuWM3rNaun
vxpy47icQZ9TtMPWHeSo8RFvivI0rcZ5kQeGpwT+7tBA9bDLeQX/OJaZHwbE
x0ei0rs6K9qYVdoEjvxuvAGShbaMb8BhVYoz1rtGSBzJWtk/3VWUQEKx2C66
045DtpU5tTNAyea94CxxCKBSo/pSLlTFOtbVRRu6zNRSuQhd8HjclQQDfYad
XtB+QsFjJbuPxL0boqJ2u6FOwrcpjvO8WPvnlmCLgTkLHPfvPhhP9+qbmtq0
/QIHuKJ5aln8Hyenn1FYeQvzSc9/ElJxtKlVAM5veGEdipdSjZsJkGGWiqeb
HFPrWONcHEkpXdnKk8BYs+U6E0Bky0Mf3KFXeAm2hh6SiSGNl76VZRFRipvA
D3rJEwE8PScLi9ZBTWk+lq6lStqKv6HsZkPSPVh8brLb1KgeTydwux2uxRQW
P+bIkNiv9G11+1swa+2y+tLzScXdAVEAU4Z9GGA0KqyGPmfTpQSOY9Nhv7zp
cF76SSe3wQE0iu6Ox51MDWds7i4OyyKW8+aC6X3UrsyfSEsCjYD75Qea6vrJ
WDYRtYKYQktthaJ5beGY6UUE8ukwXqx0WTESV2KV0M4/6J7jZZL5KrtfikTT
gdmAXGZrBnSmaAWzItWwqzXZXmaH8lbtFiUpGpNrPjNs10pFOgDrEIxVlAKc
o/1Cq0itrD59E488Y+ovYIV3kOvzNfX41X7fKbMklrXvvPFxXCBgMAVPgkEP
+rQKkwc7tVwV8hFKgeL7kONMkmyOGk/CyvBnFAzztoNby55sk3SPSCdUayoq
0sY7bmGRr/fxT/0IlTtwbhXtCMZdBm8eiC3XYpVJaoQ0ebl4daVQeJpoCXt6
En8lAK4OlJCCxS1HPF8MO5PCf3qJ47mU5XWN/SU6P0r2mgoMwsUhSOIUUYOO
34Ztkzkgcs1hx7NJ5WkKLFZ1ogBl+GlkyPhgh4llPS4CfXRBHEskCkBal7g2
sqQKZP5lDYqGT/fJZPTufmo7+X9e2B0EZu+e58HOnPh65q1sfHDE6A6N94sy
g12/ojPZPhks2X8h2CJGTprC0H6GLMFR0e8pGjMzzoqi4bwOq9varAQz8Dg9
QZ+zHVEvs6vuBI/O30oknh9n/vJtHC0nfb5y5TiK4nllpkXI9o4TNe2PpuYh
/1fLahXy1PFgPoXDujqAL1CePJDYFZx1iwVtK7aYdSBX3dviw6Q5mnFvydi/
y8NuptbiT6jYIHCB/1o8snRyjzlLE9MYpKqbeQw5y8JHov/ZCqpKFoyR6uYT
SEMQWMz1GgaWMynSDxjZ9TQi1mi9XmrfZHQMsy03n+C9yBpjfNAX3d4LHK8m
K6uOnWAUabLOxR4l0J/FxOHwlin5g3ie29fO9o2Ag37ellFPdvbcDeM879hS
9DLgAbJXQNmDtsACnY3G5t74pS1s1zpgf2ylqjuKiCTUJ2n9yl9nhk3xvP62
pe8wDVBi/teT2HedbgGksPxEjpoVzvQLe0fhwfta9xaLkhrm+GXEKe9GvKjj
FrvUCOClHUbgojJ+kXWH34DVF7/6iZg3M7oOEhzGEosAKcLzfafWue14hFnH
JJypuP1pUElmPJBJZZXOkWq8Umz9BdCXXoFvPH/j1+UKwcqk0n1GWkA2tAyx
pAodLaJQF9hNVWmJAbPlG0i+4S1Spsin7+JF0SvRuRmaHwI6fYHysmMrOVgI
0vSIRzEVMGceIrhhEbfRLSvrWE9w+hUktzkCjvsSs9gHAbmpIdZZCciBlWxs
qTBal+VmYB/XmZ1j2bRE/uhppInRnsN4FwRPpsSxlellSINo094/B1JOUTmx
IFDfsI21/ZG8v733SMhlSrlMOkoqMKYAXN/FIIsFX1r6P1Dhm2ZdJljs+zN+
5Ywx4Igl+ImBgDK1iCOj42L3OjxY97cQg573Lm1yz8pDLTbsjNHdPazXWjxV
/LVjbZRqyFMCzudxkQf6orWySMn3lFuJ9pIp/Pd8rQDDqXJVsCxmc/q640EL
8Ev9JPzPcXYI3phyijAbwaRSKt36We5hWK3rDbS6Bf/lDk2pP0X9K9FhbQTU
QQh8IKSYsLD49S93HUf9A48pm/Xobvabd/UHwi1IIaMIQ1Lt/278jMlHd4eY
5loManSy2BYOcLxP2zktm5Qqai2/QcP0+LsTnoAFQkhX3T6N0WYKHtj0dxmx
ITIHnRV7MzZ8k0CLlAZpbRODaAwPUPFIJZyn72G8gQHZ/PQIjKzcjeBxLqPK
sNfCQIcX1nc3oGWtJza28CI6z0SIBSBM1Fg2A7J1HwAI3V6sPZLmVMS6U166
ptmCiVkX0wsmSwG+WqSS4OGVu+DI3uzDnox7aKDz/IjnjNLcrxtvjHHPq2AJ
4Bptcdaeydmy6osAZZ84lm+qawnxzMxt+IxYCgU1vIntpYQQhZDyq7x2Ohqq
cxjUtVxF5d0uc0xr9KavJRA65IwL775VCLpi53CiIaNL+3PSu0C8HM+JPU7I
bw4CYVADR65N+qTNhdzdLFRZj3hm57jaVIG1neUK9xTQ0bx55EAav8GVsLQq
NeSU9nqrUGXw8P0wkNqJEE+sb2eZv+bhkt7WEyioNTvNMba1ZTpwudFhKNvZ
a1GHMdFDEsTpR79NRRKsL5n0JIxaUq0z+vO4OT/vPfQCNstT2L8x8dvl4PA2
Rq8aMYlaDo1SVJbcnaWcLANAT6yBTOUg8Sm9FWqxK1AQ6i5jz38Gs3SqOTTJ
T8E089+UFZJmoXkYjJApA8efLNljs7jfxZhv9IS9KHFH/bH8se1CDRJG034y
MLA35t/ckro7UDmGATAHRrHiuAhhqd5OLrIIA6zKSlpQRqwsh6MkpVZhsU+j
nwrdr8RaLvTulNmScZBbonZ2KX13HmeBn5e0fjeK72iKUTUh2clfvdZ0TAxi
p8dT6qFYB6JG3GJoVb24TNyf7c/6B8aQaKhBo2qWB/WHtrlLGigYzDHyLI4b
xw9sDiAXcuy2oKvxJbJ0LJ1lMCkAeJAuMHoROWQpmK8VzTIRzvSqIdg+6hZi
V+gC46NNhMeV9nCuRmleQBh1mH1C10k+l7bEMWXy5zR+CNuoJz2KHELnbhwJ
RsSPgr1HoVmz+8dPJedyP1GR5p6i5oBObkZ8HntumdCKlZ3yT1ndNlSJZAGy
5UQtkt8qOlQ8kCeC5h9858hKYOHDNN7SoBT4F6NObvqCx/WtA0lWOMhrMerA
SMwzlvSUBh59C9Kg+TCcJK8PBPqn9Blb6cG/QUb3XA9/mPHhgtL0UoRwRSyv
o+Hao+t2FRmHqwxr4h0ZeCU/N/iE6Djs2wLt12zbUbHA6YJJdJeuP89V9PND
F12oUjgW0AeJsa8xGnfBGBdqpNkT7f7KaEIm1nH84nC1pRdrpI/uoGHin2UD
Q3btt8GiXk5wHPv8mGhCoeFrj9oQyDYHhTb1TGE0xHQH0d6Gro3RNzFYFAhV
nXAFhNJiGExXaEr+rrBpNCqMTXwuCa/I0+rJ2TjaIaRRmHpLHtFsqxA95utl
soRk7H4RownmP2rikf1qL5POpf5fkxbtNC+5Gv6hWl9ZGTaOEKEgpPAXco18
FQYNH66T4oauIgVGi6oet9UGxGUm+2N6qTBOWPzZWw9CBgPkpOvADx4qTOZG
uZO1j202BGwcRqQ/T8/aH07ggvnkYKl5JUIRsgdLoU/GavJ+fCUnNoq73HZD
DyobCJHAByUUWVN9GdhcIGQgPNi2Z7eVr0jEYgW+ANnGjScO8nYMZDLBV2zx
ILwuG0KGJx9/B7W3lTzEi+ESZ7Jc1kezCrQM1dAsAzFVzNLQhABsMdRsFux7
qSVyvqqtJyptvn0hiRAfgn4y7vPjGQ6YRcFeZBwuHXmTYEvOj6NhR1PUhqya
ZxWUKl714jnYWBC8I/cdMpOtREKczwD0E0mmSyeirQM4Pk8AJy7Dvx73IkH+
pnJ37UENc/c0HSGjqfoFj6huBFCKwUK9JH8Iezks9T3rLPiS9ejBGrHz7Jm4
V3b6Q1pcc0eL8VZZ42QOEDzPfhqbikIDC/wofDuc+QDdQYtU+UQsubq6XUBY
kCClQos3y0PvQpACX++FmYVgfv/oV1seOTcFQ1otD8x5P10E3ZQrcWxMm4AC
Qlc27hpYRnb85ibwtsBwqWsRGjJz3X/IrS8gXk+L8RIMetODLiUgk9STuK/0
91Flw4gmJUtnsT97tmrHFOZpl408en9lY8bg3J81YO1wripm1DQvwEr3DepU
lK5OuyxSZtzLetpi6CGmALMfyKPuxhgQ5sd/IDqYrrWhHN9c9JEUreNpLqpx
4upyyFhrSPo9akG2rrwfks5eE23eKrLh/95YqipX4E4K/4AfOI2qGEU1SX7B
NVE4IsooQoJ4JnA69btJRQLw0PvcAiXIG3xO7UvX2dFPXGXAgF15vO7D9l5P
4p27J0QaqzRCyzEEWM1pvztJt/oQSC6kHNtTlXOBSejbk46kbv87Zq21Y6do
hZ+R5RcxyxrETtkVgp77UpnjLMfBDxQT9/R6Txw3IkkhWX1JmUuGE6JED2TP
D2X5B/FA/Cr+N6tnK7MG6julDpzlvHeLDkgQZXu7rXswDwAG20O1qa6upJMo
ZL2nF+gwCk1kFvbxFDOy6epJc+zyN4qLo7z5c7gy+UWn+iYhMlsw/7RrtLmZ
ZePgYsLUHxhR/O1/P8PmDls+pPp2ZTb9haZunkaz4gEqKABApwZejWBkrgcO
1JO6MDWJW9DZJzSwQTSSgtFbgI+0qKSTYsVRP/3O4ELeCwhZb3e+ptaqYTTq
TdeZFmsWQdG1zD5G4vWZJd0yEWhwbZ84PLbrq5wtCdu0K6uZgQ1rMAz8vc27
VpWLyvSO1eNx7qEztHt83DG2XZhqoP3QTby/10NYrlEXsE8qn+UJu4X1CuR3
a4SPY9k9unoAGBWsQFEd+QlwRUbirIsX9C6+q5LNaFm01wBDON32dMjp+iEx
EC+iFnydKoFI3DW1NTyCdfQr363TX0uvQLeESXpCcOs11aRWNtZZBfOkyLSy
pv0hd51IcmZDoyKMU2LssOeh5VJzWGeRhKwAknv0/49ssJ2wMUvAjnD3Wovf
T/ncNfqceIm8d5/vFa+IhUe+l0OXpXxSLq9fKThc7OYRHX8tzcKMkdZmpk39
Yxl6XkkMP0VUZXIOafqgFujlW9MYFHVqB24ZG+cb1wnfVd7jqz/EuhylCIC4
WGlFLQrcoMtX98vo2iOdHl2bGkGiRpqR5pfya7tyY/cYfT0+HvPaHZ0tjbhQ
uAKg5Wglz6bJHkdxv7bs6gA8dqDfqI2kNNTI2YyXu6WmcSg489XDL5/EJK0H
ffdJO3RBRSy4moSNxRJia3zT3gUlU6Im24PIZzQ6JaV415uN65+YINKda8qZ
1Qkx3FHb6dIXB9+/7RQPMASujn3FLqPp4yoCVCiiRdqAnqi3uRnyXIUUtqlc
SfUStGID7/AI/5pWRNEF2Zo6D+94NbMOcA0LP/VD4/ngd8f9iHt9LJLDkuqN
VDszwiwBiSEIoh9lYqLSbc/j4ChdHxY88j5yniLsQ8esnZXBKfmjOE/yJp6a
khgL304FJEXFute7l+74K5FhPC1MYG/1L3QP5b/mRS0T1R1jsxZWl+CPLokh
m96hKI20I8kraGTHFkfxD4KwdwKtepFsI6pEgyiGXlR7fj+YsCF/ZBLF5lfy
lZuPfZgDRKNU8D4yDOqH0Nk3pfWI8DHzO3tD8X1E+JH+yV/t93vxMcuClxso
K2llCmIX0P7B9XjyzSKxT1a1twvBnF3LHFJen1MEqsUdCJdoAzxWLno62g5c
veYBPETJSGhLZT/M/Gc6nkrpuq1rnlltPoqcfek9Ku1HFmi+8iCP18bp3n8e
nmS0PyUyTcvQGKfM/+8igVTqLzURTDUX2Dsv63VMeN9fkt+ead9SDiz8jCNo
M0rzsZsjPKf2tGO41IlB+86aSj1jGvpcThQ9GwUnLC36DCbxLGX86fL9gB4s
qfVrMkJN2STVxjBCjSYr8J0sZV3KulRMFMFhaVnUD6RIHDhuHaKXrtAX6cuN
uod47qqnmozFwin4ZJopbxEVnj6slF6p30HyPPbYsEV/oFjB/xg/ShMC/5KA
4/vuV/8FCKqUUbBUMrU6Od+RJ3SSy8zvvrpb+mn/sIy87I+ufWsEUK2b8lzy
SnpI6LwzagxRywKwEfvN5JO7xeqWfJ0070AOZYB0tatVhSz170gI/nrXkrBL
rMXkixpyFt2hXrvJrm3ka+8I8nNz+KcSakaIzW3TdKJCJlaT454HLBHEp6Wj
FPNCFn4vLgoQYzEzh/RDzDLWEImMinDpGjA51js+TU5NvfaI4ZKgLFlmH9OA
9iLdHlzSqIDGX/gDvI8cSUXwWRwzr060JruC84LCwx9e1rBf1CLyf7oc5E/Y
xLZ6VxLGhDI4bBmcnWLeioTQBXdYd3votVaShkQqMQBaFLbl7UjPloDwEcLS
BAwJXBorqIJpi8KEqPiwRG3h89+qK4BENJtcCFxrkuHqSR9xz0AkBz+6JbuY
ZTU/MurDUl/D41pAMZRoGqLWWoqRmyIpIPbJE1olACH4T0lyIYfwU1UpLtEB
eAJyfSpQJp5ZlBSD7avLSXqYOgnkJH1U1nLTFDtt8kCiWdQ2b7wyd78SLjFU
SgXq0BtIA3XPpLMrQEHIvmuUlq0sNtPnYatJJglsnRxukMPnuj8PWGfzpdKz
XJ1hZPcY5BuGKeVDxoRL/lwOTELUGBrhTb5v2gTMT2cpJUy0Tx/lpYGf9FIu
k3LBz8AgIC9RPxiX+mq/CSeKKw1VTBVEfkQUMPFqwgDat1HnHLkNhS/zI4ip
MLdV5vnnXhTvG4px5SxJ0xDl5tw8f+5SwaeVhp0K5tOxWMDTCNJzL1+vgXhS
AyNG6e7xVrKu+tZ6LtVzd040Op+efugKAlwpeVTfDGoyWXoLP/pMaQSp6N7e
wFXhoya2rw5PJ6M2V7GTt73F7T2AI5Ao/wpn9t3SRo0wLWg57kYC3vywyGDp
owpz4AAGE7O92x+BbakEbCCwIvk2lZ+hjYIBuD/cC7fSGi/gQdYtv45giX2q
BPBIXeEL7kmeNoXt5fbnMxfkSi6V+scCEttJqv2Ei6VdGUNm1aJyw21TRbFr
/kXyAvvI6jLpBDflVvrE2BaK9P+rbT85yQQKABJcqRQNhBgaSOd26PoTM1VT
QfjZTPdlCV2rw+piFdoihRzaciEZ6SvOXJfFWL6gbpPA6I5fUom7PulaAFDc
V/BEZ0Yrod7yh3lGH0JN77eUn5b2fftHECwP/Cm57NVTWTw/1ylXQG3mbDpp
4xgT0qyF4jvQRiBA8E+O5EeiFdNhgm9CDCEgj/8c6+Bxrv3jgxWKS58nJxyP
J/CxWSysE/ULgwyQuHXRulNSudNO5nL2deB3/IgXLurih772qpR8xwixNTfx
l0MWWYQnEvW1V51HvNlIm+LvUkHQapEb9BdFl6JZM3HrIIUH55A0WUCrvFl0
ViDDFaiijlwHmz5vzrRNGXDOe5TJkpLOJmk9b6Vr7XuitMHPmCjlTvCd3MbF
lqkohADmi79qA399pKtIodXI6o7ztsKDE8EFJYu1BRc2indDPNYj7n3O2dtk
y9wDGJPnEBv6N6++zLMuHMd8tyIWAFK3zPusBt7eolE8heBu3PUlBXlypSzq
d4UBibmubikHBxkVLwlFsS9dog9/cV8CH/TSrxDq9aXqA1kklEtmI03eEBP4
ZxDY5T4M/B1txhieCBAw+xgzUJhkpEurtUKKNPk4Fk/QYI0HP77YJq7YhRfW
0jzPZrLEGsRo19NfcYUJ9txD1cv6cYlJXVCt4SYoQlaJQrBGJq4XUSbCNTNR
QhHKkBAztwhGJyVmWj5O2g8uyO0jVkg7/U1VRJ+1l+f96Jd5vZv74WABtUd3
VmNBysiH7MUj+/5zo8o5eI5PfOT7SG8XSO5Z5A0MPfPzRwRWOG86wb+KpH/0
mXc5jojy2SGZDeaeZlkOdJPjVz02I5Z2GifPPKfs7aaLEdojzESgjQt7ah+L
9Fx1n5y37YrYi3YvSELGilrxXp56mfd59B1QIYysWXMWXM3kC32vegI9C1W8
Da8wTODoM48k9n+wCdtyM3HIjEeruxsdsjxhy2ey7aqXPkyniYhga9xOjzGU
5APPRQMzfQlTFyTj1EAhhdJMbzv7RI6dCbv7ds5Y+nXq9riOXdpNl/6EpRen
CqTDQTpJmPF3MOj5ab8/vdwY6yQ2HC+NXr8QoC4FTbvtxVnUc5DHrmiifw2Q
mpTOhy75LtS4iMHLJW3aX2Vgs1plWde/Ws9pQklckOGLf977wOLbARZp/SWf
xmdbXf6Lo63Nn4ykR54sYrvyzc2KvDQm3XbWyv8Um2L1a+BV87RrbksHqU4P
bigY84dm654sBkajTJg15fbOgGxyqf2q0xZ6G99q0J7mwAUiHNfXyoNfrfTk
K+31EgC9LzAnb796s+tKXdjn7QWyMbGnsxqnMNZgKoybLWAIZDCahTuhYCCR
gfknxskvCMbDNReWihHAA2vY7HPGsdG4/o+iEXL4cTEcQB4pWAlT4kR4CdcC
u9bvw+Sf2AHhKv4u6TOoa8VF62w2mLo9/Um9AcWWJzODZ94D/st4V/u3Xfyp
VGXBvRGkos0aZM8ehrdnihniAOTtZGUiRqATjpfNp3Fi6oIf2MjmDDeUH7qS
Zzzm1FCmk1O2a1pQ/4kfPYOwO0qV0nvjLna2glW+g1LujweistgYyOE8/1OI
sA7HPymczbU8E+8pcRdJJP5RBQIee7MG/Y2LKXav4nbAq4qiDNI98APWPXQC
cE+4omeHYeqmW6F3t01Z0u3JS/JwX3HNlmiDmTO8JsFWW5/GSuJRRgKyt6Yw
mnSAo4klEcfaS6B0bAmKgUhLJMrdlQ5RtSd7y8F5przVNDHmnEUmnWyhnT3Z
oRCcr8L1i+Fsca2t5iCxzw+I/cbo3kDr64N2EUvQl8qnSTyN23+Y4cVrZzD4
8P0sAU4F/+uq/tocFgxyv4Lw3uoo5da0vRtGYjaZ/7cFVbG3Vg8h9SEPFuwT
JvVbKY5G/+kZtO7ufYw/jA/MS6c57tS9hOfkd1aWX49EJoFg2Yy1i4tEcJNf
w5yQhrVMuJlQoJPdpkH/HtLmnEdgX5upU2ApYgk7fB7Khc6ycY7ngwsTWXp7
2rsnN3N2cYrqfUURqHuLNGYU8r81361SWmGcPak+oYcfLlkYW9IGBnBhvFGx
rR2c/1Pe/4l9/Z//jZRmSNFneVIW7wSC7cox0HKZsjjebY4bhilo9nQH+jiJ
T59UlvBJjW8ILEAsDdy+6bwnDA0JUGsyWaBzaQirNlLLCLIuZ3Zp/mDWwH3g
v5y1NsbaJnuSTCOof+X3Jwct+KFhtaYCx8CRVNR/mTdq+09qBayvdp/lJWlU
Od2i6zl5Fco+ZolVSELeIMFHi8A4Z5uZyVeoUrlFC8qT4bP89CJz8y+XkJZJ
NuqE9OwGvIhUQbmQC8olC2TfNzFsDpGKVYA5JJ5l3T0vHKdNEkc6OrKkthoy
G03cSq+FJ1wtI06HNiRnWjbM/S/ElFwy/yxslMSA0lNXrzbsvWYfRNrz+xbZ
sh6M03/VxfqupKwfv7f0qO2ItyWcQKG9Y/aSMY/jaDILFLAKBwNlBxTZwyjS
DicUEn/V9+XSk1RYvO1q0ZoJSAAgk1Dd8ZISxcAdswP/RKpYHINplQ5KnpTp
Ytru4Mf1bcMUM0hgDvg/PqCliVntogMAxTeM4BPpZ33FEIXwjiKm5aN4Kl22
ZesHtSz0+Fv3UlV8/4aCyA/nXcyzJ8wP3nFUhwZ/IEdQtMA6S2r7Pjscv4w6
9qVcZVWhhBGdKQOkN7cIFdOOHgWYbvEWIA2sKMqG408pe0boh0KLqL3+Suvj
XN4mROVd84T2SU4dEfQRd8iyRq+A5kZIp/tcGqOuXFnIPk7TOTto37G1t6uJ
DBXuk1l2Wlqu6p2Q1p4wFpWfnH1C1+UztfVWhAi98LOmLIEhFaNU4c4IY86p
RcD4CwHNrYBKZGCxRcjdGgOjeHKzG4Ja4AQTYh1TvIuoQnJlEQuD93kE1DAW
r3+FyOEVlP9Yt2r7WOQItvtO6VIrzhVyAXeimrYSnsZTQCYc7cxZkmA0/L/4
KZL53g7b6byQi7BhQWJHLY4FG3L+UKtll28gCqtOUiDr18nmGNw2bSCgWmhz
VvX96qvx/Ydi+rfoG4XCKU58oljEWtEo+rfUfLOOdYuD3R7SyhnD8pxxHIi1
mXPos5TlF9v8GZX8qGDErmvuzyIQg/YK2wpOFxdPsyFZXAkyVKV5ir/81lyu
4/RxqjTprwWBnXun5st8+f02yNF/jKzeIdNR2WYhtrkWmRxcTGmYTiiHgmKH
XLCb4prEW0Zv3sqi/L6VeBXqhJubA1p0LbKSkguasV5R6EZeFMwNKeiTnIdM
fQpRexkvO6kjF04NFkgvB5NrN0Zl4fRq9G5gbwi5z0y3cPiEQP4Ju/X1Nwjg
h9fahPhdi+FhmwLiIGQvQnhGSmbPIDaXBzfH5zIlrjA1l6WDHaNBctXT8fex
XVUXpLAMnJED3lH1fWfpdI3b7VN1+OC9fHnljnsTUw9z1Q7CtmNPaXq5uWic
c7TforaeDS+QEAmzbJSRuKMx5hlJ02EgVEY2fkPaYAldWbf5khavrqDSeCPY
OVcGc5jmjZB7QMvx6WVitI8ldaLFmDP9dPmP8cF7CgHW1Hxl8Ct0hj/R95U0
93odSNKpG3Rk9Q9K0w+n/DnLbJKpRVX/3HrRtUcpcRanC6XXGvajeGJDJdlp
MlzRnSmMW5ak5ZSihni7dt8g4Ov5NjQUJMu1IbQvTbvasvMFWW6HAqEkanpk
MOPrOGPHxQfo1wOfmrYkGivvXZNAz18NN9QETOVYtAk/FsELYQndHsO7rWiU
pbpUxJYFGP209SOomgOY8RHHzEf+4Yivk3QkR09zXJiyw8V4Tb3zlMRWVlT7
dvsKMTLzY/WVxHIfZ0Sg9bk4q4RP+xu5+oQgfNDQ3IzS4YgMPm2Ml+xDxUF1
AswGjVWEZ6o9HPcrFWkBh3t/xvTF+UC36ipLofhxlQv08GdTtvVpvrGgs67i
PgeWWm4p3K7pi6FteCBubUM7+xuVeFZ5vqr5uMjZYpiLN0OrFA2y9L3gDAvF
RxKAmwO9g9EAT84zGMABTF5I88Fm4Lo7p3doVJLaf7wwfytiBYkwwwO3guiP
L2lUj85LYUMVBh+TY7yEP8leNu1t3SZIiA8CX1w4SnFkAqjfpjfg4XApo+tG
20nqBvqquhAMYWiWTmsxhRDyCX5aROGZRkbGst6AyqIxUiLlkA2/ngCvugte
i3rKNgiy5jR40/vdAM8z5id2Qiz/JZL62EixFw4xhGOVt/Ejip3JkgtxhB7p
e/KuqHI8hhKg3e1x+Fn6KlB6iYdZCjXY80js674RXPZwtZEARqNRuZTJtOWo
elWGou0/xLj9YqAbvzLgtb/37+UFhGk8l79D9JvgLbn/yjGUq3xALRP//fv4
Fnzz6YWXlyAg4niYsPVcwsKPFmoJWie5ibrd8m5yU+JF/MKWfMMQwK24tTkK
88Rfe3ipyVhKRqxgK67MgGiTFMjXZL5hcr4P1diDnVV/qQ8r0q1Ru9wZD0GC
MJrOfLqC1hiRtSg7jkbUficueRXpJ2PbrxKmf+F4rZ9H6C7gIWSnOdWiyyNZ
JgogtAtIVhrZe0IjXIakNwSh4RGG14VLuv1PpMvZY2fn+WbcR9YX3r7G82Al
3bF8zuMx6pN1rpZTFC2Af7e2GHNHasAMqAC5FMOgXj6zqlQ8IQBtxtRGXj3M
NHDZ0LNPptjjtrh0QfnD8sftmmFmSftRQob8slJfr7bfEuf5vCsSntU8jEn/
9a32qZfRS42nt619q6KPV6a2j6s9qpHVUWIb1K+PuetbywMZ9H6hD4oxJH5n
Sx+Wy4WWe5hDEyiSTpyNKlytPvMmnmU9Eu7A8giRQhK3v27nuhCm/8MKPM0C
pOF9c7isxwDyCRlkypYAzE7S/4bCKsAfsTG2JajshhGocH5LKd6RnNGtqtEm
zLuiUg2rCvm7+fQPttuAiYe/bJVl1dBMZQ+b1LO6SXhaWtm1b2lVHHiMJDI3
D7dO19M15BT6BIcpDwtnG1zuWc2ttszX9tbtTaK3+oUoJ8hRkBe7F7pIp22b
1KKOyrkStfJeLW++4acpXWZYVz373zyIDHqfmS5cAic2Et/w5k4s9WyYNp4z
h441F+NOIozQQuCfRZy/4nPy+h/sV7yl01Y4WFKJqbhNJ0CL/numUN+6lAbe
oHPfbvoqIGTnReovbLWWhgMezfGqZq/a0oGD0Apl56rZF0p5BPwfIBw8k3yj
/RIw+fZ4nKhhUup96vI79xY3wycNHd7q/r3UYDuBRHwSF7vJpuDZEREZpvce
22RJI6QRh0ZlOVEx2yMwZ60f+I0gtMJ7yU+/+mI7fsTjBob+mSAgOEeZ9xjo
3BWYYU4cEhyEYKs2W9MuE56D+ZOBEpB12crGqc6Ua9NZpIgX9nWqgs5Zz/yU
c1u+d5pcMbtDYjVj2uAHn5uEz4CD9M+frNa0XIZ2eBPP7kHgWKmcaWGNX9mf
orzJKthSbIziJJosQwm/FW12HSC0Eht1NCYXdR/r5l0iJM1d9ozE+WV4i8Hv
jjU53YKyKzQoHy9pExOE5wyW3wKmI9EAEoeX+iM4tWpXziEYLhwNNq51/x+W
4MdGuy/g4qzDYq5s2buCsrnNJzMip9TI82FuqMeFQUZDR+zn3c7QxNObuQYe
dX6u6btrh5zXkixxCNWB5cIc87jOy/F+6BYcYfjeFx5NimQ+ws2HzqV6SYX2
qyO0wiUddikwOYOajNUfBGwhfQ5Ekr9293m5l2GekxwwT0N/gkMdcClRHDtu
BULp9DnzSLcvBun0Da/5Uir6/PiIHRUZ6ChHrM3++MxuVc2tPcNilTBGaLI9
U4aQfT32LuFf/ssQH6cJCQlGzkJiyftGJzTep3rC/OEm+uid11bJewuaWhTK
WmaXHOJcFTAf/ISLVtBxruSbiC+keSRjFpNsSleyHhYBezWcKVCgMzrA5nLT
rC1beO+xcWugNVuUsUXV42hoCKS7lKGGzjTMNYIWTYZN0I9NrxUddCCN03Y5
8S2kLPVruJqR0YEkYdxOobg1frUTe56pAavGO3T3pxpLVG9xiNXK2T4ZEoAl
67i2ASH0+QKvSKmJSnk35Y/uiHzbMmWjfZvXMvaeQQi0BpzAd6EWCqeWnjov
W8NMKk+b3+5cREzOpoQqLOnXXiH0axY2ioA57I8T1OJOpUbCyyKuUyCp0EDb
MPy/nUdFz4GE1w+LSxuY5Fl/NpAlByMQxHATXyRehPmQBi5ngtB7rGxSDIXh
kk2GtPTM+jR1Y5n/c7RyA5jYjFHHYdWuy5CuNpvGT4eoipwoUmJSE7DaFgHC
VaazGJRf4xH4khJaTd29WaTTeXhrP1Xaue0JR+4humd2nd/d3kObBEREsnP/
iWRyzloG2Tt8u+L6PiiinFnap+420WUk/FI1kz59uoG5ohmXbM4ROj+myC3G
M6ujI7Waz5xeEWfghVCefjgtc764b0rO4j30Klk+LDb6+PUlmx4EZSs0jEhu
w2uL7TPD/C7U+eijF+WTktrEyw1CU7i1kaF6yvIe3Gy6GKcJZ1IiXWhzpvqR
yB7mdgq/cyhoYVYcTRcpsOARle2nyF4o5faEDIS5fp+IKCI37S7BlmvZHCno
jnFhb14p8DSF68nMkkfnEIwsraWI1bAg6/P+sxtOem3Lh3uo0az2ymt+FyQf
yhL7/7flO4F8UhGGxyy9Jw2b5kn2HWgGzL+3gx6hwWVe9Orh/ri5Gur37Kuv
SAReQQxwnoREZJQtmQXk+Cr0SUqua/ExjklKzMSK3zAqWB2sYjpMkGrKAK80
LRyUS3nlJi7uCYL1zlCUfStl/CRR17sl+UyLBACi7G41veqtkE2DvApqN6WQ
UnKPAp7z5wzGOAwe3qivW3daYDg656s2zW6KC2NcwHTn6JTvjKkgTV6v7TPm
zx2wrxTAq1o2c1gCISpqlr9A6iuwKj1CbO/6lEOZyXQOGRFFM9LSRNW7KNYB
yqqYAUDEfXrsrJ5r+JNZ5UqCieRZ9a8xXq2WA8IdO0OsFEj8tZLFzJHCWl1d
wobNH1/E9PiIJEbC+lxXi6nuVM7NyW2qVG9T5RneOF7q9Br48u/co6x66K0q
SMMjNnnKqvye0Sh6a4d5B/h4F3qmV+lU8FMhDWLk1qzE3YJQMUMXNa3iZ34i
JLETwOLxFiUlVwMR09M7H/YnqQf0oJe7lYlpUxsBu+q7RjClta+yihC8//uf
PRbtGx3yOZWfDP0PM6xCFkixDSqALLAtR6dHkZrPA0BbYy+OpWq3rj22IRWE
bI5BcmUagmQhlhHbeariQjiyhyyw8tM1jL4LjN/CeLPnubt1mR/MeqGMbNti
DdS/iJ1FgjO1wxJmlsqMn76+VH32O76OyWdrRn+9O8QvjeVG8ijGbCluMCeM
kp1AQgrvp+tBe/kx/7Iozel8LnMKYShBVaQI4txR7pQ2jyGswtP3mEcThA/I
5oT9efqQGIgrMpBBJnKw6KWTQYIhkjJjRK2S8qYG/5nKDwVijzSOkQwoobVO
ovWA942RBy0+weA2A2N1uHde0MGWij7Im6iHCkuv0MsuE9x7dxbSoqgN2jDR
JflIw9xDOEao2d66rBg+pDJTR/an7NZrY9fxI8WYpZV1Tu91I6eYfZZe7mEq
aYooprTE/bIFaWVyC3zp3xWtg2Tn+dsGclfsIWg3np+o0PAu5cSAoZqWdsYa
KkDGRIjWdH298MY4tSRBKhTilhVvkzqksRxmU8Wqm08YbcMkBDuXMH7MkA1O
Y1MUWK3KXChT/I1fVUhWwKeshZ6K6qyARpVBzEW0oUYDVKbHhx4bMz4GKHHa
rwWMcCIaudvz2rSR0FNEfFtWYlyB1ed/M3VeIlY0mKtzwpuaewPAecomNdS0
EvXggz9lHptkCLHDIW+aLpmSp2zQY2IpgXIPty9t4v38cRY3N/EWsl4nGq6H
Kti/yHnh7V3/5w+XkkpIizabrmp89M3FiZVdwBFflvwHTurpifFYlWC7FomL
A62lp8GjmuWHLghVzC8gJayPUk3YMJN3yqClPTCBwMzVz/JGnpkPjP4ftVX+
1gci+KjGcLLUp8+3QlCKzN6PgFkEPjq00azFCCyQE+V0KRIIh96uIlhmCpQE
vbm159gc+GVzrk68Aj0hToxEpUIbzPJ7ccPXBuxcUlg5iB5SLyP+KSXIl9fK
HgWoxTIDA990aJtWh8+jeruzLJxet00EOOH/YGW9XfKgFXK+dO+pUg6wIyOj
C6KOJnlrwUmgZ/iYCmM798Dbl5iDHGty9o2VR8YJVgbpsVlkreDItWaumyDS
kSCmgh7KEeXw/RYSOBGqgVeCMvDvgM7KnbCSGV7djizlwGWwbJ8MZMCkhpTX
Ke535mWFHWP55B4ODSKh3SdJ/ijThyfwAutj7cvC89wnDaXXDh566hsffkE0
RGjdNdd46QMK5RBAVwM1+CPV+xbg08u0UyH7ebM1QVUUopvGNNSwT2W0BdrJ
YO0OIqTcK/eszg5xwdf1lCnJy5VCwwtqFbhz0BjG0OXtJ+hvDeoTzkAXpHxp
ICV4GuaVM7ysP8RZXokKQOctdq1uRTFqdmlCZrRx9c35aUlEGyuWXTJRiQN+
R64/ccFK7OzXRCYzaBz0sKdJPCI7Zo0wuVhIkOu/gLd6j20K1y8mp4wgcGJp
crrJBNTPy2IpZJH59srBkbix6VpGhWmXChvZzppg/rsWFVbLPnF2Ih4nZ5Zc
XrIRvrFesfUBl5vqSG+B/3spYnff2tCRwH8PS2sOH0Ssw8jOIl5p5GC7EqiU
fgR3fmykrQw4dxzHqmufecXHrc4S07Vk3qSZZFdpIr0R2Yt0fXOB7ZvwgJg0
zyBzkIvQ4oXOVVY+wrgDJza0LrjZYilZSgZozYB2iO+GZtrok0vFQGtq2KLp
iMrDSj5v4Y0M+/8bZKsrYtdku8hhJ/wMTSz7oXJt0EZb3D7BtF8ruen/Nu4m
iYs9EzR7gRhfAYruPt/83eMWxBewilg2r3v2aqdAVfpJKCJ7FyXUJCtROTW9
UkoDz7oJx2OHd+N2uLO/yStaDf31RNuBmrGEtDc7OTmr2h2Sb3WP2kAlcuqx
Nm4b0WELuARABZ3C2E1VaRgGTditqBOOvLfyxg+nk7KJTpzJP2PCcGnPZDwx
OGokvRD9ESm1TrzMibx5xBr9/Ym2U0GE1pmVl78u6R65zoZgCOFVvY4cGlfX
pHZlaK00l5DYMmlJZz77kiZHCNlX2uZqT0MY2FkKsG0zGoEFfdNiPcIA8GRO
ityJPLDJgRUh70bbjMsho3H39Np2AifO6/0TIZC6ZQAzvL7odLO012O0cYhb
nyBxy1IOXxTLc/aTmYdXiB0j37TKbtIgIgiFrjBNvS/rbwAlMMr/RPv8jBAJ
2n6aFuMMsBsGuuvSY0fxTOqtBg77KRHJ2FEMLfjlBQA38dtSKCfani4D9tDb
mIwUsJfGsstsSeabzG4BA+NZefdC2CQojVGGEijCgSyyrSl1sJfktXK2QF1u
bpZHCwDgqT8mLe+naDixhQhDFRvQG2yswmp2VJg0gftee2GfJLwIRjogtsbc
NIy91kyGmEckVb48pdasaDRe6EIC77FLYwEbqU3YKl4aP238vdXrsaO67mnH
el2z6fpOX0xV/tUms5Gb2mp7yQmS9oG6ZkV968ruolhBv4eXEe3QBPjSiD66
QFKgEqM/looUSR0E+tG4pk6mqf6+HPOd0RcaLe49j9f24rzOxvIFJPX/VCt6
N6MKuOkGYfhXZ1Wq8Pg9W3kHsFxCFfEBbYXW8TFGbSlWmZa0tUSgSpRmMzHU
r5OVnpjYTXwtidH2iS5eA2M7ASlB9EubGUlcK1ZVAk4PJRoqrAyr2Z61KMhX
u6HSxefiBbVnv2bkSAUZfWBqkjjwwgfIo/I9y7AR9OlulO+jflkCgiWwrTFs
YeHA93ycjXtMbDHa7Px7zh/ypKQAJuTeqV1BV50wADpW9wqUiUxnoI4eYAU8
d5yoM2rqAAXyUCRhuE+JqRLi8yJf1tuTnADpmIj8WvLvUW5xqRgc9+WjOR9/
pce/qHL94NVMkbECvp+NQIi169hff6Qn3ihK3zfT2mWG7BQ5S5hP+npJdAvd
rAIbfBdVHNIi/6TASIvZ9OgkjMT6serBvOwWOJuVrRofNDkDwZA1wKk61DVt
Hpj+QgsHUoWaVyUNwyeu2fzrZCSuhu9BzWq8VZakHxdfLlTBCNX7p1hUTq9d
xsG0+nbUyDlABa/J+7N+puJ0ajKkplPFLVE1koH7Asz7DyILfoevacXg2xu6
zIhu1arPomi2ab5rtLsYjo7Mhivjxd0slvtcS5TQ/kpjVgjzFwlVwehfqJZA
F5HE0HoB+EPXrjpv4dWGw1+Fu2qo0lI9VbAdaVrpt89vef1VR4IfzL583YgH
II5ckF+s2diJelgIUKtWUiYAdI2rEdUJbys4lgo1nFHbtOKBYyK7B9zAtrsv
IKhknqh1G0MXrJXW2sJ73A0SJObks9X848BzofA7sixm6gpx3zbmAGqL3aIm
4I+wOLim1PC+m5k2HyMBtGubM/Poi1uz1Aq0dgRJbXzFPiXemfuX6G9a1Kb8
c6ufggj4N3P4kpSUcG5IM9ovtoxDmsSD7P6K6Gcs9cp4MDzbuPZMkMXX0Hcg
HHSnbrm7TfDVNT7bkkp8dtHmlyQdzbUM9/mk2/719pJvByvMfrOR8s1DvMkF
2KPpLsjGxMnktvvi1ger0AoIGm0fCsASpKG+1AIWfbNDL0xF7XpPnZjnYP2A
E90GMVUALGm2xIm5ZZ5RyXMh10NO+9WxMTZvCjm2Hx4cPIqUv1hh7GEWbPu3
dpjwERjnVRWNtd+FXOObpwc1VqtQSZaxw4dQFRG41KPzr6Ggw/YtcczX23Qz
1tjgaK/3Uiw2Sp+QkPZxLZINWVvCT6s2zGUBCJHNYDTZrqUqMZ4ef3C6tt4d
eKeWt+kw2rD4i/xK/GW2qzMxQiIJA+MHeMO4BMNdzVAs+ms429a/1FAqsEvm
EMLUOrG3/zKpsXfRMpTQSzL8EZZaNjod2Z9JUGcrJkk2bnZeQ4V3Vo9iXibb
YpFelgQhouGhJKa6/VviwZGF0fUmFwEqymceM6fMpi/PtXvTWr5J/HBBGulV
v6G8cNeLt9Z8q06Ly7B+vSNpHxazV8H/hGnu0yf+pqog4nYsMW1scLuWAW+1
I6X4whBvD6g+3E8w3FPJkPHd4hU/ERpUBPnWka/NGe+F9dv/4MHACP/s3prB
gWBqUeWBkSaGhlSkPJzJXEKMy8eRvmq/a24K1xQLBk+CHELMeLzuxg77jL53
H8vryxeSLdsMceZON3wTOQL8RUfNLnfLQhJy5MczxX3KvL6pCtSZMcVbLu2j
h5Ha9O0qii1hjrCnA9qssXjbkGtPEl3smHoq/YtY53QnuZZf3wHdTrs57AOi
MvyPapyZaJtc2TcMpXrkuh6IDIgvVWNVYpUOEOnVzKTYF9cYkQQ5yyLCrfbI
UZULK2qElS8Q0c/pBCnTbZS2nqHOugOAm1jIeunzT5K6ShI5RmeQ2ooTqNEY
h5EAEzKcBHD2jGyi0HnvfAihO5+N/HQrgRiKKid0Ym6WxlN8J7pdh/NfaYaM
vehjNBNqOQ9Yy3M3fSeGPOHjAt1iJnxTGwoGYs9NwuEUHvyZ/J62ealRt8a8
wNbONkNOqgycPlX8YsITpMg7oy1FxfWUSR38nTubz476t8++f0bu9F3iVfYl
rGPA9xS9vK9DgkQqEE+OCEWDpd7UvuF3BI5DZcaTDE9DLkITW+WPont2BnB9
aYsVDCIH6V5SRHP+RYSNxgicvAZzUw/5/Suwng3E1gtyMwtN5Gf6J5e2KTzh
3bZSaq5sCicyeyK/0FPuNOkm4VLn3slvDwGmbe6LPtnZDv+T2jut7QPCqGEI
SD1icCKFf+pYLO0cJ3/C0mlWOqAy9ltlayFW44/Gb0Txk3f9mJvNHD94I0S0
LHFKc0/m4Kxw3nZe6Y9Shv5aNvgZeKmnlf4K0cHdM2tZX/UC8n3o3WC0s+0Y
g4eSUSP6gHIUpald7B3ju0Fr1oJhkjVz2cWAUP1BvsybtBNBEBv9c4v9JtUZ
oXfH/WTWEHTQ1SnLl7Wouw/E45gpTEsAtvhPIbYzh6rIFbuODmWBynBFFqJC
/z8IxJapWoJG+ElfVGhffoW21yxC3nD1/2TINboKVwa7aA3x+4nfyz7krFdv
wTtncZ/DRSeCVG8B5KaGVZBjEnJIwqUJu24KyTGK3aNOk7VW2KOnyvjBFbBV
Y36lxVixopgNPWegCNzXTU960Cx168T3Rnc9dFpTEA+mBvpIVZkcqMQ87znz
LLuE3/FeT8firFNKyTw+RtQOsYFtJ7/UJxq6T+HH7ByupnvOEIP6upn1gHAZ
M263ZPa4akPu3DKy5ruSw/Y7rYxukmj7pYf5/2ROGBgtAOi4yJSfZ/bY5VU+
ibQTcRi3QqA/fP3nN36Dkv/fAnrLn9btqTeskSKZ9hsALL29a2qE3ZakQfQj
FwRVRHcmY+tMvLmzuQXDgzKM7+lyjqY0YQl0nQLfuKo0CNUv+6vVWrlUtkU/
nrHLmoSEXnQNho2Z+tBMJ9u5NjrzbOlLqGpvFgBoVL5Y+q5N7pERKLk5XNYR
Ra4jF5rRS3zbQgo9FvD1/U2dMMuc66IqFSYBHyHxH3eSE4eZsUNB4se/I10n
psc989X31uv1axf1LEC6lWxvKZimYyyaiDdTBS71GPjYfxd3/X5f96QJyhxv
8INA8rC7RCQvGrgaTSla+m4OUa/kGuxrVw+9sk3TFY41VlEICB433UUW9f9d
eTG6rG5QpSVLCfvRo9tGAwfUYXIMuPNZF8zZcBtVC6AlujE0wuuDoPqlhZWj
LSTxy9AeUiG+44IrVfi9/Xf8kLAD7kUAWOOCk2H/tVB7zM0DJEqAKuH2YjlV
GK3+eh8xv75fIJWxA3vD6qLLzfp+GlP+vec7Ld6a87JGWgiNliN2Lbe4xmwM
JrCiZTZnB56OH7ZdxDzbCxd1x8xHmZ+TlNkcH4GasCiQaMB4Ki3VwisEH4gR
7GFYyaf7nGOoUhBCKjMM8+LplL82eOgbksI0iFf0wfXegZO3YjzslOsxBglw
9WxyGbG6VZUEUJy4HNwUHSsblOr4W18S+pp47mAbgs89NW4ZMWK5xBb9JM/J
560I66q1zXAs3G5Nzx4qyo+dKZyVx5C+eBn8hTBLhmj91h2qXAyBMmPfLFnC
riJWO/z5zww7K1eQ+j/JE5YW+vLqIP+4rXg32PMRknxNcCsFjJC9w5I0lDgT
xcjYK0V04OE9XuiZT0yd2XXiBDGeZ1QaLPVPVoVJGbJnFQAKkfyOT0POjE4/
uxiy1Ej0UTvpi1ah9nzpbPo/og3JtTcHSsqnJLKtE8ea+If9uJGkzIXkX1Kl
F+QAFoSbMLIYMvRl5d4mkLLjhg7GxNkvnO2ACySbMtHFJqsrqFN8fdKyggxp
3nZVN7HtjH66NZt8l3sx4IQcew+jKBHp7ROPSqXb6eH5W0p5ALNVA65LRnHY
Mmj3nDF/GuR1dj/R/EjNGXFBlRzAQfqHWjf5K2ShA98+1jk+0bK2xoAF7GCd
iGgOw+LhFoPg7xl41YsX1t1FYJlztDtS736rk6E38ePAW5taMce/owcmj1Rc
dyTfDY7RrDaXSk3CHXXDitJ7WOVxq1q3ISGvsdErmPrG14obaWGhSsP2AUD7
xiGfFYxJWnrh1K1ccD/vCBZhUJ9mTeeQs4igy+7fXkoA5AyJ2ynV62J8HRET
ikNrh1SfuisrqndLm3/tbSfEg37Xe8uXMuDt0GamJWsHbdFvdBQfvUNPu1wY
FVor2IiE+7RW9tylW8E+rDMmFvXcrGrWl2KU/bcJRIrDAbsas4VxkC5++T8Z
tKvBKiaIh/dVe113kZPY3pcoKSRIR3n0mIshg0vxyo0otlstUNyLYJlbCn7p
iyCwWBZqy0EYyDHifFt92iPYHehcxrNyRlV8jJlFsJ4L6bVZJjWRFRa+QaWn
keGIJ1uNsIJxbumFTsdXbfhrrgKkqaP5WR3lw7MMFlubPj7KBxzjT839OscE
DC0jKLh3SEVfrElymCmAOuCg9KITlbMCj9x83sjAFxERifQcu0QY2CJt7Nsq
wxx6x2V4LRFWcskcrINTDAMVLJVuzoPmlwuToCUmJhU4z1iWfJZi22pdX4nc
WU2PX3GLVeUGs+ZPMlX/YK+YDzS8peThasgXGHLFmqIlKC+vEdPJX09w7z3G
sowJkPZD0LNOrxaGH/cwVLbc/xWHVCNCp3nhuExLksFDWR755UcEBbuQGyBW
5u427uwtNEvpflzTHOFMrBvMHCQdGzlbJTZN1c4eXT4VCNNithgvvYSh9ye5
TrsZNIIOqnC3s2+gLDtZ4IYc5f8pk8GCuYKtgLquxwdWWgXDaOcpOEFtIR+k
vHS6O4Fa/X0ear0AQpRwWrpKM4b+h7czYJnNM0MELZ3LGAxXyDyU6zIcn60B
+PYN5MgjCAg9rVrqxYbimOYZd6Jwywj/2JjTbWwBKd28u836qf2uc5nLIH3o
oic8bUtlatCXkTAQ3a6Rv1i7TaI2+D90I6FerghbrThe3L/wW8R0tI7uh0p8
r8aoGgXj1Skx7sn5DuBeETHXxEP1CnYd6RlpSxBzhLRtBINEk8i9i5+WfdP5
NGZuxdrnaRFmYLR2vnNLflKUcpsWPGdSNw2l97i4brdW9VZrwKRE9FaGUfjp
YmnYfQoK0gWlgVZqvprbcSlRKA983mpJxOn0lTAANJscEyKL+cS63DasoJ+M
puGlxghk2wyHqJRcTQMYNYoV8MJWoeU9GcEeC75gvQ9sKfnXdsLuDZEs3ZII
ynl0ajcJwBn+4vDtwWuanKEJP0Wi7pEsXhRY9IFjHY+7KPaFUx9WQPoeVpEG
dmjatgWzM9Vol8dyMJvurqhrxujx0FwG28Gdwr7wt9yVHIMslyPV18lW1M9i
Js5D42CAZIiNGJ4Bf9I5CYeYQ2d/YtoRL59GrM9WFvgQ2cfmi8+BAey/YCLn
e64D3m/1N+6o9F/O3V26z89yXi98tIaz1g+lERgm6Bq3yBz7mOpQ9dwNPyTg
RwuclIskJ6sqCP5Za+bE/rUJ1wBC3xsD4M3TD8cVukrzXW+xdvGpAVJxYWCX
0nt2wPJdmI1/FXMCLYxGTDbUTvrB8ZF4VhckcaXt/Q0jAO+0+CgHNMOsDEDg
Vyjy16Bf/j/M1DnwW9u+tA0maGW++sDDcI2y/wj4PuAJoZlYno5aK1K9sIA0
ObY3f3TDB8YGMcZXnaLilBfjPaJiJ4QPVvD7G9zxija1rKS3yD1tn4g+yWBI
dcwD3a5V8qtMaALhechLSjT5vlwIIXi7b+PtmUriiEzX0LQg4dpB3lpT8MMx
3CTLyBmbKuHXvC3ceOiqTENy9IAHfhqJ5PvyNtjZSDaEZs7MpViqlqVTYpmJ
dTMKx2RTftoHe20voFUEsfMGicycHabBUc1KpN6rBkeHZ4o1rGzuno4eAFAk
38+XjHTmvO1CxKJYPcmuAkWroT7x8UgGbJ6uQ45G77hui6dTTsBhyCImxquD
9O2PBQWJbv1GjhY0pXcQGQ7rB4Usi3GLPCtbQ7y5q0qWn4SvivtpVhi7rFGD
csb/we4346l9wVLNJH2dTHJa20ovaowLc/5a+kJlkcbzKZPVyPkuRPkKD4++
CsCUlg/aEepQe8DCxd26p0Ihw0oLmAkh14Q2kIhHjuWuKkDan1Llnf1eEOm7
VUQQ5JV6dT82dsxZZBebZl9A0C51GxsTpz7vGEzTK/xZTYep2ZoTDdBrV8DZ
TdYHjqNI92wQGt6tM6OOOcnYvUmf/X/woFtnMVKpiqsGgi5dUJ1pTrgapZd3
ng0U7E3mpWl/+kxBPuCSpGEmdX9xj8G1GGQlmEqRzhCEhcs/tbAYXqn1hQP4
xu18X+AxktzFmo2XErnE0vlC4jotsWvGURsw+qYhPLHDHxqd6ubodz8S6/lr
ywpPP6wqERpxppBkwdnRe2kOu3q9CINILGJGpfciP8nS9eskr5HwfeOc1K/Y
8nRFZvnLdz4xtlzUPaJ/vkX6e4Mq+60d1tEdWJBpROs5nHlkAtZBXot1oHq9
B84KtQFgx6OoLT0jZtrhgoZHAP16l6GCJLASOs7roA6bDsK+sd7TX47mSbEG
+ahjmhfof3lQwLoW8D+liRfNemoPDioApurAYROSQOEqR9NvGiQFGKZBvwgK
XEe9FtKFeokBggICNW/HN0ibpmeycBBIY/k/kuDAN+ewCU8RHBF7v5f/L9Z0
qhnNf4fLEh5xODQj5dhC/J4yfbbOv6m5CQ0976HgWN70CU0pz4FsyePMKDQv
q0Hl2mMqEpcGJX/dyFZMHXJMWndqZLvX4xm+3oDMD2tHHHBDppg7Xc/NtotN
8AyQnfoZjuXt5szB0QDbcLs/1MtvGiuTtv/B6L6pI4D9cspt/uIxchczzgmp
2j+vcNFAA+57MBmX4zY+Yhk2wwyWwHgSvdjv8prondojgc8oEWY0Ug8h4Wa3
JTpux43nv+GqJ43RGS5Ok5ANV3/KSADucFqVO0H+Msfe9mcC12eB2N63PJOQ
nEmtCI+PgTktGO1sH2cF/FxzvXYbDIS8xCzCUR2Fg2lGZAQ+EOJmlSlOaWyd
wE6vSYYnOYnVhmO67Mvf50PoKDaZa/Hp6ojn5wtvkHrUL81c/blmLrr7W0Ik
ivhu4yD6NQElPbMOK33k5nfr64e0q1uQjqY1not386injS4QcELDIaEMNcz/
PNZ6YOwKAMBLq20RVNLCWfb36i+g1BgFJ80WS7SqUL++cGBD1znQcf3K2VL8
byIGUV8OvhLwUU6lwoJ5U/IRHoQy4oOndUWQ3xxOdSK1plqzSNGLFek5r5d1
p5+CfuAdDX1/es5uNI6nynvT298CSDYnOgbNENk0BU60J+NFUD7jq+srTaHD
uLb3/e1G0zgqc5sMy3G0uhoH+5xJRDWoRhMM7mjLdijrWhzfie5dNWwSVnHF
ANQ0cpY/mvKe0hyQDjth76nXnCH1UUAtrRU+x4VzzQRNhREi7RkPILoBPrCG
c2+aLAQ5ruGHVOj8i80/Ur4vNYIsNViMWd3hco9jojK5K9Wfqqz9QjUXeOy/
kKVyuf+kzFJiDK98VWMwrdKs03wcBeKoaKFpp4JQ+YxA2RBskYXPHUFlJeBN
2DelRhpxA7FDRYsuUklwz6OMoZlXaGbpVd8UkTsq876iXIsbdfIGUfiOWa3Q
ThCYQAOTnFCh3wx75vfpEg/2N6/8md6PsJTRMQ5LtW1aNju5BDlph15exdP9
XdiQtq/E+PawLbdwSfaEDA6zdLcCX7nz3fxdS0BWxfSeAd7OGJokn/mDORW9
+xJ7NNeHG/9Esp4qa7X7WAErugz+BHQJNGhv0wbyaXFia2Hb+pC5HgEFDeiD
I6TnHc9wH3u7Tc+SFNW3drXEZUtjJ8O4l08aXYW9W0cMZ+SMvscedYVwfopc
SKmVYkSLgq5plVmsqg7ANICg9IYo++7SGxVTC0aoC9nmuOa6LR5RC2X3ql+Z
QSgs0AH1xj2jr/smISqSkNrwKwPN8CuQyFd09xsckGHxi2rPXs15TkLjN5i9
3zvZOzvvLybSZXwRkkcU+hEmdbvLO81JSa30wqYK9kW28vIx7CZyAjxoRmMe
QEa5I3OXqYNyiml1olZ3obhh+ZmzB06sd/wKzIvgRSmxl5rLK+uE1Vzfhgwx
8e7ZYOvWstajlZgdMQsXx+2AHUr9Ev5etTGGrbzEJHzVQPdQi8C5DdIC+XJK
GdgNRoH5c/udk0gtkcumRJW/ITP8d75MEjqbmNLq2n1NDpO+Vgt9zh/fmjqU
H/HikftM9c695mJR/cD6lPVc4XLXTQp7eke9Qz9RUohoSmn2t+CBECY6YS/x
K5AVWsyc58g8RsN0VX4b/WfLNz3tVuUWy+VzMKI83gafpRSPzBPaQ7gEe7se
smc7TnABwxU1haG9RQBCTaKuarxQ62z8OA5z6+yT0d4JVbIV6tv0TxKxccqI
rDXmeF3Oqc/02/VRzrRPNigJPf1lZ+kWoSeE3rYumK5lllWF2Z0vKcJgkbdm
17vyl+g/jevLcr5twp1FfulJrGTFdTfzx8V8UK1DW9mI3v/jwjGJdVYg6ENj
JXRqMB0gm5gGyO72vLySUuL+Know2vf8gBiOkbvfJxwusghLCnn99nViKfb8
8gYDjYX6iZIh0chjHumtL0jKfVHOHWO4ewND0/8qw4wvXGktloznxvCavsBh
CjsOUo7tv8mPXnMwzgD7cl7qu2UX7MXGbk2C09Jzx7nw9F1Ch0K4JOR5gmI+
hdYGVleVrO1fzJL4+L0w0FVH0DB+7rEqmviNII8DQO4wYfjyzvLwoR6TGWh5
Li67I9VuCiarYGH/L+t3OY0641ghC0MRG+oCBX+jOljuT+amm+xvSO4S7CDQ
0c8EEMvIrt0TEAF75r1OUrHbseB6/ezCqoUHTytJNT8j2lOI5Vtghmr2xtNI
ru+n8rzm2PD6szk3nnDHZQd/4Ojr6+oYxOaqmzNfE30CCmmYyw760JkK9PLg
dHRJ505C28OA4Q5cQyaxDeOZNrl7q/AJ9IU/BNhYaekTTrOMUqzT8uEHS14L
FtB56T0k8Q/iCQAkOyr2JACsVN5pfGPtK23C2UPZkPnbs6Bbycyu/lF18u0X
ZVHNBFWsFsAPxElEiND1cXFoW12pWMfsAhBiJI/niSRhLQz6BmohtkFCMzh5
JWDpMRDDJ0/9eHTttpRWXIlk0SyYrZcUCappeLOx/JTupxVDaJpB5PWlwZAt
fGjZxxB2tLW0aUJZtoN/ddWglVhbZyna4zoy3GEkPBmfrLfU4B9KCWWhuAsQ
dDO33K0olFeh9m5VwIBLSsmdWvY4C3kiWo5KQN2s3Si9ZEypnpCn/aaBqr2A
OvcZD+s2+Hmxm0nrixw1GHRue2xv/PA4BxCp4n4MyZlEivNPdKVLyEA3n/9X
BdAihH4O9coO3H1m+4JPAaVmGwwS2t5N2myLDn6NUpv8XKLph2i0sw7ffkmy
G8z+V7d8bqyUpjy0EbkEw0oE6LEzq+IvxQJnANHAiTH5lHZf7i758zW4hX7J
TO08yBvvYjYf/rziGnE2iyVRUCbP66BvS+3M90lxald59ufqr8fBOJ2WyZBJ
sDqIHl3U2AY5NtETRUgcGJ5aFxp00SU8mr/P3ebLI6bB2H01j1lMeO7oK0gX
m762SwX3/0/8wqn9lpdnjwHFc6KS0I7V6r7bmsJpoxbzG3yxQWFyJK/IZ8AF
aje+N22BngZcB0hHUucP/miYLZ8a1J7sH6cYy0xrC/LrBkmRxNFgtopLDLTx
lmRSTMc6V7uQnPwGNn8wdLNyjnzRaCVdvbmQEp6YQ/FY+iH/nbufsNdA7yes
PR7Vb98ajebuwNie/kWs5sU5472Ugf3CFKwLGB1OCx/7/hO9loACzNrYnwT1
Rl+K5djBX2zkoja7Zur+BZH4u4u6vcbMpJCCSRyhpcrVtri0dacaFSoAH6rr
3d2PGbNQrVeUYX7pW754VvVvM15LwbCgvQAW6k5Ai8RxM6oTfomKSrmlM6U8
vkIKXn5gtEkfvX2NxIoShb0GdYLB5oje1BoQfHNlh0dI5nVI/m7S4p7rsz+c
v5yxqHbcT2Mj7J1SHLXVMVOWTOuq6yWXe+JBVb0lOZmTcC14fAW2w/wRSePb
iYsk2B32ovJo7Hn5OvqS8gpAxeMuQmWyViS0/MahnVs9P5sXSJd2xUIQ3ubg
Ta4i5QsVkkaLMnVtIbrsgBOFSLyTOouyGNjwBo1wmol3KDFweWNzglWCQLSh
PkVFaIRgrwDKyco8EKPzksRyfhCpIsl3DoCig9trUi7sWnsqFS0+zFVXCYiM
7i9CI76k/ti0pEH3nWeVQfuxdWqooU1BXBtMC1sqVXwU6PyTym1qYm3TVOm7
2lwLvK3vEAB3Fdeqgc0FOvqqQW873isiaJ54zlEHIMQzIGtdaNaocHiLcnZt
GzIBSRz5cuRCCj6C5O7Jf5EHr/SD2nF1S3WDGMH/k3Ko1aDwqzXEUkvCvB3F
+ova+xyBZPyNXuvGZhoGcg9aa+dO4p30cH7rlRF2AEjjM7ymckx3sxUUD1z1
0pkc2kr5K0FeXqQUjSiUrf43Pu3kQQxZmmBgdMNLUaD4jkJZS7k8TcE4Z5ng
S8H35RnxikgP7uwBYJ+/QtcjCEfwbv58hQfdmEWjdtrcnZ4TDGEPzxHDGFNa
qIR/HyhdICj5Qmb8CoptjykQqgKQR+gQAmECHMiVgRjG22XvSTlokyf679/L
DureTcNBI3JTN74EnQm+EUtIxXtHtz3t8AZJq0QMo5mGFv4A691878s1Son/
iKKO9CtRyC8M3FpGNQx0p+qydfESoPQA9QpGMhf2U9auFAhpvILfflJPlnLQ
C/fn0OANcLoTmvo7nD+LLas/hweI3rPHOlrXnErt5RMb1+snlVnqQj2rE2JD
zZSo1QuqpFKyI8ZyfaaDgne2fVfYUYLGcKfErR2CTPwGuUGBZ7R4JzfCK/hl
gSeV282tn/R+laVgzAC/yuz12zCGWqRd1nLq2hVsw5ma7sFcUH0sAyemG1Jf
6XMZlYaNVSkyu8rrGgq/88qQN+vY0y8RanhCVXO96pS0Ybc80GLg3AWGz7CR
NlWRlP6AthmQMZoQGYzyLDajdH2zjn8VBJjubK367V+lBGTi1s/SIP3bxA5A
/0g9OR3CcNQl4C846VDNTWuyPv9T1hsXVfiC/qBzlL/reO0B/tayM5ip2sU+
iBAuLIvQBkkX/uEUkjBz/VFHc50I9Fs9cOx+OWOAJH9vUVCLTjBWtnesP+Rz
gb7itsliSUQjpjJhSgI2/2iXhRkgszyACCQJ6u5n2tKKMY/w/wIfzDLlAHon
vtBvxUryIKIQZdEtwtxDPHMleA02dYHug4kpfkY9SyAkw4WSkIFs6s3PPI72
/3V6aPpnh1rLMPxMy1XKICRoMW5ihnTGZKHB71pgM0Im9+HiFvAjrQTwAqxp
5XKESQShlAnuDtxJqP+bLXc34bgYbtiKKOnQALy112H3yndLvyY+7JGoC311
/IjndDnGpXdF81VBcRtndw/Hdg+zXcxPuKmfXztnxZxU0lY5bdCbk9npAKGZ
wTC0RJ6yF7x2p+hPhUHYetWigbkWMth5pckWqhEaGULKda2SgqKUon1Duc3h
337epqsx++/NVuOzRj8GQpwo8xLb2oRtrcVMMxuEb531R8bwXeUZFzH/+BFM
QxSmNqE3L1PtMp9iK9bpJ+H95Z+F+rkdTRvEL76svN3nAMdNL/o84vKcuKas
TsF2ITAHGEhkFow8voj0ERcFzc9e/BqoEKpRvfFz9bgrZxlA6KcG8d51DtK+
xN1A471FMmuTKwTWkWxtUS6nps4jOvfBoLHdKmfhbj6oXriurXCirhqkdMD/
6zZwLm71gnleLB4gVqi8zPGon7XozvbvWXWgImazJsM8+ABju4Wv3EHcbrJ8
P4hoU/adurw5HVFYDn/LpaJ61VykzOAQdL/Q2IvENFE1vswVK5tU1aGITr6c
Z5I7m7ZS2TMHxcBuPAUhkevzl9lRfIj9bcZH1cfhbPweDV+mGcdhZgb0eZMm
y2c4ni8nxRMN0B9CXgikcWZa4rUIhsHRcubev1Bs81xFGGU+fddUdb+tlRCg
I2t0ziOKsRka5dVPLflCDyCgAAoknAyroST5pP8Dajks0MRIlP3JxCcrX/km
jjiI+VsH9I9mva5L+SsrN8ZVZXPycrhTJn5r2HhRxJY9A+23zu5UaXT+Nxf3
k58SauSllM0BFCNmQ3FYRgmJtHwOac+s1BRs7pU/lppasWVngGgARJjjvLC9
p6srnvaSmo1sp5rzw+ltvYPB3nMxvYz/24rLmybFgBUU9R+Mw4vayfaUEsK7
/jtszhxpBPb3z7VfMRisDj+woYezx+a2VN/FSFKS+95IGSLaO/B66hUFlMMS
zediGSsq7iqH5FlEg0wxcMKD1DRAy8zZypKlko0s33fMgt6CE7VSnZoEyyUy
ZWY1MbFaDQtly+ACsHyDXsY9Rc4EzWgtLVYL/HiwtXhiYbLL7TJF9ONYB4s9
XHdn7qVOF6ODiivy52Cj8EUKJFDP2YpzFx6zUV8dxar1Jz/E+X12Kz+YCSHT
fW2u++qMZWw7u5jni7NLFWqDy6GmeVXLqDR1VShZO4xqYUjVfDeNdOr3ffD/
vM+pDZ7nEbyykag3MhGhpDThrGlEf+0myJNvkq328r4XiyQVu4vJfiAiVr8v
p2fFGUtHglIwq246e3cRUGt1j4s4kGZwEmDqM/5V0PTy91bX4JLz+VO8r9A9
DEnNrQbo0zcRmyOBLbltkBng6tezpWUFJ+ibeL7StH3zxDP3ySBah3Vpn/Y6
MmiaTGAxjwY2qhZh4WPKwoP1ivTYFbIzFUGG2EIzWfEe6cfThSnCUChFMD+M
7eCkVkoBGsmYTkzIktfpJz3o3q5Tny1i8Sx5eAzhq7KmxD79dI15Clqni+EP
Ov2S/cIo9ajKsYNZdLa4hji56Vo+Pu2iIQhzpaW3G1cp/l0VKbZ/E5OQrb9v
Y1yhvICXPbQz2bvORoIOh7XuJQLfHpBkoKLhJtK6C+1uagvckCmGuGc4YGh5
FXPcxpbTHAB3i4wGBGM5ZEh16VOtKfWtE9Kc0fZ5sCSbXvu/JJI0lhYgcJCm
6mof5dXV0VWrZ6zMM62O8z66cU587YZ0eQt9o/Nx8LotoSu/eGeQBtHBvfKE
bK6aWWHBQSXK1a6pTkhqh56io+foZAt5G1pJQpXM6+w9u7/DjPCaX3HCrbLh
e0i8FsfZcGOwHp3v6TU2PDG9dI6jua9EORRaZjrLbnmleTbS06GGRsLo7+qg
uLJbjwVwkR4cOCMuTLYEGlCWeH8OV4WixfFLgYNS4o6Lwu+JBbKZ9WnoogUv
BEF+xjlH6DjLa/GTCCJXw87rf1wTiWDrMmqcPwZLYfxOg2lrTGUEidVRjALM
8PJoN+OsMgtDS4Nt1bko9Xtx98B0OBCTxqcohhScMYQtckkKuDk/gJuP59Px
UTpzDr+pQvPUkfU9HCuQ4cMbFC1YpGr5jROfrpx8WWOdzmfBjlBQPaHZh6WQ
F5wuNv3yLodf7rEsVfW8wVZu3xfrrzNLtnKz/AsaJsHd9ctAQrX2FaXvA8yN
1+yGsf6feJkIbEMYLv6uL9t2lU/5MfIzF9/vMhFJ+bl/vDoAk3C0pnR0AlJ/
S7GInFIeXmVhrfIlXKIGM9zxuEm+qs/1sVa/KoVWOfxczaWNQPNCJ2NQfrbA
CmezkeAQHRAH9XowkrjFsnzhC82/LZg371Uc3ujmmHLkL8Ey68Kug1Or8/Tx
KPP1HQkuNL1H89IQKzCqzH76uChJWlJiy+nHWPW0SNvqj5QpyNJ+cJ0MFTrd
KJgcX0aM0d8Iv9wHzqVsrxbIKjUTfF90YU01uQK+k0uscGzZ3g2J8LmCf3z9
0H9Cxx7FtmpM+nNLwNfizrOl20JZfAQy8HUOfG1bTS2bOCYo8+Zdq0PVoPKO
s7JypKRj+e7dqJ7qLfoQ2nNCF64gfxX6cxzzbND9uW1i3alcqujW1nWh0GJ3
9GhrBiNcLf1ttoQGsO+x4y6v01Ibvv3pCFdSkVX9BV7JWfKrc94jYQBnBzUy
hiNp5XUIV3c5K5QueYjHQ84h3BzBtNZ4TP1U5SSloVc9PeKZ0dQMWRqXLtSX
mZ+KId4jnziKM5l0CXXQHmlIIxdHgh6cGfv8MS5hOsEafUBfpDXiFFSLP+FV
1FbsO5osMo8X8biX7j0xYuHcmhkbgM016D0yHhEVHrMuFC/ZZ+VJLJSS2d6v
WnNYdHH6gloetMkQ0ozXWUkw0/hhDnbWwm/ZdYF6hb7mAJJF6/zZdP6LAsHh
7BVLuUMJBbVxa5d9jYf+U5/Nmhb6A/hjZ1JGKSHK3u0EWcF+cIQklEAGHRcy
kHTkpqhQaimuoyhwvRWa4GlqtIqQi7jZxNq1RmOUJvBH4jGuTTOlwL7ERkrB
NyQ7IQelofZjS4JJ4jANtcjpyW9PlbAQYOhFkP96T8zNeN0mYHGxwZzUnNSB
YWk+/t5lRftfKJI6e14jIoZPMCsV6i0McSgp752eUreH+m4H8aHn9dq/zY24
UcLOQ8aEd7HjPRDLTphJzBnQ3TVg1CWLFJsUoCcs4K5xpkuQg3eUEHIYpUFl
W9lUU3nATb4Ha4XCdCjR014pzHAMlemllF5psDnRYQAY7EBLqMcjeN4tJQjb
4E7XfItqM5muWgCV6HWTFjuXE0OvkRizQtZQKFt2Yp4p+mMYMt8wIKzK5Kuu
KKiPfqI07ND+YPh13VvTGzAgiY42LrGLdfnh3TxrtmV6JHZ9lY+uLD2I

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3GEHxwzDtPq0nyTLeZaNv3DO6+6wzTq3RJ1qBvoWVdSLsIKycdAyejspfkRa435slS8igaozJOGjZWrAaIPpTWqYHTQ/l9s7tA/2U2x3Ex02LDAZSSnxdDfU+tYUIVv3p/Tw2k/v6dx8E22r1paQAXS5149qn7zwEaKmtBdy2241taKvvDtPbzlnfM+BgOql/QWEGAQsMbloA5Bcm3NfLSoPXaZpBLJ9kbMhhp1qX2sQQumrOLgTsa7b72pobUJDIwIX2zmD95o0cnoH0nJb/59hH7y3DIi1QMpXVeQfQ8rN1Bvy7mDE7nwgR93Y3OuGN+9ggHnGfg/Fy65WEM9KrVxNl8py8npoIh6zKND3WJuev3tJgHSPghxfpR9XLoHhIvmMW7sieypLjFgMW938AODXPpzWOPzNGRaI+pWIMw2bHMDAxaH/pFrtUCUDYv1OfLmTpCC3JjwJkfKxmCAv+I4LiZDeoYUvhWzVVM6Z52hmCqJ3/3R6Ql/UbDvrf6ENmFH4Wi+6TGQTnfcPRY7V8B3/NryRwgB7VDaTzv7RVtzc+XaVoRy4lc/8p1y23eaViuFdjy2ff7tV6tt4BfrbcxKTLE7Hgt2SuZTxrmhfJVFuwAGDTy9J1k/1txpGox4Xlx2S2Ttr3xPaesdoY6HcRGdl4052n9cQydnY9s8Ww8aEm9NQwULGtXwWW3GGdxq3Uj86LJv0V3qlvVwKqn0LghpMvJCnf8d1erzKq18L4US5I/GGaUonvfymtA9wUkNbBTGGxukE83L1SHRkKHR1Ywf"
`endif