// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RrqGyVR3zsAlJ8LBASmNUNxZSEQbQCUf02sKGlYqQ0etyeynMo8erbL465zl
ayyfdjwig2cL78+jw75s0Z6B5FD+ElCb/Ic0E3W7mKQ681yh7VJPtDMDkwO5
yW6EFx33hO+E5nBmvb0+RhBh+dCY51MK3tLANYUE4WskCvSAuWPj1XaZktx6
tuRvScUs8todudXnZMfrn1zRQXvUpdfNNGuqMay9ICY7oPmKwdIhqirlI+MC
okRaI2b3wzm7FE9BqKEzHWkLx7B3IcSR5kJSit97n8eyxIV7ZuVCOSYovHzX
CDpHshI/IaMbHBSr4DPU40zNjbBh27yI7/Uxyg2jdA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UNfjfHC+bYNUFXTkOSQwNnqVfY2DybRXZBRjX26Z79zil6fIk2Wd62vUVSto
2IA4LqAklU1O63PmN9aCEA4R7j67aAVBYP5Dtm2fliue5N+y3TkKX6Mrs4O7
ygGeW1T++5/sLVXq8GSl35l8jcYeUm2paIoNknc7XbrAG8QbacWSx/q4lNj/
Q55nfCdmNdcHuISaH5DXE4ZJN1WSq/kfSSCS9USpkESZdjbFFkffABK4Atx0
eafGRyTaZpNf8PxgrPW/1XrJ4u+QzXDA0C0DyO72ODFa1N+XrSlBJtcOMfsg
koW3o/vLAUn8BLkMfUG3LJTeqGALxkxzcvMREsrvVQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rMi/BpUZ1PbU+ON97E2p9sn5dVhXr1IZOUDM/qA1JN3+coMsX4o6KXe0o9yN
1n69WEw+Ib7G3ruaTE1BCE5t8AQdt+gH0jgM3Z5CTYOomG97ofpdECZsTJGr
1zhPvGZOhpNI3iYAJqQit6adb6dl2PxGiddk1yfgkhvu0pSIV9bJmIUaNEUO
8p3O2T3F8nz6ZdNw8xJ32/UnqCBZksPG7nQipYrebdmV8RaGf3qRuxiRQJDm
2FLfIxB8vSuRZ9bQBfgqa49C5R8IKoKZa+cN1xulOd3aTARcIJnO46XCEOTa
9pzGpOmIRQyFy9L7lYFgw0EyNrFdHR3OZmojwEx9Hw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cslzjDyBsaxQKrYQpuRAzfkkEeh9FDA52hW5WdBgVPPpzKaqC+iSX5kvDhEP
8UrttCgeqz9CM6eid7PrJrIeobEJ5dCf+saa362IOayopgELBsEqEJk+BnbJ
+9Ao6jJH8ey5tjDWLsrHlHlH+fJRaClhwHlm+qupNhLiozhcTqY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kaTvI0nJjRP7NXWeu2qZWN9SM1P7IJYIdc+7U85MeNZAzGvFm/PHplk6/yAB
zdxapmY57nV73F4u/dlnajAuaOLkMk35KUSLW6VqE4mCYhTbC02wf8NlQ/aY
DJSNg8vt18OFXfo/btXcsjtw5dElq7eS49R1NoBY7uXF5A21OENMX0ATgiRA
phKhIB4kjsxni23UUKqsw5kHo6hVlz0Mu9ayYEUoO9A4R0AHsE9vbzRyc2Xv
8HwPHqvPctACBBgaBLPEOLNLiojrJ8Si9/DEUbKjL0QPVqeIGVs9pcGpNs6q
FinyQAC9okKc5ug67uH9nR6XS59N6jMfUcQPca8mHoafzhpCAZ9RlsM/CyHa
URmPIfZIZ3jJ/fDgEMcHf8UCBHnReDudexEbI+zSSoF4/Nlwsxu/n/FKXifY
nZBOZYUibwMFYdZOc8IUfj7fZYvKdw6IphvHY/qxbvfHjiJ8iN2mFGa3Hb1N
Q8qV2NLnewXc4JdoIz/j2n1PeUELTpr3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jLHMgv3VQPf5/Nf3V9dZ+j9iiiE0iZc3y2KTORvamoFXEoHWdYimaoRUY33v
rCRLn1+5THp1Ig2RGL+3YFLDDNzL8LWMP/PxbtajE5C6IdcntEsPuJu3UoLC
1Y/qju1zxfIDbaDph7EdQ8nitAdM0fNa/KEQ2auLUf6jjtn2mew=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q1ubwsyOha9vzihJIsyZYVnkp/20u6RZ7/iFc2PS+yFDjTur6PLyq43/MEwN
OR9FKpJkLcj84FyxyaTuKnwrcAQVNWa+4u80BCVU5de6ZjezoA3vEG+YY90U
+LEj/bRbW3E7P/TOa5h3K0pEcf539T1WSSWdJWLI2yRpOlAeBjI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13648)
`pragma protect data_block
7Mj7tE+gHEiqvu1NcH9EuY5U4Wt7+G7J8PKOkuS5rBc+FDVZB+lfx1DYZ5DS
8EotHVG0+BwVw/GewZyizZLWdodGqDUUJK9K7g5MmQHGYaHlmx7t37MLTsX5
dEEVxiuZDgF4rc2OeL1YZIyAWbswfiJFNOuWuka1tHgM7mnOUtsytvSbt4TI
8iXDI9++s/edr8SxGOpMk2+txlizQMutnP2T3vXilDlP43w8cBHrST0IwiXN
5Z9Ig9ykBglfFGBUz/WcfPukCceuFqxNrZjpggpfyMsFlBafsVivMjNKkwso
4FnO2kSHrE+1lHs39kXu6Em9mLy9WuVBcHopKj5CxPoiteLtWZJQUwhuPtm5
G2NjWypPBl1y4Fe/vwBgA/qrBCdBGVZjcxis9zYV0ZWZbFYImz/u6LdeBiOB
Z4tmtq8g50GGEFC+VFchnJpdV6kiEidHteTKCMfMet+UQqXfJY7f52J9cKU+
GzVadS5i3K59dXDKM3A6mO25NILn+G9PO0pUDjVp9vdE5jS4we29bXOMAZjj
M65Bg3smadt7qbDfy+Yk/b+pUk/lkViYWqa6u5iB+dPTBNiuShIXb07SC9IO
eTVEHiwYQF0zThw8WvQYqHc6Mwpi+/SzqV8bEZe5ob6xLh+FBEKp8Oy6tQ9U
fUUzVfnvw7gK+sHcHQ/DPN7T/W2vger+/vXOc2LCPJfoyr9gyuwyFIiVRVFX
kf33CiY1mkyj+QRtg69zEmarA/xS+jhCp6ShMBENeq5Y8ddySyOAwlvMEpDm
X0d1BkVnx/+XU4WGDl5xA0eHwAdSaFccJPtjE62Nukwq0rgkoc0F61xvXi67
a8OkKNkGVFd1xY/l7U3uWDYxOHb0NqmJ4vLixqDr8T9/KYS2gm7QSIMhTLQ0
lRoEfR8CQnOaQhokvsuiCjqt8ilh0dBYKOtrwcX9gr9d1wlZ1CDreWbpv2p0
4D6j6Gy8TSZByx99pGuvceDjtYEVET2f18BFuFCpeTBYENph+7aNk0rsX0mS
MeVzlRgdEXCCzdiXwOy+58u36JWhz/wKHWqEjysf0aXErwNqiv7BRXZiIIx7
p1WUE7juMzG6sXDfP3t9eiAZRuQSEmIeSILTQtbs6bUqN/TbEnxOzn7XgGEE
s5m2sd9CR7SP7qQrQwO+AsayWDFeHgACgZLWFhkdMiWKE3daRVkfrm5SquyW
bgPREm2wtKIZQL42UujmBaQqwc4iGSR0TvdTMCuB+bzkHj36jIgZy/yXbpEt
eXda8pRutb55kBF+tvsEx9QldzDVl3xSkIpT4ZJvtVsMvdTI+BzpG8yuuGfS
+oQNSWM3DdVrhrp+UmVf70graqEX1dOl0RVDegMUFOgt3os1jthCp9P6KtQt
+K0reSyX4s6BQF0VktSn7pygN5s39HUcx+P2GiNkOv6nCZ1KBSZe5ej+WLj5
ol2vlCP1d83ieY5ksbZtcbZFyyhTWc9Iwxf4c3gt6SRld9o4U+QdA7kdOW1O
OXrTAZItyhz/vsp8VGiqQGt6TmGPL4X6/l0wiwkJNc+MMoi3a8GdzbcAnVhy
7jL8ULtAFrOtfA65uUHlNQ8J9l0KLHoG0ClXDaQXgojcm4lzLY5KtVpb9ffv
lzpIEK3swdtDv0PYN0LG6eL4TszKLSnpbPO3PSoOGDkU2tMASSxxCeXGAGTV
+WC1PLgIJbrT8KhRvbRy182+Ngs4/izYBkVTrWpVlc23U37EYE/5OjuNP3kp
CChxOwqh3N5dMjKAkQcMlfKKykezhyfU1/V2FFtiXLmVV4k3nHgG+lg68VUM
q8vRJQK1os/6TjyGgXU4iWtKQKnOGsGtmvDIbeF4uueJdVQjU1Mt0n/H68xk
t1/HEpwxrG4S89n35Xse2d0RKfRId/f0hrFHHsQ+gyrkz6VofTG4wvjS9y3o
Q+laiOXg58c0YeWNEUKYxwyX19jMfVsgP6wHTflV9ClxY14bXcBSShyCv0y1
HyDT5fu+Y8ifAq4VH9ruDG7YNrGG/yMOx57rO6enKiRNuFYZpnyOmgyTU0ya
ZWHFrGHb3BmZK76VJdmhvRPJuHSP8OsaKry6vXlttDUD+taPsbYbZfoT/jZ+
4evJKUIB8gxI+c5OJkdYOy+BQhBoL7Wo9klveV/m8aEA1MAIYbPZa2cuU1/R
Z7jsjrQjar6W0JdozZi9amVdLCG2buHjA8xRubJGFp//Tlm/Ru6GMSTqWmR1
NaFRZaqLymGo/2MO05et7sQKKzCYXnGysp2dlIRTlH1KXSFgT0tLXmD30Aua
5cbJCg2iEHK7MpE0ya+oEOirjdZbRTHGs1JsUIqbp1ic3HuFxWyp1NzuIpVe
DUaVQgya/jNziHdAKdN1Bimn8hnYI/uW96KKbzK8RpIo6yG+imW1TMXZ4JOU
6hqJmT421nsRk+D3swc7eg0QoTEL94bsauFjT/7tFwAUkCYDyjrWLtqhf2Cj
fgFtJ7yVMUmsbhk/Lo8nlBcpo44eYFTeOuNG73FJIsXlQFClBZ2JiYtslE6Z
uz7sv+nT284Yw26mC8uCo//4AZlxb6EjbBywF1pLLCdWr4O0Nnjae4jbY1TU
BSuSg04OKiK0ft1GISFR7mXAVWMP6SxG1JxhWxKouXEkOkuMOn0jNPGptult
UNUP7r+4uuBzfvPtIkN/aS3R8GUKMyQaIRy1cNFF9iWp4e0e8BD1pEv/zTua
1O72AEro3TCTyhFLn/HWIardZPiwWt6sNlHrSSbRXzRaHr6VT+YY4+Q3MCS1
ZWpdXRj7daIZfUqPOyFPCexx/H2XjjRAJ46dyjHAsB67mcb0pUsIaMlrkj7C
+E/+nNyT9lIpxBdcCb47Ar4bQmIAoWUJU5XcCL93h1KQxpKLt1Du+iu/fJzf
oAZOH5ABq5kbeNKUVZLJq0RldNelVZ32+V5SMa9WMlJ3pmC4UYWuUybbaT33
bcFx03dgcCYVJ8/qviyES2P5r+e8DQwKWvuJQd8Cqzgxtdfz5cqPv78TSUkT
nsSSo5teMKhFQByukKMgTzu/fD37qslrM3ZilPTPPq8IoXFAA388WRmTKE05
g5OJp8IuNcQGWQqD8VdrJaT1DiP8Mej2KgPC2fQQuJQvwMh6O+UUoGxt5mwU
IuDSnrHdeNlxZYdAX2Opd0MOGfLrOYOfptKODKUyBj5NLrhV7fOuhrd+ow/t
whc5svpAJwwpmVyXgd/OtXfgKCRWOk8JyrWwXyqDNibqA11vP3oDhSC7ddrG
KD6FRlB4wNSaPVKgtUCPExwQvcpTuu6V4Qo/6UEW/lpJsn7RVVTpwNSBZ+tN
WpF21OhMH2SiGNb4oM13UXfGeJuUbm/MNFSzsW+2dxe1V55tUNiNXjVNoa2r
6wmTNb9oe6b/saHcyC4ngcoGRKO8zqbV1s78fc3KIhZ7L08d4QWIDkAimKQC
SZjtOMzzpoFmzOUYR7Dw+L9/xzdZWLbXn73K6Fe1Tx3YDtmMC/y8a9r59csh
vqSkfp/5e9nrSuOvrt+JxsadlMdAWL3OKiB9aRGyzVNSyj/OoahYEIBQY5tr
uGJhwrSHDFZEcr7v8IGZBttB24+7Yn0L5blv4g8RLobif7dsdBbVVQ0Qa8w7
2nyolv20PshGRYp6+65ehksW5OnQ9CF/dULfoXzEWvcWExnr3Ch6AStk/e/1
8nsNm85jp+57J7HuPGLvyhbKjKvZNgYoEyCzWfdaETg9SX4wMjdplLhDIOEJ
lCCqzR0iFKY8ksPVHjnBHlOsHsJQl9yEbEcmpyXXRqL6Kr0uq5vHNSkD815J
FbMIdQ1pfMh2gmkCM9qWmvempfoO+whXgL2kZgV6hGz6UxRhvrxNhneIbirw
9twS0f99Q5J83lbmtO/GKgAujtnjJGZXMG+p/n0NY2ulv4+0GTWsazEYaYP6
Uue0v3kzNvxpVXC/037R+uM4xHqEKW5sx2MpAs/cpW3ZceUTI7K9iuah6DMH
ApzQgKWwoCKi3LRuKuDtJvfQrrSrgXC7VJOOJ5HyCyJ8kfnOoMDs/bxcOL6M
cGBEow29OxNEs9dKTE7zd35VAAkeMmUyxtScOun5wtIJnAXEYHUgcGoXUid3
hPtmA4ceaXF5pUHW0zV46lAB1rP4KwLkFQcl5EnOO3TQ1b6vkOyFquOWEuSo
NMhipMh7EnUhZ7gJCGrxycEB+knnwTIqhwwj2vpFSdzFXciF92TY+7urid6A
/KlI3mk8wGMibzqtVjQ3CYWq0UlShJ7x0h7qvO97E/I5GCrDjol+D8mMSbfF
6Ck/mrJz5mV+xtM+awM6FADVgK8jUivMnUbTp1jh7SDUOWbTqW+bo2Murs58
GLLAOF1z/D3EVHP0FEXUa33s0WtG4gi1uO12zW/Hg/f+hOW9g4qHxbYElGaS
tzfeQoA9qL4ozHjrsxgUk+CpQk84WM25laeVBVHyhYHWCLoH4/MG3OHyxvzD
+5vPKBT9/rnDa1IVzemPkMnSjyIR9sW931I5FBUqZSshypMG0kfkkyjMufS4
PDF+4hVF+OGKCWxS2K+Edkkp7671BVKucUHOLwYbzybNAyFlRGp2xPv2NlcM
EBHHxssKAb9RPSAlmxxCMHAPlYu4Y82TKfnKLrXySpq4KEVXUWHCBkyHODtM
4okpE+X9nSRIMcGIQX1137uAXe1xdSBFJAAKUqV9ODhS1W2JNBqCSwHuvwds
M2C1pCa4fye7A+j/ooJWyhh3lP7Nt3v5zl7+rGfY6msDHrMs9nE7wKpNBmZx
CdlZp+1wfOYtu212U/DbOoLNBVIXz35FLQgTdGT/XK1g6XtBdiK1bQc+6IAb
vQqLJFF8c7nYdn/PM2Kc0HEqjPzyenP27guEaQ7c+QN9Bq5oRT9OZTbuO16J
KnksseMocWZ4Uke/aEOpxRqRsOkSs+EjEGvadI47HyLJfPvq5nEbJ+Ne7vSe
kltAJmeGhVOKB88rErJi9zjNEJBjT01T8Y0KkUMuw1U6+6yzWl2D0ldavqAA
eKUfaZEbUpfauFQAtbm5j3J7RdqowTV4e+w7Zf1wO0VnUKd/psQyBKy1z9Ku
u+L8VfokIlWWI3ga1Rhlbp+KNvCWntPisN/bYbxC+wfzWi5IOBMxUkEZk2vg
8M1jUUlXNFrYAaMOvfFnq9rXtjTWL3RKgdUpfTbRRrAyJjWL9mdsDH6zdPcj
oRKzpIX1aKKHsBF3aXuCuZQDL3H6VDm1BtSzBUvKdHEmfIyLs95Q1ZPKZzBQ
LlN5aLMzQ2CReTWjM1QCjh1P2GFBWdG2KP5TQolJj6Zz8+4+dgd+G4UPC+rp
hZkM2CpCOKmDHmCQIaBKfyrAnGvqvqG/jPnN9hcyH5ZnW74fPQz0Nry7d0Ml
0zXAwobR6IQPvZcw+VUd5p1Alf9jAXbG+qNcP6w5dgF24sjNH7px/upiz8/s
7KvI/hyqjL+X11bwG3db2x6LAyv3ijE6/oacl2Y/yMP6HkcqnNpnDZAujzvm
I2bxxUBayKIdR9OvgBls0DHbm3iFd013kWBdLOUqvR+tlgwV2vGOt8YI0hog
cRIWjOetHvdB5RiaDzeAEyUWc8gAWLzvNf2u+RoU+NzzhVidkI25GVOgJ8Yt
J6oQFEEZBKQIt1MfCDnayGpg8La6je2hKWdcAIw9TfZx/aKnj8H7O9wfzA2b
UdvuAUPMEKu35GgK8mwX+6vXTY3xh2inUbw3ERprfbtYhpZc0R+GMLxTcsqB
D0aEIdIzuHBe5LxS6ZGLnGxcYqTOIVE/h2pV5HIDp8nr23Gh6/6x3PF0x2cm
veq+U6V91yM+jeJ96yAUQlnTYILUAtI00MK71YuNbIZ6MVhBjN22Sfg2u2dI
zUVVP2IOVofAbpxhcDDMM7OoajR2Bl3F8KQeYhpWoJiaoPZXfk5uikF7XNdz
Bfp/ArXKekdRiX5sLlojD9CLKzEz6aN2r4rub0zDptjOq7N0ii3QRhvxUtkk
MJ5v1ZlJeYmVan7lPf6AlUkVopzrbul3YzbIvGvbV1P13JD43sRtaIbyS8/e
4xwWiNnsLiK4+0C6HMi0w1q6vunxTwF6uKBDElYWBv6Ervp4qhUhAyvipcaz
sZNCxW4ce3l3LAcIqSvkZCz8C+5OYAOWycDcuXqjTieHwCvJt/NTa6r3tpbZ
sNKpgIvqtKWX1B/sHb4r6PjRBTVn4EF/5FMKWVz4hfY0R82V7aII+c703N67
ABbNcEYITDxWGj3aaiVj8lX9f3vr99NRgmoNaX2yb18ZLD/wUR8TF/ko/ITu
sDnTeMC5zJmldDcbrz6LM/dqo9GPhCLRxjX/EhZErqfvV4mQUk9yA10XTGUC
MbojdaI1kSuTONqgao8WWLNk4Sv8UK1PT8BgKDrWRNMb8tNYB7e0Xo2Z4BZm
bvLKz0wGlArfjuHbbXmkR2sD0ZQ8aEJ0CRO89r6Tr6APsJtg9C+2fPiXuGmZ
We7+Rsy+wkp36iaRJdlM5bxV/3P7dYw+wLqgG+kktbkykyVO+6u/+aLuMO9A
Iuxot0dnxyB7H/svpVU5Zw7lgW1yeZmDsMls1VK0VRulaf/FoPK0Cl60ApJm
D6cRprcaa4Ep8IAiFhP0BSGA3rWF8whuZ1s+g07maywfxEd8NB2zCGQXX0qF
CSRIqqDBovn3FPqo9O/tXtk9YxhDi58WE38vrpPgSookpJmOPyjINLA7nydx
oD8kh0DfC9sC03cFPnarV6QKmKGw0ueMcFNCR5cWg0MtKg3eFaJOHggjxR5S
eU/r0p9WxpVoDzoA0UjGjSzr8+KzKzZvo6rBCDwB86NvWtT19hiHEPDo1FkJ
qHF1MUwTA854OjMl1Ww5valk5hvjWglI3kjYAZhByaMei6BzpwK/7P7v65Hc
4AzGuewWLpmkjCdNhO+5BdaOEGs/WmMl5Zw+Bd3wUCmDscG5IvouzO3Un5rS
kIRufrRVbc0eMZ5E5Fkyc07AgxbWPzB0sKzxDMhdtV7H6Q3uY7ndgVw5nEDc
RhWhLEI/XEP6gn/qd34pLA7npw3kyV4LwW4F9BC1LDMKmVRaVpwxudCSV+K1
itE/fGdm0MQ9AGmyr2ZN3JwPra8dGbp3aeghROdLjVbNnGzQ+8GqlbxP5H5z
Tp5L3oLkJce/4WpjQxIBZSsNyQ2Y4FazGXCqDHtjPf13P8woMwqjZDmt36Me
MbD4fqqwEHEkvGLeob6Qctgr5n5QJMUAPc3dTNwgtFfknM9a45wSNR611Q/E
noPTWItoeyiqGX/N5p/zxPnRv3/yjdfDd9NG9w+TE1or3wz6TnGnFB+EG701
K9QaHFzg+DPWj0oqh/YJ4jyl6FUyJO1gBEdP0AmHPHSWaiN0OMHfeRK4yYGh
ecRO/MFclMtnLSto+tCUJ+ExF/QnKvN5UAPZUyO8uhHk84tv1s2mbKLEM1M+
X4ly0cWJn4K8AU28hFyp4qHyAb5aly/JR0T57Nph7e42D1/RYW/BmQkCTnTW
WW1MVMzkOApN8l3sscOjmeHuAJvlnPL3Wc02MPQAO8n3fynrE1lhFYynZDTv
4SVEHSW6uQw45u0LH/7hruAMY6JqmTRb9rlseAVc/iYoOpLZ8e8YkQnT2DKa
M9DFemEYMsCOw7XFCoYy0QUlozO8IqP/UOo6YdrjqWymXRXUAAOPehQhvl31
R8y95Mf6Zt2hpmKtim0sqE1tylzIuEYJYZveVaXLU/2wEjupbVpWPqjzypJ8
oMgpp8OsIMnpgdxxbaWkgGVvMylITpf4FB39H58e7H3aOIyBq+/1MXZKnO4H
/zqRDKmnFRSC23oGq5ZqWRBT77JaVAXrnsuUTa145osEBB58HvQ/664hwsy5
JIl8WyewDRvFIlHiR62fRxcxkvpnKcQc223T5M3q/+O4hBq+hiSzphWApkt/
TpZ9bKAzggPLPYv+yF3A86ZHG0tTJYJfMgzmBBiXfKob3XWO5FFKzQyeqcXq
YIBZEMAvEqrohOOFysM5lE06D7E1c5kaL+2CPw9j7kUwA0vD3k3GeiIl7eZd
Gr+U7vaNTN/BzwgKgpcHM/9C6nuk79+cN3mLTdcF7lrslNDnU8Ox4gddZQNK
Ey3P9xoKCCeUgWZ0sp7KpHTikt9VDS6YsmEcSZQvxyZr9PhulLVGrGgry9Zi
Sn/9XqiajnpeNbokOz315bhUiAcUsyOHhmFwW6S4VgNT0gTGGPjk6vn5Rcyr
zgY3IiQLvBWXyWZWs+ymKdojynuzz2CNC9HsOesflNrsB6YYkp0uETN5jH4T
60w3IU6NTmtE+KLBhW6Z8nFnCsy175Q6UmBpwOQSD5KZ7jbidAMZqrVAeNVB
wqiuE8oY/8MQaEelcSXjJKT2uWQSNY3VKxvU8/sLGuTZzHXoeZCMktFy3lRX
qbwjk3GSxjVgdhSi2AjiZlvY/C7CPLWQWRG0NES/o0pf4nTNv0Gb2hvE9tIE
bp2K5Z005MPS+e0eIqJl7AFvwxRlk//vo2u7slVxvwwNKuu/Ii1YhyYqgFk9
xuHCqN7Shc77uiZsFi0OQlJk2I32EculcWkVLyypyLzRwDi7IGWzWItnI5sC
tMj4IZ4vWn5KhS4+xkA0j7cxAzCiDB4CBClTkGtffuUkFk24jmg2RAIq0OXW
3iSNI32w8j8zPkALAazUvakQyz1tz+im8BxiEO44IJD+6EXDwB42vb0aLcLb
MnhTwEtnWvdSQtRkRoa6wPg2Q0vf2HoHtOeabz+ChTL7FWsxb3jA74sY59J+
eGMYGJnbzAS+Z5J7P/L2+NOaSbrsDtUX3BBtq0t5lKC+rRrfpewT1TsgHJUT
iL3z37nU6gsgp0lsdDeVzLy6VzqrRy466pArCXob/b72CSAfMPl/xi89e37o
RBgGf4tBmWRKsPGVwJSGDY7XZ0kAENEBhriq/immYY5qURtb62BjqEhon8Dj
7LgXMHMzK/NpWDoYC2VH//mNreoi6OlyHFdn9Q4qN5inbcrDwfVHebV55Gg5
109c2dvYCtVzldi+oE4UC0xant6HmgI0ih93z7JZZ84m1pK61pqIfONnenog
0P+/RjAWAa6lAJ2AMaT7EtJ7x8L4eoXyEsZL8Xk62RKwXpwjORbubutV6shU
bYuNDumHQTX9jJAbIyPrTOYMr2K6w+arjAfz7xi7c90ZkbiLF7uhDtJop1KW
k5w7BgNLc+LJ3XawmFMJnI25wZD2TOW7/PIps9GIftT4v3qegaoLA7uYnt0L
Sl4YgWZW2Tf8p2vdS/L2HSl2tCVo/KAXGMkwqAIG3JgWlFqaVYQEO/nGYWDT
u/4jZETRlCTKiY3xKJ89qh8lUYVCLwvm/NoI8h8RfTe6QpA/9SwBfR8DySXc
ZS/eK/SynSdEw6UFxESklVXIjNkf4JIFBupUrjc6P+yEl3HtKjVh9syxgjL0
cuHA+8I0gitJ7Q/og+7VBHUz03VjRIghtVkxBstsUCmmxbfucKsR4cOruQWs
QU6mVEAySFYYS9DWo3xr2LCF0Iu/oz93DfuOcLYXeqPJxn+4S5aZUU6KA/0k
+m39WhuexDFzgzDGUBZsimKUicU1rL+gY4IFQN/WFmHgHn/iX2gwwk4yr94Z
Jtlp0DdEoD6osParso6y21UQbM1mNyLAYY4luPbkacMkkZmRh0LRkqjioUo8
vusqSuKg6ocTsW/fM/gd20hSpViMURs4+chYuCUIP+hBaavwLWG5fDZW1w0r
YRregA10f1Mfm19PtrLmF66Nv/Kwaph2h7VyYYSbV1mOsa7kdnMgVrbEmadZ
Dbq0mfGVGSm88w4xmXdMS4kDHMRsW68P2M8nUYEjtb6P6C9A/Rq/j2H3Mrla
YnuYOPSWoZXpNfc82Z0IVgFBYsVNVuxkSx3LKVp/HOH2k4sSyNwL3dvswF4P
vP6kBjlvwAyzq9fr8fFbEJeDOi5srFImAhDbetVkyDqjqfzklalcGktViwlo
2xtQGdpZ+b7nYOsWE3dApuxY32D03z1eZyp8wqI2TqCYfNrI3+wZX8b1Q3xU
EmIAEth5r5XMLM93VDtbnJj9gQ+6nfVFvFbkn/javNxCX/4QB3jX0SRRoAIJ
nJ0Zqc8XUBwSBeBVPcnNS7v6Ei1wMULxsws36QfsXnjPnyfALnessEW391db
/++gOViEgC8BiNmOL8PazZyujIaXIIe8RXQasYwRaNn1FAT3OGSMnMLL0Rap
utZobgqWSoN2p0fGg7j7XpMZvjGh8G5HppfkpQja/o8dKP3RShwFZ0PLy0vt
hAn0EMrncLO0lko6aRci3HQAyGdqFP+nsjFMDQJx+P8GyO/j6m4GxRoSf9Lt
ub4IiqeKhVM0v8JQovbGSHq25p0aca1bB5uMLG+bfk4q2q046qTmO2TaPpU2
tYWPurwpQO98ojK/xPRynXwOay+YlHwMaaNgmuIk/+bwrWXoHV56zAO+gZwg
2QvhpO+xnoqjFe1nHUzWDOemqmLxdXIYd1k/3DgFOkSss0O7QZiEMuIlPlJt
BKdwtrCakmUimsBPO93qhAZOJfYtC1cFd6YEkXi01cKue08Wbr8eKF0ZZinJ
qY48zvCedLa7/3wM+4Eb1Mfqa5EkDzU95J2UeDGOIrmaicEofRtoMd79/A9K
JBYdtnUaA1316Xrv9BS363p9WOkr175z70JRW5fvmmHxSGoNX8OtVU5xRK93
lTnaKM+KMQYhc8ZYT/fIcQEWsijmy3JxmXhVuKQqCVuJyBAi24bXJJqQQIJg
0RErlvh3g/8uKPXxqkKhmfqj08HyV16VQ/+yUqpwqD/gKd5DpxF4bBUnpxDj
/gX/yRX338E5+Mg1xE9TfpDvYAGAoq8Nm6lmmaSnHe3ySVHxAX9Np9P+qygs
rsS4lSk4+efL3DzcNR8zjMBJ3H7MAPWEaHOO8Emc2C9QTRqyvekZchHpdUs7
jEt8W7M00yheiFWL7cW9lsmhjDC3MTlSOwvL4LCDKoc7EyaWf3XdfuVUbLq7
gA788u5/GlrW6n9my/0X2qdCrCGsA0rN33RoybPx0gBHS7/6xcZhfLesuwua
sqCFqPEUffiOK6aGeBQ+zIfBddVuzN3PMYk1tc2IrY27eJ/ZGq2Zp/vv21KR
gO1A2RxzBEB1rISmu1TXidYQPBXS+ldu+br+Brzjh5j92Lfl8dkx3X0N6SEG
nvza8mSIwjNXt9Ix/gHJcomH61rRPW1QZiILiigYs7AGB04s3fX6azHRxtjk
r587eAusfvVQB702Y4i/qZcPDBQ6QSBz32nbRMWf7cgkj2iBON2EimEG82/q
7FBd4MbozmYUKRDI+QB3+zn3qy7QqSJ67cG7uJ6SW2BBHh9sBBHGg4ANsVeA
yv0DPfaUYeTqHlWQl1UxfR8oYtVrdfzAW92o5TeGu66BLltzTbaugzK/ws22
wDIx4sm7m7XmO2M58HL43k2DjUOV6ERvA2fEwRH4QiNPaNz+Q0mhXF9a79VC
KXy8QwyC48DYjBfanf8wCJY1Kng1MmE7NqjaVXVTmMaOw8sQHZScNdERYcuK
jYHa2dXqukUlb1/CLJqQaXd8veaOzVzuN1QSGC75Jx+lupSsiCvA5rJkox0s
sGCyW/D3g4By4AIpGyaBLvsdxeE4F6m05QkYyLwc9FIzdeaAUji5IeOLTute
wIkJSCsML2S06VHc82rHSWL8I36XR0OvZh3J6je0znyWdwkj38gsfNUvnkQc
H6CELLDuOjo9JsjQrpnivO7xGn88eZXIFWTj28KhY8841ldNNnBinf8Q1HYe
u3l2Rfq5pRlQyfrZqPrfnx8y/yRtW6GFNjQeHa3b+uf4tMupIIRzhKw7QcbY
CU88fUDDBDoHAB2dxoBZd76XE1xVXwfNIMSq363Q85Kijd5G3ImLaqSF+V9z
BcRzSmAG+y4F6bvjm+HD/lTqJQPYQ7E2i+XdfRyB1CNyKS1KWsZMs1ioPyxX
3Suyi+W6ZpDphGL4/jqNMPEJYKd9R1QWmF8FZvSaZU2AJjVzkUOjFaVHVzOC
u2bWJOvTG3C5/t8R2/uS4APsw4SLBggpGzW35NPGhTcKfjzyWewqekMhYlFn
NXiXP5Iiu5eoS/JO0ausp5fDRBPnDnoFJOkTJ8P0qg+vJH8nlY9xtZqET1Py
zKcLu7KoSmm0nz1Cm/01xkD9wePDlarG6YkdOqlD2D2lQKF4MT/FUJ8tHmN6
i9NA/4bVJBamGmZnpyV+1Im8h1Kwyk9lCWlUwhxTGYgMmoWkLwTpMJUQkfVW
spvesekKj243x1S7X3avPSXzGWbeoTvYDjCauVEEzL3Tf386oHd5PcuQOyhf
qS1a66iwukEd2vS1L5XwBlxUONKjceP64PgD+u0LTIJt83entqXq/8yLQ+Dj
QV32/oePVcy0VFsj0KwDSMYm+iW+Q2ksrEcRhp1SbDZjudqYJAvrc+gH+lJA
VkCVUJErmyekej0lMuROOHNq1rJkY/9EpyAGN0TqBavQFu+9SAuds4y0oeyH
MnVp0r9Os88DishACANdy1BsLSqHgOQ2Dgp1mfm7b7C1DvtjhW2y7g6X5/bC
U6ygGbCU50BQkSiid44Ts6IQjqtTjlJQQbhqiIx2SKu20bmku3mF2mdLRrvC
u9jTQTOGoB2vtYtM0qnu9tV9Pp5NTpdUWItEzXf0nolzrgkHzj7UDT4Ni9FR
BVbkRFgjV60r+qm7Epxy6coLvlX8EktMBPEAjMtVh33d0y0XHJG8m4uMSTLy
wmaXVstZhJRWMHfjgI6YLtusJi+G/Lx2GhbYHRnELe8fLblkHZ343qQ3/OOg
5nd3x0tndC0Ay5zd3nrR8vcZ4lOJkJDpNHeGg9g36+FFH0+xHMw9rHlryFWu
6KjmxdXWLgNPWdMe3G31hhlDtXbiU9xgNmKYPLMzidkbCxKmMl9/p+XL7oGU
f/oDXANk1rQNEaMvvlACKvYfXo2F1/UqhDgZrcq2ZpCZ27CKslNK6bUZea7F
+p0MFxaM1mEuvr/CbtZJiSxTEn6S34Jedgw051cFwqReVXJfmEELKrlvjIVo
KG6JmSMcgU3Pq81QdC5pq5bEWvskkOqw9ZPtHef/csnbdKStRvVx4gvTugiP
DwOdgRfK6n1oX0OGPLOyEnD8lyfAJIySHKTQiFlZjudBkYtK4XUdwP+G+wAg
ydxf/Daq12Y7Oi9OVm5cCWIvV/7WGvnRb5jiAenOs2w7fSDtB0ETyFvO9m0+
4s3NFun3veDDpjlfblOqIsrerAiyw3ZhkAe9B2ee7yNHBVpDG0ZL52OXSeh3
bqlVEL5E/Ea6hYj3srzqOU6vFx5t5gAReOMLkiQVgk4/JCK062KGhHGo+cO1
iY6jb2KdABMBT7j69PLKj77pVRLJwBnCvWqT7B3H+i3nI2/a8i698hRa9jNa
xLo4PJBWw3L1obKx6xbt8wr/8Bzo26TBp339dGFywXXLrFZlVbdqOeX9RmwS
4W/40MvTPw2Z9357MZL4bWB+GDONcqEqgUHR0N9WOcERq3Ya5hAMsqQKqqgI
hEsit2NZe2aisrXZKnmlUonY0aqKqXir4Q4bOnlx/3mJnGycCf6UbUoHTNtV
j56u0PfiNw9YwQ7vDVdpjUxlfWH1mZFVHXrcNTh7I5tBEbp4Ef+BEsQf5T0r
y0iQ4Yri57lPpRFxdXObJm/aku/3Jl1EiHyQf7BAFmYk3/NYXW86DEjE9Z2E
F8caiAaCnEeyc/Pajslivw3c34eKCmYnVJshtVScwv+MQF2gdApETtE5jR0c
O4SKqcED0ZzbFsmuNASfm8ycFnrBSW+1lmAObSEQgECXDcrMNATKll9q50vt
Yeuo/IkTql+kIdLS8XirP0HaNFEtNzdBG9qT6+/LIm9AFKWjHor9k9fYOCnX
WQncp32f0O8MD6Ja/z/jjJ9dL5rjmTiimCmXVIzggJp9saPstmqCi9KpeLQq
dRc+QyN4+VXwgHXukJHxmsD/J6vDvfOX2vshJKkhGxnDdGY7u9eW7K1jY26Q
qrcLfK/N63k3lmo6/+3kHZTd70cAXRKRTcsZIi1jtjyGWmAosGAHLoE6cxGk
sKH8POUIkIwlOiZ37WG55Oxm1l6TE+U0rmIQY1wiHYwXsZx8mjuZT14drYB/
0Ap1JItaGWyrGEdNtDH6awTfwJQQFhCpdEIaBnvoKQihYHiXMQG8RiLHvhbF
b97+wJYJVFyd2mZNh+haNlRIVfJ4L8tmdCQuhJIymZt5QhBvbW5stqIVTYOL
5CDsNUHg0p7IuY3s8AreoR7jCMagvwe5yeNOnvBeNqUAMbky/tAL9XuTCJHR
7xgTccpDCyvqRtnLuBUFeybblQTc8s4+VorsfudJsipvf8uyexvsJbzAVTMX
1mBTgdSVt+UMnvKAj9hMmS3OBdHAHKrGijy51f38hrOqvuG3oxsd3OT93u57
MrSQXfrg+HbAtbXjQI3uIo+AsvAw8yFEwSikoil/skYO9IXWlzojuSfQXk7a
X3YEBX9d4W61TrXXc9p569PTLVYm+lrarI4qCmh7Yy3Mujxd+k30l8fRq+gH
JnKqykdGEbq2HQ0bSP2PcgtUgJutFgHVrb2rPuxbKd8OaqBWiixn+IdWWMe2
zfIj0AztoStoGK8PIFsoSpn0DkNmvuhdn6dZOpVzpR7ZNStOpnVDpcpL9ziT
wb7PaSV/N8IWbLtWFuVchwaFo8AYgkPCIcn1+DmRx0geW01dP6vtZd9Gef4V
5E9gQMAscsuO0YAIPA+RIKQEXGV8oUD3hMrLIdO+9qBPbMSQVWAPWJWx6V++
hwICS1BcWOEGN/9ZgEZu7Wd8RBpdpdeZYWE383WXPOZibsc4Ue2CMmt1a5aS
c87lN7pgW2X4eZ7JjnHtUPXacvu/LMOAFZXb5Mn6k4CUr4WA3Uw06m3cBmlm
ec+TeSYHWAShodDIYBLSBho64SPB5ts5oS9rz5ZiUwEU5E/7jqgTGICxGZm5
uFqNvFnkyBp6NYaRSbLeZ6QDOJGKmMGrj3JD/ZXgPxFFFItHpMpZj5Fw42Xn
iiTByEpINHPJJIgt4O7d0/DSokiUEc92z4HEGLq4ZNf55gBdkLHtR6nb6T/I
2bzTw/j8Yxy+E8x+XWsXTMQZ1CdRa+kPz5rHlFQfi8HzP/LfkD+uFegeFstE
jEsHPrMlVJMTIMQMHPwgtgmezKAdpszHyET4fM5HtBD77Vhe1NIAnZsPB5iU
JcEIwcEMQBH4sgoqjO0pBN5uNWuoAQxw7qCpi4gzvnU6lShdqsiRKC3v3Dtt
lPOn3MyJAFUoF6L/J343CqUVvMA4WOjOPIXExQEjYbVuSuA/3nKF5Nphfl1q
B7dbdOpTzF6kSMmuHmc9Q3/qZ0rzyQBoAbc+fZWgLv9sdFT8/8MGNO4bPCSv
4/Dw7vrk+guRRpdULqGZVern/LDYvhF8ttKvEkdjDo7paXe1udOEh495PI+Q
0VfEzZwB3oD9sAWE3vfptkI4NXDkW/8ce6dBXYNFBPp2CSYTdwGtEwlIohdP
uVkmjitcC9CAIFDywabC0eRx2itiyell4toBLVD/zg6UPja3u29t8S5GwaOc
eoqnezVl5bwvzN2r3/9sePCqtvU3PqjDISqh4MhxrzHII49iOrnCS2maxIoV
mc8SYRWlGhssS2Tmqafji6HhjpqO3CC7fXd83JC4w9qTUePRhye7UuWVzgbO
d8zWkKSusi7p/Vzxl9fj/+iPh8n8sDFE/DMF/ILYWg46QkKanIIXhjUrTUQM
VAFbMfmJgdzfPlFMq7QqXJF4eAzj82E/5Ywy7cBKlacp/GWSmq0Ejg49Dtdx
ie+guOfAs8pfo5WkrITlVjDxEp7T2J0Z5IDlvDfx3FUTdEVqsDvb1hKhE4sD
wv4BG9FPrTDpRzQfMuwn0gUDetnF1rT1nOVs+4StSuHJCHB+hkvQF8zaQ3xX
tSc7SwbQeudH2/KA7r2Ua/axLq4qmaRc9S1ZLk2NUq75bbw8BA5sOBSmPgwQ
SHb2fuoGauHJK2zcARLYozYZMB+05UzjgKxZwsLMPPQPCES4Nacy+1O0HU8y
eKEQpbZrMkNE320IGv7NUPOcdKO7e3IY/6KIOsQbe/5bM4bIf2Xj7nteH8P9
QW6yqXg9KorAhicv/fI6isGE67gqA1eJ4X8buoEkwV3CL7DDuHGJydd6kvcn
il6qivj67wOYfQHcsOiBQUvUolhZ+xtYpMx/NsKK2RXfhhZiwA/eOD179Kr0
d/aS7VPJHx64mFekMEDVzweUZQje1v7CujkvP2FjZbu6/qw3ouub3Rifej4V
+wFRdtzN0sT4EuoRVzeAhHXG7LWkwYl7csep7XmfGGw3j6IIphaTXNjpBTaH
zDeikMvRq42Vpug3WZpjN6ETCKlntbfNH5oxWQnlrtgtYPPAuf49DkJNoaMw
VW1dLtDTqvfcwzfD9js8HvNjkR45pEtvGwFjARpv1S261t7PTnVaxZ4jk8ha
jc0eR5qH1KzGqh/5l5BThcBh8jIV/r0t1gqo1rYxwp0ki4/mSeFopV8eHUp2
zZLnwxnWlHyaAXz9VbTNi8IAnF1ltl5IpTESivZGfi8rpCfYPMlkkjlmq0X+
tpnZdzWqmFZcNuq7XPR/w0IiaQq8u623R42EtDoGJbD1eaPvUrcITg5fFVmB
3scrO5mmMKuAmGSR+QzvClEtZhvpXBNthk/mgJyTO5YHadA483L9AkQ/WkWd
JYFPbvicR6oXM2O8IALdAffvjGtLV0fiNdfYL6h7HVQfIbMnzuC9GqBAffKl
huqTJc3o0DBL5T0SK3ch7VWHfABWJes1pja5tVzpfM5xJgceUoqjjwU598Xu
pfXDqSdD4hJM2AodxhGzVBC4NQHULWFZ3HVtEJh+P4qwn4t/ValfrsLTK4yF
T9JChJmVsib2vHo9LFKhrX0FwDV9J0p+XPqe2F1vZGSNC2YXGt9cSgBjYIMb
6JBCcpqRVHpKPMd78HkOai+G+cHcJIlD/cqjAxsB3yPYR3XkxnjJqpthzfIn
NMwo26XIae46c1PPece7SC4jyHug8kI3xAB73nzmUauTM8NkWsu8JIazBh0f
rqtppET5x6Nbz4AN2q7LZytyRB3bnz0xBePMtt/9s3yOSEM95yvdv90UDuTu
3zQjloSMJw5Aw4vcY4fxZTASYU2peI6i1drQeO9sooKJxcabM8RePRCmcm8b
JtlMvArFISYrIZYtfw2grg3kVKKGRLx0MX8wIfIzpvg5U7NZQgCi6Yx9Ru3Z
uj50a3Obhy23RQKB7duZeo4eC+GLGTYwR3lCz6RJbbGhdE6nCQivt27I0jIR
bFeDiWcF5r1A9gcvGpScmXG/5mHsTHF1JUsMZd7xz0aiiBpYMvA/m3Mv95Qd
zzXsAyk41sCe9aClMdhqdP4/S4LLi/rNCSSr0bPghyJ///6jjQiaX6IJVnsL
dkAUHHmpGKj8VEuRubHepV7hcIQsAjsXuCJX2oJ/LNGYeEaxoUWPdf95WXLv
sMhGzMSyH7pxVg3b1OPtTLHXczknAIaXN2PN9WgwRzJFoznldD7q3py/CfOS
qEB81BayyGxDeTA7JljZPZEJGVhlkG2nPdBAMd5Bm6m2VtgXTPIvRSXcdZc5
+HGpbyF+ZXsBZWpHT2W9LT/MS/MjgUIibcARQq0x28WAHfhHCmJbj99k4yP+
XmELTgVG5PT1rFQVigjDo84IpiCTf5Wb0EFgeK96K96h22B0RKcd5IHCAUtP
VCesrdvPlztkJHvy1eMB6dOF1f44UinX1BmitRKuIMJP5L+EG8xGG0muMzIh
gd1UpQab45I2c7/xMUKt6dI/XrbgMjTYG8ToHsCiZ3QQX6lPG6SxfEbqn8iT
1Sso/WnM5PKeqbZthMbJgLpJlPR/ok5W6MwlxHVAS9jebtIaWdkjT33XNSUu
8rgljUVVoGKokpZ0V9PUo19WVj7eYDeGyZEr9qDQghvGVoOtpCDZpwY1/LLC
LgcPyd9qwXTBCcC6xZnC4GeesV0KRDXaxcnTSm5stLTggSMKJGL8E1wOpzma
fPNmDRl2ZzL7cwxpEymFpIS2oP/7/16M2TGRoXsibISeG09QZw9QGRTaHnnz
p4wBbShG5e6l+s/tLd4UxsYREN6aSYjcE9s0p5ouj8pYdlLtoThZZC87KBAw
SIQyDnyqKgAiPDi76gYFiVGMspgLJxHyhLG0yNfD1bNzG4WoA9XHZue4hXmu
6kh1x0ljMHvNCmWk85Bxn2iAmTpFxkhC/4wdfxyEyvcEOrg7BOtfNgAlZMMz
WgwVyBDghGjPoX1z2w==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "6ILtXxwzhwHEl3Q1IZ8Aoaw+a3ni57H4pSJ4X3f8I7yWpedZqdD3iZXXkX6phyUDKeHSBNnWISAzDEqycEtj7YD906oUhtfGdJvEx48mhAll/t0fbYL4tQnW40OB5ne7y6mbLhFhLGUFjKH7grphQCr90QOHE5zC7aUC4Gu6SXregmsplYioX8ZT8NmT5dscafpBby6ftWSAgQWwtp10AtGkl+gXAht/Yenyktn0Vx9aq/5LFSFf2A7CfhzzUbnbV+gDwi7cTtVc4r84JfB0HIizfxr74UKmKhGeTScA8yFvim7ia1Yg6hE40EOFiJmOE6Lw3jxtwXhD120clpmSSBn7lKo2tsi5IGgYIpoTDqEDqKQoaKsbdKTa6U+7BJhgQhhhEQbR9PYzLM8u4QRwAGml0Fj1sWgSMH7DZIj3SYCB4uPtpowfgbeNUeXTcIlb4Zj3WximVbOtEoQc3HHL0rW3skc24Bp62taScav9ktUy5Mu2iaSga0bzqQc5HIKzKUiHXUIBwPEZ0Hmiq2kkO5+o7wKphQ0gLotp9u8GPxO5kOHd4GNLFk2T4mSfh2dQBoXL5K8wqkouLzOfw8oVBwDz+9k9nNqX0yxozetQP6lU73IfuJAf33bZ7VCMINk+LWuDkm+rifsXJAM0CbUnyf7LuNjwgaeNBNIVEp9Yt+2mdAjwxTwFbPrd9iFisgo7MNpN55nrjEN8XcgOrVZDIMMDojHBmwvP0w+t2RrsaV+M9jwhrWOnF1vzuir+MNSiwuOfUz6APQURkOPWm1jzCCctZOTaw9NoEs88v1uQdzWR4gcRhCKegJVVZlc0zQNrimWQQcxf8LSuj1qN2pZIQ79PR3/2BOw/8LffT8O89tLfff8ePZb9qUQUFebYdJrsEdY9DI/Q+dlk6oHOUNYF0hLWeYB1TGjNPTK3yH1HBizH9Y5u/suewwi11BmYKoitVvJRioQ6vaFv8j6EKYMjb/tQ9n9IuaztIWDT1zjkO7TZh/BVJM/tfp/YCITcQ8d/"
`endif