// system.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system (
		input  wire  dut_refclk0_clk,                                          //                     dut_refclk0.clk
		input  wire  dut_hip_serial_rx_n_in0,                                  //                  dut_hip_serial.rx_n_in0
		input  wire  dut_hip_serial_rx_p_in0,                                  //                                .rx_p_in0
		output wire  dut_hip_serial_tx_n_out0,                                 //                                .tx_n_out0
		output wire  dut_hip_serial_tx_p_out0,                                 //                                .tx_p_out0
		input  wire  dut_hip_serial_rx_n_in1,                                  //                                .rx_n_in1
		input  wire  dut_hip_serial_rx_p_in1,                                  //                                .rx_p_in1
		output wire  dut_hip_serial_tx_n_out1,                                 //                                .tx_n_out1
		output wire  dut_hip_serial_tx_p_out1,                                 //                                .tx_p_out1
		input  wire  dut_hip_serial_rx_n_in2,                                  //                                .rx_n_in2
		input  wire  dut_hip_serial_rx_p_in2,                                  //                                .rx_p_in2
		output wire  dut_hip_serial_tx_n_out2,                                 //                                .tx_n_out2
		output wire  dut_hip_serial_tx_p_out2,                                 //                                .tx_p_out2
		input  wire  dut_hip_serial_rx_n_in3,                                  //                                .rx_n_in3
		input  wire  dut_hip_serial_rx_p_in3,                                  //                                .rx_p_in3
		output wire  dut_hip_serial_tx_n_out3,                                 //                                .tx_n_out3
		output wire  dut_hip_serial_tx_p_out3,                                 //                                .tx_p_out3
		input  wire  dut_pin_perst_n_reset_n,                                  //                 dut_pin_perst_n.reset_n
		input  wire  dut_i_gpio_perst0_n_reset_n,                              //             dut_i_gpio_perst0_n.reset_n
		output wire  dut_p0_ss_app_serr_ss_app_serr,                           //              dut_p0_ss_app_serr.ss_app_serr
		output wire  dut_p0_ss_app_dlup_ss_app_dlup,                           //              dut_p0_ss_app_dlup.ss_app_dlup
		output wire  dut_p0_ss_app_linkup_ss_app_linkup,                       //            dut_p0_ss_app_linkup.ss_app_linkup
		output wire  dut_p0_ss_app_surprise_down_err_ss_app_surprise_down_err, // dut_p0_ss_app_surprise_down_err.ss_app_surprise_down_err
		input  wire  iopll0_refclk_clk,                                        //                   iopll0_refclk.clk
		input  wire  refclk_xcvr_clk                                           //                     refclk_xcvr.clk
	);

	wire          dut_p0_st_cplto_tvalid;                                   // dut:p0_ss_app_st_cplto_tvalid -> pio0:pio_cplto_tvalid_i
	wire   [29:0] dut_p0_st_cplto_tdata;                                    // dut:p0_ss_app_st_cplto_tdata -> pio0:pio_cplto_tdata_i
	wire          dut_p0_st_ctrlshadow_tvalid;                              // dut:p0_ss_app_st_ctrlshadow_tvalid -> pio0:pio_ctrlshadow_tvalid_i
	wire   [39:0] dut_p0_st_ctrlshadow_tdata;                               // dut:p0_ss_app_st_ctrlshadow_tdata -> pio0:pio_ctrlshadow_tdata_i
	wire          dut_p0_st_rx_tvalid;                                      // dut:p0_ss_app_st_rx_tvalid -> pio0:pio_rx_tvalid_i
	wire          dut_p0_st_rx_tready;                                      // pio0:pio_rx_tready_o -> dut:p0_app_ss_st_rx_tready
	wire   [31:0] dut_p0_st_rx_tkeep;                                       // dut:p0_ss_app_st_rx_tkeep -> pio0:pio_rx_tkeep_i
	wire  [255:0] dut_p0_st_rx_tdata;                                       // dut:p0_ss_app_st_rx_tdata -> pio0:pio_rx_tdata_i
	wire          dut_p0_st_rx_tlast;                                       // dut:p0_ss_app_st_rx_tlast -> pio0:pio_rx_tlast_i
	wire          dut_p0_st_txcrdt_tvalid;                                  // dut:p0_ss_app_st_txcrdt_tvalid -> pio0:pio_txcrdt_tvalid
	wire   [18:0] dut_p0_st_txcrdt_tdata;                                   // dut:p0_ss_app_st_txcrdt_tdata -> pio0:pio_txcrdt_tdata
	wire          pio0_tx_pio_tvalid;                                       // pio0:pio_tx_tvalid_o -> dut:p0_app_ss_st_tx_tvalid
	wire          pio0_tx_pio_tready;                                       // dut:p0_ss_app_st_tx_tready -> pio0:pio_tx_tready_i
	wire   [31:0] pio0_tx_pio_tkeep;                                        // pio0:pio_tx_tkeep_o -> dut:p0_app_ss_st_tx_tkeep
	wire  [255:0] pio0_tx_pio_tdata;                                        // pio0:pio_tx_tdata_o -> dut:p0_app_ss_st_tx_tdata
	wire          pio0_tx_pio_tlast;                                        // pio0:pio_tx_tlast_o -> dut:p0_app_ss_st_tx_tlast
	wire          dut_coreclkout_hip_toapp_clk;                             // dut:coreclkout_hip_toapp -> pio0:coreclkout_hip
	wire          syspll_inst_o_syspll_c0_clk;                              // syspll_inst:o_syspll_c0 -> dut:i_syspll_c0_clk
	wire          iopll0_outclk0_clk;                                       // iopll0:outclk_0 -> [dut:p0_axi_lite_clk, pio0:outclk_0, rst_controller_001:clk]
	wire          iopll0_outclk1_clk;                                       // iopll0:outclk_1 -> [dut:p0_axi_st_clk, pio0:Clk_i, rst_controller:clk]
	wire          pio0_pio_master_clk_clk;                                  // pio0:pio_clk -> [mem0:clk, mm_interconnect_0:pio0_pio_master_clk_clk, rst_controller_002:clk]
	wire    [0:0] srcssip_o_pma_cu_clk_clk;                                 // srcssIP:o_pma_cu_clk -> dut:i_flux_clk
	wire          syspll_inst_o_pll_lock_o_pll_lock;                        // syspll_inst:o_pll_lock -> dut:i_ss_vccl_syspll_locked
	wire          pio0_pio_initiate_rst_req_rdy_initiate_rst_req_rdy;       // pio0:pio_initiate_rst_req_rdy -> dut:p0_initiate_rst_req_rdy
	wire          dut_p0_subsystem_cold_rst_ack_n_subsystem_cold_rst_ack_n; // dut:p0_subsystem_cold_rst_ack_n -> pio0:pio_subsystem_cold_rst_ack_n
	wire          dut_p0_subsystem_rst_rdy_subsystem_rst_rdy;               // dut:p0_subsystem_rst_rdy -> pio0:pio_subsystem_rst_rdy
	wire          pio0_pio_subsystem_rst_req_subsystem_rst_req;             // pio0:pio_subsystem_rst_req -> dut:p0_subsystem_rst_req
	wire          dut_p0_initiate_warmrst_req_initiate_warmrst_req;         // dut:p0_initiate_warmrst_req -> pio0:pio_initiate_warmrst_req
	wire          iopll0_locked_export;                                     // iopll0:locked -> pio0:pio_pll_locked
	wire          dut_p0_subsystem_warm_rst_ack_n_subsystem_warm_rst_ack_n; // dut:p0_subsystem_warm_rst_ack_n -> pio0:pio_subsystem_warm_rst_ack_n
	wire          resetip_ninit_done_reset;                                 // resetIP:ninit_done -> [dut:ninit_done, iopll0:rst, pio0:ninit_done]
	wire          dut_p0_reset_status_n_reset;                              // dut:p0_reset_status_n -> pio0:Rstn_i
	wire          pio0_pio_master_reset_reset;                              // pio0:pio_rst_n -> [mem0:reset, rst_controller_002:reset_in0]
	wire          pio0_pio_subsystem_cold_rst_n_reset;                      // pio0:pio_subsystem_cold_rst_n -> dut:p0_subsystem_cold_rst_n
	wire          pio0_pio_subsystem_warm_rst_n_reset;                      // pio0:pio_subsystem_warm_rst_n -> dut:p0_subsystem_warm_rst_n
	wire  [511:0] pio0_pio_master_readdata;                                 // mm_interconnect_0:pio0_pio_master_readdata -> pio0:pio_readdata_i
	wire          pio0_pio_master_waitrequest;                              // mm_interconnect_0:pio0_pio_master_waitrequest -> pio0:pio_waitrequest_i
	wire   [63:0] pio0_pio_master_address;                                  // pio0:pio_address_o -> mm_interconnect_0:pio0_pio_master_address
	wire          pio0_pio_master_read;                                     // pio0:pio_read_o -> mm_interconnect_0:pio0_pio_master_read
	wire   [63:0] pio0_pio_master_byteenable;                               // pio0:pio_byteenable_o -> mm_interconnect_0:pio0_pio_master_byteenable
	wire          pio0_pio_master_readdatavalid;                            // mm_interconnect_0:pio0_pio_master_readdatavalid -> pio0:pio_readdatavalid_i
	wire    [1:0] pio0_pio_master_response;                                 // mm_interconnect_0:pio0_pio_master_response -> pio0:pio_response_i
	wire          pio0_pio_master_write;                                    // pio0:pio_write_o -> mm_interconnect_0:pio0_pio_master_write
	wire  [511:0] pio0_pio_master_writedata;                                // pio0:pio_writedata_o -> mm_interconnect_0:pio0_pio_master_writedata
	wire    [3:0] pio0_pio_master_burstcount;                               // pio0:pio_burstcount_o -> mm_interconnect_0:pio0_pio_master_burstcount
	wire  [511:0] mm_interconnect_0_mem0_s1_readdata;                       // mem0:readdata -> mm_interconnect_0:mem0_s1_readdata
	wire    [7:0] mm_interconnect_0_mem0_s1_address;                        // mm_interconnect_0:mem0_s1_address -> mem0:address
	wire          mm_interconnect_0_mem0_s1_read;                           // mm_interconnect_0:mem0_s1_read -> mem0:read
	wire   [63:0] mm_interconnect_0_mem0_s1_byteenable;                     // mm_interconnect_0:mem0_s1_byteenable -> mem0:byteenable
	wire          mm_interconnect_0_mem0_s1_write;                          // mm_interconnect_0:mem0_s1_write -> mem0:write
	wire  [511:0] mm_interconnect_0_mem0_s1_writedata;                      // mm_interconnect_0:mem0_s1_writedata -> mem0:writedata
	wire          rst_controller_reset_out_reset;                           // rst_controller:reset_out -> dut:p0_axi_st_areset_n
	wire          pio0_pio_axi_st_areset_n_reset;                           // pio0:pio_axi_st_areset_n -> rst_controller:reset_in0
	wire          rst_controller_001_reset_out_reset;                       // rst_controller_001:reset_out -> dut:p0_axi_lite_areset_n
	wire          pio0_pio_axi_lite_areset_n_reset;                         // pio0:pio_axi_lite_areset_n -> rst_controller_001:reset_in0
	wire          rst_controller_002_reset_out_reset;                       // rst_controller_002:reset_out -> [mm_interconnect_0:mem0_reset1_reset_bridge_in_reset_reset, mm_interconnect_0:pio0_pio_master_translator_reset_reset_bridge_in_reset_reset]

	system_intel_pcie_gts_0 dut (
		.refclk0                        (dut_refclk0_clk),                                          //   input,    width = 1,                     refclk0.clk
		.i_syspll_c0_clk                (syspll_inst_o_syspll_c0_clk),                              //   input,    width = 1,             i_syspll_c0_clk.clk
		.i_ss_vccl_syspll_locked        (syspll_inst_o_pll_lock_o_pll_lock),                        //   input,    width = 1,     i_ss_vccl_syspll_locked.o_pll_lock
		.i_flux_clk                     (srcssip_o_pma_cu_clk_clk),                                 //   input,    width = 1,                  i_flux_clk.clk
		.rx_n_in0                       (dut_hip_serial_rx_n_in0),                                  //   input,    width = 1,                  hip_serial.rx_n_in0
		.rx_p_in0                       (dut_hip_serial_rx_p_in0),                                  //   input,    width = 1,                            .rx_p_in0
		.tx_n_out0                      (dut_hip_serial_tx_n_out0),                                 //  output,    width = 1,                            .tx_n_out0
		.tx_p_out0                      (dut_hip_serial_tx_p_out0),                                 //  output,    width = 1,                            .tx_p_out0
		.rx_n_in1                       (dut_hip_serial_rx_n_in1),                                  //   input,    width = 1,                            .rx_n_in1
		.rx_p_in1                       (dut_hip_serial_rx_p_in1),                                  //   input,    width = 1,                            .rx_p_in1
		.tx_n_out1                      (dut_hip_serial_tx_n_out1),                                 //  output,    width = 1,                            .tx_n_out1
		.tx_p_out1                      (dut_hip_serial_tx_p_out1),                                 //  output,    width = 1,                            .tx_p_out1
		.rx_n_in2                       (dut_hip_serial_rx_n_in2),                                  //   input,    width = 1,                            .rx_n_in2
		.rx_p_in2                       (dut_hip_serial_rx_p_in2),                                  //   input,    width = 1,                            .rx_p_in2
		.tx_n_out2                      (dut_hip_serial_tx_n_out2),                                 //  output,    width = 1,                            .tx_n_out2
		.tx_p_out2                      (dut_hip_serial_tx_p_out2),                                 //  output,    width = 1,                            .tx_p_out2
		.rx_n_in3                       (dut_hip_serial_rx_n_in3),                                  //   input,    width = 1,                            .rx_n_in3
		.rx_p_in3                       (dut_hip_serial_rx_p_in3),                                  //   input,    width = 1,                            .rx_p_in3
		.tx_n_out3                      (dut_hip_serial_tx_n_out3),                                 //  output,    width = 1,                            .tx_n_out3
		.tx_p_out3                      (dut_hip_serial_tx_p_out3),                                 //  output,    width = 1,                            .tx_p_out3
		.pin_perst_n                    (dut_pin_perst_n_reset_n),                                  //   input,    width = 1,                 pin_perst_n.reset_n
		.i_gpio_perst0_n                (dut_i_gpio_perst0_n_reset_n),                              //   input,    width = 1,             i_gpio_perst0_n.reset_n
		.coreclkout_hip_toapp           (dut_coreclkout_hip_toapp_clk),                             //  output,    width = 1,        coreclkout_hip_toapp.clk
		.p0_pin_perst_n                 (),                                                         //  output,    width = 1,              p0_pin_perst_n.reset_n
		.p0_reset_status_n              (dut_p0_reset_status_n_reset),                              //  output,    width = 1,           p0_reset_status_n.reset_n
		.ninit_done                     (resetip_ninit_done_reset),                                 //   input,    width = 1,                  ninit_done.reset
		.p0_axi_st_clk                  (iopll0_outclk1_clk),                                       //   input,    width = 1,               p0_axi_st_clk.clk
		.p0_axi_lite_clk                (iopll0_outclk0_clk),                                       //   input,    width = 1,             p0_axi_lite_clk.clk
		.p0_axi_st_areset_n             (~rst_controller_reset_out_reset),                          //   input,    width = 1,          p0_axi_st_areset_n.reset_n
		.p0_axi_lite_areset_n           (~rst_controller_001_reset_out_reset),                      //   input,    width = 1,        p0_axi_lite_areset_n.reset_n
		.p0_subsystem_cold_rst_n        (pio0_pio_subsystem_cold_rst_n_reset),                      //   input,    width = 1,     p0_subsystem_cold_rst_n.reset_n
		.p0_subsystem_warm_rst_n        (pio0_pio_subsystem_warm_rst_n_reset),                      //   input,    width = 1,     p0_subsystem_warm_rst_n.reset_n
		.p0_subsystem_cold_rst_ack_n    (dut_p0_subsystem_cold_rst_ack_n_subsystem_cold_rst_ack_n), //  output,    width = 1, p0_subsystem_cold_rst_ack_n.subsystem_cold_rst_ack_n
		.p0_subsystem_warm_rst_ack_n    (dut_p0_subsystem_warm_rst_ack_n_subsystem_warm_rst_ack_n), //  output,    width = 1, p0_subsystem_warm_rst_ack_n.subsystem_warm_rst_ack_n
		.p0_subsystem_rst_req           (pio0_pio_subsystem_rst_req_subsystem_rst_req),             //   input,    width = 1,        p0_subsystem_rst_req.subsystem_rst_req
		.p0_subsystem_rst_rdy           (dut_p0_subsystem_rst_rdy_subsystem_rst_rdy),               //  output,    width = 1,        p0_subsystem_rst_rdy.subsystem_rst_rdy
		.p0_initiate_warmrst_req        (dut_p0_initiate_warmrst_req_initiate_warmrst_req),         //  output,    width = 1,     p0_initiate_warmrst_req.initiate_warmrst_req
		.p0_initiate_rst_req_rdy        (pio0_pio_initiate_rst_req_rdy_initiate_rst_req_rdy),       //   input,    width = 1,     p0_initiate_rst_req_rdy.initiate_rst_req_rdy
		.p0_ss_app_st_rx_tvalid         (dut_p0_st_rx_tvalid),                                      //  output,    width = 1,                    p0_st_rx.tvalid
		.p0_app_ss_st_rx_tready         (dut_p0_st_rx_tready),                                      //   input,    width = 1,                            .tready
		.p0_ss_app_st_rx_tdata          (dut_p0_st_rx_tdata),                                       //  output,  width = 256,                            .tdata
		.p0_ss_app_st_rx_tkeep          (dut_p0_st_rx_tkeep),                                       //  output,   width = 32,                            .tkeep
		.p0_ss_app_st_rx_tlast          (dut_p0_st_rx_tlast),                                       //  output,    width = 1,                            .tlast
		.p0_app_ss_st_tx_tvalid         (pio0_tx_pio_tvalid),                                       //   input,    width = 1,                    p0_st_tx.tvalid
		.p0_ss_app_st_tx_tready         (pio0_tx_pio_tready),                                       //  output,    width = 1,                            .tready
		.p0_app_ss_st_tx_tdata          (pio0_tx_pio_tdata),                                        //   input,  width = 256,                            .tdata
		.p0_app_ss_st_tx_tkeep          (pio0_tx_pio_tkeep),                                        //   input,   width = 32,                            .tkeep
		.p0_app_ss_st_tx_tlast          (pio0_tx_pio_tlast),                                        //   input,    width = 1,                            .tlast
		.p0_ss_app_st_ctrlshadow_tvalid (dut_p0_st_ctrlshadow_tvalid),                              //  output,    width = 1,            p0_st_ctrlshadow.tvalid
		.p0_ss_app_st_ctrlshadow_tdata  (dut_p0_st_ctrlshadow_tdata),                               //  output,   width = 40,                            .tdata
		.p0_ss_app_st_txcrdt_tvalid     (dut_p0_st_txcrdt_tvalid),                                  //  output,    width = 1,                p0_st_txcrdt.tvalid
		.p0_ss_app_st_txcrdt_tdata      (dut_p0_st_txcrdt_tdata),                                   //  output,   width = 19,                            .tdata
		.p0_ss_app_st_cplto_tvalid      (dut_p0_st_cplto_tvalid),                                   //  output,    width = 1,                 p0_st_cplto.tvalid
		.p0_ss_app_st_cplto_tdata       (dut_p0_st_cplto_tdata),                                    //  output,   width = 30,                            .tdata
		.p0_app_ss_lite_csr_awvalid     (),                                                         //   input,    width = 1,                 p0_lite_csr.p0_app_ss_lite_csr_awvalid
		.p0_ss_app_lite_csr_awready     (),                                                         //  output,    width = 1,                            .p0_ss_app_lite_csr_awready
		.p0_app_ss_lite_csr_awaddr      (),                                                         //   input,   width = 20,                            .p0_app_ss_lite_csr_awaddr
		.p0_app_ss_lite_csr_wvalid      (),                                                         //   input,    width = 1,                            .p0_app_ss_lite_csr_wvalid
		.p0_ss_app_lite_csr_wready      (),                                                         //  output,    width = 1,                            .p0_ss_app_lite_csr_wready
		.p0_app_ss_lite_csr_wdata       (),                                                         //   input,   width = 32,                            .p0_app_ss_lite_csr_wdata
		.p0_app_ss_lite_csr_wstrb       (),                                                         //   input,    width = 4,                            .p0_app_ss_lite_csr_wstrb
		.p0_ss_app_lite_csr_bvalid      (),                                                         //  output,    width = 1,                            .p0_ss_app_lite_csr_bvalid
		.p0_app_ss_lite_csr_bready      (),                                                         //   input,    width = 1,                            .p0_app_ss_lite_csr_bready
		.p0_ss_app_lite_csr_bresp       (),                                                         //  output,    width = 2,                            .p0_ss_app_lite_csr_bresp
		.p0_app_ss_lite_csr_arvalid     (),                                                         //   input,    width = 1,                            .p0_app_ss_lite_csr_arvalid
		.p0_ss_app_lite_csr_arready     (),                                                         //  output,    width = 1,                            .p0_ss_app_lite_csr_arready
		.p0_app_ss_lite_csr_araddr      (),                                                         //   input,   width = 20,                            .p0_app_ss_lite_csr_araddr
		.p0_ss_app_lite_csr_rvalid      (),                                                         //  output,    width = 1,                            .p0_ss_app_lite_csr_rvalid
		.p0_app_ss_lite_csr_rready      (),                                                         //   input,    width = 1,                            .p0_app_ss_lite_csr_rready
		.p0_ss_app_lite_csr_rdata       (),                                                         //  output,   width = 32,                            .p0_ss_app_lite_csr_rdata
		.p0_ss_app_lite_csr_rresp       (),                                                         //  output,    width = 2,                            .p0_ss_app_lite_csr_rresp
		.p0_ss_app_serr                 (dut_p0_ss_app_serr_ss_app_serr),                           //  output,    width = 1,              p0_ss_app_serr.ss_app_serr
		.p0_ss_app_dlup                 (dut_p0_ss_app_dlup_ss_app_dlup),                           //  output,    width = 1,              p0_ss_app_dlup.ss_app_dlup
		.p0_ss_app_linkup               (dut_p0_ss_app_linkup_ss_app_linkup),                       //  output,    width = 1,            p0_ss_app_linkup.ss_app_linkup
		.p0_ss_app_surprise_down_err    (dut_p0_ss_app_surprise_down_err_ss_app_surprise_down_err), //  output,    width = 1, p0_ss_app_surprise_down_err.ss_app_surprise_down_err
		.p0_ss_app_ltssmstate           (),                                                         //  output,    width = 6,        p0_ss_app_ltssmstate.ss_app_ltssmstate
		.p0_app_ss_st_rx_tuser_halt     ()                                                          //   input,    width = 3,  p0_app_ss_st_rx_tuser_halt.app_ss_st_rx_tuser_halt
	);

	system_iopll_0 iopll0 (
		.refclk   (iopll0_refclk_clk),        //   input,  width = 1,  refclk.clk
		.locked   (iopll0_locked_export),     //  output,  width = 1,  locked.export
		.rst      (resetip_ninit_done_reset), //   input,  width = 1,   reset.reset
		.outclk_0 (iopll0_outclk0_clk),       //  output,  width = 1, outclk0.clk
		.outclk_1 (iopll0_outclk1_clk)        //  output,  width = 1, outclk1.clk
	);

	mem0 mem0 (
		.clk        (pio0_pio_master_clk_clk),              //   input,    width = 1,   clk1.clk
		.address    (mm_interconnect_0_mem0_s1_address),    //   input,    width = 8,     s1.address
		.read       (mm_interconnect_0_mem0_s1_read),       //   input,    width = 1,       .read
		.readdata   (mm_interconnect_0_mem0_s1_readdata),   //  output,  width = 512,       .readdata
		.byteenable (mm_interconnect_0_mem0_s1_byteenable), //   input,   width = 64,       .byteenable
		.write      (mm_interconnect_0_mem0_s1_write),      //   input,    width = 1,       .write
		.writedata  (mm_interconnect_0_mem0_s1_writedata),  //   input,  width = 512,       .writedata
		.reset      (~pio0_pio_master_reset_reset)          //   input,    width = 1, reset1.reset
	);

	system_intel_pcie_pio_gts_0 pio0 (
		.Clk_i                        (iopll0_outclk1_clk),                                       //   input,    width = 1,                   axi_st_clk.clk
		.outclk_0                     (iopll0_outclk0_clk),                                       //   input,    width = 1,                 axi_lite_clk.clk
		.coreclkout_hip               (dut_coreclkout_hip_toapp_clk),                             //   input,    width = 1,                          clk.clk
		.Rstn_i                       (dut_p0_reset_status_n_reset),                              //   input,    width = 1,                        reset.reset_n
		.pio_clk                      (pio0_pio_master_clk_clk),                                  //  output,    width = 1,               pio_master_clk.clk
		.pio_rst_n                    (pio0_pio_master_reset_reset),                              //  output,    width = 1,             pio_master_reset.reset_n
		.pio_axi_st_areset_n          (pio0_pio_axi_st_areset_n_reset),                           //  output,    width = 1,          pio_axi_st_areset_n.reset_n
		.pio_axi_lite_areset_n        (pio0_pio_axi_lite_areset_n_reset),                         //  output,    width = 1,        pio_axi_lite_areset_n.reset_n
		.pio_subsystem_cold_rst_n     (pio0_pio_subsystem_cold_rst_n_reset),                      //  output,    width = 1,     pio_subsystem_cold_rst_n.reset_n
		.pio_subsystem_warm_rst_n     (pio0_pio_subsystem_warm_rst_n_reset),                      //  output,    width = 1,     pio_subsystem_warm_rst_n.reset_n
		.ninit_done                   (resetip_ninit_done_reset),                                 //   input,    width = 1,                   ninit_done.reset
		.pio_subsystem_cold_rst_ack_n (dut_p0_subsystem_cold_rst_ack_n_subsystem_cold_rst_ack_n), //   input,    width = 1, pio_subsystem_cold_rst_ack_n.subsystem_cold_rst_ack_n
		.pio_subsystem_warm_rst_ack_n (dut_p0_subsystem_warm_rst_ack_n_subsystem_warm_rst_ack_n), //   input,    width = 1, pio_subsystem_warm_rst_ack_n.subsystem_warm_rst_ack_n
		.pio_initiate_warmrst_req     (dut_p0_initiate_warmrst_req_initiate_warmrst_req),         //   input,    width = 1,     pio_initiate_warmrst_req.initiate_warmrst_req
		.pio_subsystem_rst_rdy        (dut_p0_subsystem_rst_rdy_subsystem_rst_rdy),               //   input,    width = 1,        pio_subsystem_rst_rdy.subsystem_rst_rdy
		.pio_subsystem_rst_req        (pio0_pio_subsystem_rst_req_subsystem_rst_req),             //  output,    width = 1,        pio_subsystem_rst_req.subsystem_rst_req
		.pio_initiate_rst_req_rdy     (pio0_pio_initiate_rst_req_rdy_initiate_rst_req_rdy),       //  output,    width = 1,     pio_initiate_rst_req_rdy.initiate_rst_req_rdy
		.pio_pll_locked               (iopll0_locked_export),                                     //   input,    width = 1,               pio_pll_locked.export
		.pio_address_o                (pio0_pio_master_address),                                  //  output,   width = 64,                   pio_master.address
		.pio_read_o                   (pio0_pio_master_read),                                     //  output,    width = 1,                             .read
		.pio_readdata_i               (pio0_pio_master_readdata),                                 //   input,  width = 512,                             .readdata
		.pio_readdatavalid_i          (pio0_pio_master_readdatavalid),                            //   input,    width = 1,                             .readdatavalid
		.pio_write_o                  (pio0_pio_master_write),                                    //  output,    width = 1,                             .write
		.pio_writedata_o              (pio0_pio_master_writedata),                                //  output,  width = 512,                             .writedata
		.pio_waitrequest_i            (pio0_pio_master_waitrequest),                              //   input,    width = 1,                             .waitrequest
		.pio_byteenable_o             (pio0_pio_master_byteenable),                               //  output,   width = 64,                             .byteenable
		.pio_response_i               (pio0_pio_master_response),                                 //   input,    width = 2,                             .response
		.pio_burstcount_o             (pio0_pio_master_burstcount),                               //  output,    width = 4,                             .burstcount
		.pio_rx_tvalid_i              (dut_p0_st_rx_tvalid),                                      //   input,    width = 1,                       rx_pio.tvalid
		.pio_rx_tready_o              (dut_p0_st_rx_tready),                                      //  output,    width = 1,                             .tready
		.pio_rx_tdata_i               (dut_p0_st_rx_tdata),                                       //   input,  width = 256,                             .tdata
		.pio_rx_tkeep_i               (dut_p0_st_rx_tkeep),                                       //   input,   width = 32,                             .tkeep
		.pio_rx_tlast_i               (dut_p0_st_rx_tlast),                                       //   input,    width = 1,                             .tlast
		.pio_tx_tvalid_o              (pio0_tx_pio_tvalid),                                       //  output,    width = 1,                       tx_pio.tvalid
		.pio_tx_tready_i              (pio0_tx_pio_tready),                                       //   input,    width = 1,                             .tready
		.pio_tx_tdata_o               (pio0_tx_pio_tdata),                                        //  output,  width = 256,                             .tdata
		.pio_tx_tkeep_o               (pio0_tx_pio_tkeep),                                        //  output,   width = 32,                             .tkeep
		.pio_tx_tlast_o               (pio0_tx_pio_tlast),                                        //  output,    width = 1,                             .tlast
		.pio_txcrdt_tvalid            (dut_p0_st_txcrdt_tvalid),                                  //   input,    width = 1,                  tx_crdt_pio.tvalid
		.pio_txcrdt_tdata             (dut_p0_st_txcrdt_tdata),                                   //   input,   width = 19,                             .tdata
		.pio_ctrlshadow_tvalid_i      (dut_p0_st_ctrlshadow_tvalid),                              //   input,    width = 1,               ctrlshadow_pio.tvalid
		.pio_ctrlshadow_tdata_i       (dut_p0_st_ctrlshadow_tdata),                               //   input,   width = 40,                             .tdata
		.pio_cplto_tvalid_i           (dut_p0_st_cplto_tvalid),                                   //   input,    width = 1,                    cplto_pio.tvalid
		.pio_cplto_tdata_i            (dut_p0_st_cplto_tdata)                                     //   input,   width = 30,                             .tdata
	);

	resetIP resetip (
		.ninit_done (resetip_ninit_done_reset)  //  output,  width = 1, ninit_done.reset
	);

	system_intel_srcss_gts_0 srcssip (
		.o_pma_cu_clk (srcssip_o_pma_cu_clk_clk)  //  output,  width = 1, o_pma_cu_clk.clk
	);

	system_intel_systemclk_gts_0 syspll_inst (
		.o_pll_lock  (syspll_inst_o_pll_lock_o_pll_lock), //  output,  width = 1,  o_pll_lock.o_pll_lock
		.o_syspll_c0 (syspll_inst_o_syspll_c0_clk),       //  output,  width = 1, o_syspll_c0.clk
		.i_refclk    (refclk_xcvr_clk)                    //   input,  width = 1, refclk_xcvr.clk
	);

	system_altera_mm_interconnect_1920_ciglmda mm_interconnect_0 (
		.pio0_pio_master_address                                      (pio0_pio_master_address),              //   input,   width = 64,                                        pio0_pio_master.address
		.pio0_pio_master_waitrequest                                  (pio0_pio_master_waitrequest),          //  output,    width = 1,                                                       .waitrequest
		.pio0_pio_master_burstcount                                   (pio0_pio_master_burstcount),           //   input,    width = 4,                                                       .burstcount
		.pio0_pio_master_byteenable                                   (pio0_pio_master_byteenable),           //   input,   width = 64,                                                       .byteenable
		.pio0_pio_master_read                                         (pio0_pio_master_read),                 //   input,    width = 1,                                                       .read
		.pio0_pio_master_readdata                                     (pio0_pio_master_readdata),             //  output,  width = 512,                                                       .readdata
		.pio0_pio_master_readdatavalid                                (pio0_pio_master_readdatavalid),        //  output,    width = 1,                                                       .readdatavalid
		.pio0_pio_master_write                                        (pio0_pio_master_write),                //   input,    width = 1,                                                       .write
		.pio0_pio_master_writedata                                    (pio0_pio_master_writedata),            //   input,  width = 512,                                                       .writedata
		.pio0_pio_master_response                                     (pio0_pio_master_response),             //  output,    width = 2,                                                       .response
		.mem0_s1_address                                              (mm_interconnect_0_mem0_s1_address),    //  output,    width = 8,                                                mem0_s1.address
		.mem0_s1_write                                                (mm_interconnect_0_mem0_s1_write),      //  output,    width = 1,                                                       .write
		.mem0_s1_read                                                 (mm_interconnect_0_mem0_s1_read),       //  output,    width = 1,                                                       .read
		.mem0_s1_readdata                                             (mm_interconnect_0_mem0_s1_readdata),   //   input,  width = 512,                                                       .readdata
		.mem0_s1_writedata                                            (mm_interconnect_0_mem0_s1_writedata),  //  output,  width = 512,                                                       .writedata
		.mem0_s1_byteenable                                           (mm_interconnect_0_mem0_s1_byteenable), //  output,   width = 64,                                                       .byteenable
		.mem0_reset1_reset_bridge_in_reset_reset                      (rst_controller_002_reset_out_reset),   //   input,    width = 1,                      mem0_reset1_reset_bridge_in_reset.reset
		.pio0_pio_master_translator_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),   //   input,    width = 1, pio0_pio_master_translator_reset_reset_bridge_in_reset.reset
		.pio0_pio_master_clk_clk                                      (pio0_pio_master_clk_clk)               //   input,    width = 1,                                    pio0_pio_master_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pio0_pio_axi_st_areset_n_reset), //   input,  width = 1, reset_in0.reset
		.clk            (iopll0_outclk1_clk),              //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset),  //  output,  width = 1, reset_out.reset
		.reset_req      (),                                // (terminated),                       
		.reset_req_in0  (1'b0),                            // (terminated),                       
		.reset_in1      (1'b0),                            // (terminated),                       
		.reset_req_in1  (1'b0),                            // (terminated),                       
		.reset_in2      (1'b0),                            // (terminated),                       
		.reset_req_in2  (1'b0),                            // (terminated),                       
		.reset_in3      (1'b0),                            // (terminated),                       
		.reset_req_in3  (1'b0),                            // (terminated),                       
		.reset_in4      (1'b0),                            // (terminated),                       
		.reset_req_in4  (1'b0),                            // (terminated),                       
		.reset_in5      (1'b0),                            // (terminated),                       
		.reset_req_in5  (1'b0),                            // (terminated),                       
		.reset_in6      (1'b0),                            // (terminated),                       
		.reset_req_in6  (1'b0),                            // (terminated),                       
		.reset_in7      (1'b0),                            // (terminated),                       
		.reset_req_in7  (1'b0),                            // (terminated),                       
		.reset_in8      (1'b0),                            // (terminated),                       
		.reset_req_in8  (1'b0),                            // (terminated),                       
		.reset_in9      (1'b0),                            // (terminated),                       
		.reset_req_in9  (1'b0),                            // (terminated),                       
		.reset_in10     (1'b0),                            // (terminated),                       
		.reset_req_in10 (1'b0),                            // (terminated),                       
		.reset_in11     (1'b0),                            // (terminated),                       
		.reset_req_in11 (1'b0),                            // (terminated),                       
		.reset_in12     (1'b0),                            // (terminated),                       
		.reset_req_in12 (1'b0),                            // (terminated),                       
		.reset_in13     (1'b0),                            // (terminated),                       
		.reset_req_in13 (1'b0),                            // (terminated),                       
		.reset_in14     (1'b0),                            // (terminated),                       
		.reset_req_in14 (1'b0),                            // (terminated),                       
		.reset_in15     (1'b0),                            // (terminated),                       
		.reset_req_in15 (1'b0)                             // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~pio0_pio_axi_lite_areset_n_reset),  //   input,  width = 1, reset_in0.reset
		.clk            (iopll0_outclk0_clk),                 //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("both"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~pio0_pio_master_reset_reset),       //   input,  width = 1, reset_in0.reset
		.clk            (pio0_pio_master_clk_clk),            //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
