// system_intel_pcie_gts_0_intel_pcie_gts_pcie_hal_top_300_un6p7py.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_intel_pcie_gts_0_intel_pcie_gts_pcie_hal_top_300_un6p7py #(
		parameter       ch0_pcs_l_tx_en_atom                                = "FALSE",
		parameter       ch0_pcs_l_rx_en_atom                                = "FALSE",
		parameter       ch0_fec_loopback_mode_atom                          = "CH0_LOOPBACK_MODE_DISABLE",
		parameter       ch0_fec_dyn_tx_mux_atom                             = "CH0_DYN_TX_MUX_ETHPCS",
		parameter       ch0_fec_error_atom                                  = "FALSE",
		parameter       ch0_fec_rx_en_atom                                  = "TRUE",
		parameter       ch0_fec_tx_en_atom                                  = "TRUE",
		parameter       ch0_fec_mode_atom                                   = "CH0_FEC_MODE_RSFEC",
		parameter       ch1_pcs_l_tx_en_atom                                = "FALSE",
		parameter       ch1_pcs_l_rx_en_atom                                = "FALSE",
		parameter       ch1_fec_loopback_mode_atom                          = "CH1_LOOPBACK_MODE_DISABLE",
		parameter       ch1_fec_dyn_tx_mux_atom                             = "CH1_DYN_TX_MUX_UNUSED",
		parameter       ch1_fec_error_atom                                  = "FALSE",
		parameter       ch1_fec_rx_en_atom                                  = "FALSE",
		parameter       ch1_fec_tx_en_atom                                  = "FALSE",
		parameter       ch1_fec_mode_atom                                   = "CH1_FEC_MODE_DISABLED",
		parameter       ch2_pcs_l_tx_en_atom                                = "FALSE",
		parameter       ch2_pcs_l_rx_en_atom                                = "FALSE",
		parameter       ch2_fec_loopback_mode_atom                          = "CH2_LOOPBACK_MODE_DISABLE",
		parameter       ch2_fec_dyn_tx_mux_atom                             = "CH2_DYN_TX_MUX_ETHPCS",
		parameter       ch2_fec_error_atom                                  = "FALSE",
		parameter       ch2_fec_rx_en_atom                                  = "TRUE",
		parameter       ch2_fec_tx_en_atom                                  = "TRUE",
		parameter       ch2_fec_mode_atom                                   = "CH2_FEC_MODE_RSFEC",
		parameter       ch3_pcs_l_tx_en_atom                                = "FALSE",
		parameter       ch3_pcs_l_rx_en_atom                                = "FALSE",
		parameter       ch3_fec_loopback_mode_atom                          = "CH3_LOOPBACK_MODE_DISABLE",
		parameter       ch3_fec_dyn_tx_mux_atom                             = "CH3_DYN_TX_MUX_DESKEW",
		parameter       ch3_fec_error_atom                                  = "FALSE",
		parameter       ch3_fec_rx_en_atom                                  = "TRUE",
		parameter       ch3_fec_tx_en_atom                                  = "TRUE",
		parameter       ch3_fec_mode_atom                                   = "CH3_FEC_MODE_RSFEC",
		parameter       ch0_xcvr_rx_prbs_monitor_en_atom                    = "CH0_RX_PRBS_MONITOR_EN_DISABLE",
		parameter       ch1_xcvr_rx_prbs_monitor_en_atom                    = "CH1_RX_PRBS_MONITOR_EN_ENABLE",
		parameter       ch2_xcvr_rx_prbs_monitor_en_atom                    = "CH2_RX_PRBS_MONITOR_EN_ENABLE",
		parameter       ch3_xcvr_rx_prbs_monitor_en_atom                    = "CH3_RX_PRBS_MONITOR_EN_ENABLE",
		parameter       ch0_tx_prbs_gen_en_atom                             = "CH0_TX_PRBS_GEN_EN_DISABLE",
		parameter       ch1_tx_prbs_gen_en_atom                             = "CH1_TX_PRBS_GEN_EN_DISABLE",
		parameter       ch2_tx_prbs_gen_en_atom                             = "CH2_TX_PRBS_GEN_EN_DISABLE",
		parameter       ch3_tx_prbs_gen_en_atom                             = "CH3_TX_PRBS_GEN_EN_DISABLE",
		parameter       ch0_rx_user1_clk_mux_dynamic_sel_atom               = "CH0_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch0_rx_user2_clk_mux_dynamic_sel_atom               = "CH0_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch0_tx_user1_clk_mux_dynamic_sel_atom               = "CH0_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch0_tx_user2_clk_mux_dynamic_sel_atom               = "CH0_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch1_rx_user1_clk_mux_dynamic_sel_atom               = "CH1_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch1_rx_user2_clk_mux_dynamic_sel_atom               = "CH1_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch1_tx_user1_clk_mux_dynamic_sel_atom               = "CH1_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch1_tx_user2_clk_mux_dynamic_sel_atom               = "CH1_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch2_rx_user1_clk_mux_dynamic_sel_atom               = "CH2_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch2_rx_user2_clk_mux_dynamic_sel_atom               = "CH2_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch2_tx_user1_clk_mux_dynamic_sel_atom               = "CH2_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch2_tx_user2_clk_mux_dynamic_sel_atom               = "CH2_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch3_rx_user1_clk_mux_dynamic_sel_atom               = "CH3_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch3_rx_user2_clk_mux_dynamic_sel_atom               = "CH3_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch3_tx_user1_clk_mux_dynamic_sel_atom               = "CH3_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch3_tx_user2_clk_mux_dynamic_sel_atom               = "CH3_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch0_pcie_mode_atom                                  = "CH0_PCIE_MODE_GEN4",
		parameter       ch1_pcie_mode_atom                                  = "CH1_PCIE_MODE_GEN4",
		parameter       ch2_pcie_mode_atom                                  = "CH2_PCIE_MODE_GEN4",
		parameter       ch3_pcie_mode_atom                                  = "CH3_PCIE_MODE_GEN4",
		parameter       ch0_xcvr_rx_protocol_hint_atom                      = "CH0_RX_PROTOCOL_HINT_DISABLED",
		parameter       ch1_xcvr_rx_protocol_hint_atom                      = "CH1_RX_PROTOCOL_HINT_DISABLED",
		parameter       ch2_xcvr_rx_protocol_hint_atom                      = "CH2_RX_PROTOCOL_HINT_DISABLED",
		parameter       ch3_xcvr_rx_protocol_hint_atom                      = "CH3_RX_PROTOCOL_HINT_DISABLED",
		parameter       ch0_clkrx_refclk_cssm_fw_control_atom               = "CH0_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch1_clkrx_refclk_cssm_fw_control_atom               = "CH1_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch2_clkrx_refclk_cssm_fw_control_atom               = "CH2_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch3_clkrx_refclk_cssm_fw_control_atom               = "CH3_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch0_clkrx_refclk_sector_specifies_refclk_ready_atom = "CH0_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch1_clkrx_refclk_sector_specifies_refclk_ready_atom = "CH1_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch2_clkrx_refclk_sector_specifies_refclk_ready_atom = "CH2_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch3_clkrx_refclk_sector_specifies_refclk_ready_atom = "CH3_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch0_local_refclk_cssm_fw_control_atom               = "CH0_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch1_local_refclk_cssm_fw_control_atom               = "CH1_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch2_local_refclk_cssm_fw_control_atom               = "CH2_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch3_local_refclk_cssm_fw_control_atom               = "CH3_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch0_local_refclk_sector_specifies_refclk_ready_atom = "CH0_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch1_local_refclk_sector_specifies_refclk_ready_atom = "CH1_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch2_local_refclk_sector_specifies_refclk_ready_atom = "CH2_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch3_local_refclk_sector_specifies_refclk_ready_atom = "CH3_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch0_tx_bonding_category_atom                        = "CH0_TX_BONDING_CATEGORY_BONDING_LEADER",
		parameter       ch1_tx_bonding_category_atom                        = "CH1_TX_BONDING_CATEGORY_BONDING_FOLLOWER",
		parameter       ch2_tx_bonding_category_atom                        = "CH2_TX_BONDING_CATEGORY_BONDING_FOLLOWER",
		parameter       ch3_tx_bonding_category_atom                        = "CH3_TX_BONDING_CATEGORY_BONDING_FOLLOWER",
		parameter       hal_num_of_lanes_hwtcl                              = 4,
		parameter       ch0_duplex_mode_atom                                = "CH0_DUPLEX_MODE_DUPLEX",
		parameter       ch0_fec_spec_atom                                   = "CH0_FEC_SPEC_DISABLED",
		parameter       ch0_fracture_atom                                   = "CH0_FRACTURE_UNUSED",
		parameter       ch0_dr_enabled_atom                                 = "CH0_DR_ENABLED_DR_DISABLED",
		parameter       ch0_sup_mode_atom                                   = "CH0_SUP_MODE_USER_MODE",
		parameter       ch0_sim_mode_atom                                   = "CH0_SIM_MODE_DISABLE",
		parameter       ch1_duplex_mode_atom                                = "CH1_DUPLEX_MODE_DUPLEX",
		parameter       ch1_fec_spec_atom                                   = "CH1_FEC_SPEC_DISABLED",
		parameter       ch1_fracture_atom                                   = "CH1_FRACTURE_UNUSED",
		parameter       ch1_dr_enabled_atom                                 = "CH1_DR_ENABLED_DR_DISABLED",
		parameter       ch1_sup_mode_atom                                   = "CH1_SUP_MODE_USER_MODE",
		parameter       ch1_sim_mode_atom                                   = "CH1_SIM_MODE_DISABLE",
		parameter       ch2_duplex_mode_atom                                = "CH2_DUPLEX_MODE_DUPLEX",
		parameter       ch2_fec_spec_atom                                   = "CH2_FEC_SPEC_DISABLED",
		parameter       ch2_fracture_atom                                   = "CH2_FRACTURE_UNUSED",
		parameter       ch2_dr_enabled_atom                                 = "CH2_DR_ENABLED_DR_DISABLED",
		parameter       ch2_sup_mode_atom                                   = "CH2_SUP_MODE_USER_MODE",
		parameter       ch2_sim_mode_atom                                   = "CH2_SIM_MODE_DISABLE",
		parameter       ch3_duplex_mode_atom                                = "CH3_DUPLEX_MODE_DUPLEX",
		parameter       ch3_fec_spec_atom                                   = "CH3_FEC_SPEC_DISABLED",
		parameter       ch3_fracture_atom                                   = "CH3_FRACTURE_UNUSED",
		parameter       ch3_dr_enabled_atom                                 = "CH3_DR_ENABLED_DR_DISABLED",
		parameter       ch3_sup_mode_atom                                   = "CH3_SUP_MODE_USER_MODE",
		parameter       ch3_sim_mode_atom                                   = "CH3_SIM_MODE_DISABLE",
		parameter       ch0_xcvr_tx_preloaded_hardware_configs_atom         = "CH0_TX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch0_xcvr_rx_preloaded_hardware_configs_atom         = "CH0_RX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch0_lc_postdiv_sel_atom                             = "CH0_LC_POSTDIV_SEL_SYNTH2",
		parameter       ch0_sequencer_reg_en_atom                           = "CH0_SEQUENCER_REG_EN_ENABLE",
		parameter       ch0_rst_mux_static_sel_atom                         = "CH0_RST_MUX_STATIC_SEL_HRC",
		parameter[3:0]  ch0_xcvr_tx_prbs_pattern_atom                       = 4'b0000,
		parameter[3:0]  ch0_xcvr_rx_prbs_pattern_atom                       = 4'b0000,
		parameter       ch0_xcvr_tx_user_clk_only_mode_atom                 = "CH0_TX_USER_CLK_ONLY_MODE_DISABLE",
		parameter       ch0_xcvr_tx_width_atom                              = "CH0_TX_WIDTH_X16",
		parameter       ch0_xcvr_rx_width_atom                              = "CH0_RX_WIDTH_X16",
		parameter       ch0_phy_loopback_mode_atom                          = "CH0_LOOPBACK_MODE_DISABLED",
		parameter       ch0_flux_mode_atom                                  = "CH0_FLUX_MODE_FLUX_MODE_BYPASS",
		parameter       ch0_tx_sim_mode_atom                                = "CH0_TX_SIM_MODE_DISABLE",
		parameter       ch0_rx_sim_mode_atom                                = "CH0_RX_SIM_MODE_DISABLE",
		parameter       ch0_tx_dl_enable_atom                               = "CH0_TX_DL_ENABLE_DISABLE",
		parameter       ch0_rx_dl_enable_atom                               = "CH0_RX_DL_ENABLE_ENABLE",
		parameter       ch0_rx_fec_type_used_atom                           = "CH0_RX_FEC_TYPE_USED_RS",
		parameter       ch1_xcvr_tx_preloaded_hardware_configs_atom         = "CH1_TX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch1_xcvr_rx_preloaded_hardware_configs_atom         = "CH1_RX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch1_lc_postdiv_sel_atom                             = "CH1_LC_POSTDIV_SEL_SYNTH2",
		parameter       ch1_sequencer_reg_en_atom                           = "CH1_SEQUENCER_REG_EN_DISABLE",
		parameter       ch1_rst_mux_static_sel_atom                         = "CH1_RST_MUX_STATIC_SEL_HRC",
		parameter[3:0]  ch1_xcvr_tx_prbs_pattern_atom                       = 4'b0000,
		parameter[3:0]  ch1_xcvr_rx_prbs_pattern_atom                       = 4'b0001,
		parameter       ch1_xcvr_tx_user_clk_only_mode_atom                 = "CH1_TX_USER_CLK_ONLY_MODE_DISABLE",
		parameter       ch1_xcvr_tx_width_atom                              = "CH1_TX_WIDTH_X16",
		parameter       ch1_xcvr_rx_width_atom                              = "CH1_RX_WIDTH_X16",
		parameter       ch1_phy_loopback_mode_atom                          = "CH1_LOOPBACK_MODE_DISABLED",
		parameter       ch1_flux_mode_atom                                  = "CH1_FLUX_MODE_FLUX_MODE_BYPASS",
		parameter       ch1_tx_sim_mode_atom                                = "CH1_TX_SIM_MODE_DISABLE",
		parameter       ch1_rx_sim_mode_atom                                = "CH1_RX_SIM_MODE_DISABLE",
		parameter       ch1_tx_dl_enable_atom                               = "CH1_TX_DL_ENABLE_DISABLE",
		parameter       ch1_rx_dl_enable_atom                               = "CH1_RX_DL_ENABLE_ENABLE",
		parameter       ch1_rx_fec_type_used_atom                           = "CH1_RX_FEC_TYPE_USED_NONE",
		parameter       ch2_xcvr_tx_preloaded_hardware_configs_atom         = "CH2_TX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch2_xcvr_rx_preloaded_hardware_configs_atom         = "CH2_RX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch2_lc_postdiv_sel_atom                             = "CH2_LC_POSTDIV_SEL_SYNTH2",
		parameter       ch2_sequencer_reg_en_atom                           = "CH2_SEQUENCER_REG_EN_DISABLE",
		parameter       ch2_rst_mux_static_sel_atom                         = "CH2_RST_MUX_STATIC_SEL_HRC",
		parameter[3:0]  ch2_xcvr_tx_prbs_pattern_atom                       = 4'b0000,
		parameter[3:0]  ch2_xcvr_rx_prbs_pattern_atom                       = 4'b0011,
		parameter       ch2_xcvr_tx_user_clk_only_mode_atom                 = "CH2_TX_USER_CLK_ONLY_MODE_DISABLE",
		parameter       ch2_xcvr_tx_width_atom                              = "CH2_TX_WIDTH_X16",
		parameter       ch2_xcvr_rx_width_atom                              = "CH2_RX_WIDTH_X16",
		parameter       ch2_phy_loopback_mode_atom                          = "CH2_LOOPBACK_MODE_DISABLED",
		parameter       ch2_flux_mode_atom                                  = "CH2_FLUX_MODE_FLUX_MODE_BYPASS",
		parameter       ch2_tx_sim_mode_atom                                = "CH2_TX_SIM_MODE_DISABLE",
		parameter       ch2_rx_sim_mode_atom                                = "CH2_RX_SIM_MODE_DISABLE",
		parameter       ch2_tx_dl_enable_atom                               = "CH2_TX_DL_ENABLE_DISABLE",
		parameter       ch2_rx_dl_enable_atom                               = "CH2_RX_DL_ENABLE_DISABLE",
		parameter       ch2_rx_fec_type_used_atom                           = "CH2_RX_FEC_TYPE_USED_RS",
		parameter       ch3_xcvr_tx_preloaded_hardware_configs_atom         = "CH3_TX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch3_xcvr_rx_preloaded_hardware_configs_atom         = "CH3_RX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch3_lc_postdiv_sel_atom                             = "CH3_LC_POSTDIV_SEL_SYNTH2",
		parameter       ch3_sequencer_reg_en_atom                           = "CH3_SEQUENCER_REG_EN_ENABLE",
		parameter       ch3_rst_mux_static_sel_atom                         = "CH3_RST_MUX_STATIC_SEL_HRC",
		parameter[3:0]  ch3_xcvr_tx_prbs_pattern_atom                       = 4'b0000,
		parameter[3:0]  ch3_xcvr_rx_prbs_pattern_atom                       = 4'b0111,
		parameter       ch3_xcvr_tx_user_clk_only_mode_atom                 = "CH3_TX_USER_CLK_ONLY_MODE_DISABLE",
		parameter       ch3_xcvr_tx_width_atom                              = "CH3_TX_WIDTH_X16",
		parameter       ch3_xcvr_rx_width_atom                              = "CH3_RX_WIDTH_X16",
		parameter       ch3_phy_loopback_mode_atom                          = "CH3_LOOPBACK_MODE_DISABLED",
		parameter       ch3_flux_mode_atom                                  = "CH3_FLUX_MODE_FLUX_MODE_BYPASS",
		parameter       ch3_tx_sim_mode_atom                                = "CH3_TX_SIM_MODE_DISABLE",
		parameter       ch3_rx_sim_mode_atom                                = "CH3_RX_SIM_MODE_DISABLE",
		parameter       ch3_tx_dl_enable_atom                               = "CH3_TX_DL_ENABLE_DISABLE",
		parameter       ch3_rx_dl_enable_atom                               = "CH3_RX_DL_ENABLE_ENABLE",
		parameter       ch3_rx_fec_type_used_atom                           = "CH3_RX_FEC_TYPE_USED_RS",
		parameter[5:0]  ch0_tx_pll_l_counter_atom                           = 6'b000001,
		parameter[5:0]  ch0_cdr_l_counter_atom                              = 6'b000001,
		parameter       ch0_tx_pll_refclk_select_atom                       = "CH0_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter       ch0_cdr_refclk_select_atom                          = "CH0_CDR_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter[5:0]  ch1_tx_pll_l_counter_atom                           = 6'b000001,
		parameter[5:0]  ch1_cdr_l_counter_atom                              = 6'b000001,
		parameter       ch1_tx_pll_refclk_select_atom                       = "CH1_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter       ch1_cdr_refclk_select_atom                          = "CH1_CDR_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter[5:0]  ch2_tx_pll_l_counter_atom                           = 6'b000001,
		parameter[5:0]  ch2_cdr_l_counter_atom                              = 6'b000001,
		parameter       ch2_tx_pll_refclk_select_atom                       = "CH2_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter       ch2_cdr_refclk_select_atom                          = "CH2_CDR_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter[5:0]  ch3_tx_pll_l_counter_atom                           = 6'b000001,
		parameter[5:0]  ch3_cdr_l_counter_atom                              = 6'b000001,
		parameter       ch3_tx_pll_refclk_select_atom                       = "CH3_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter       ch3_cdr_refclk_select_atom                          = "CH3_CDR_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter[17:0] ch0_rx_dl_rx_lat_bit_for_async_atom                 = 18'b010100000100010011,
		parameter       ch0_rx_dl_rxbit_cntr_pma_atom                       = "CH0_RX_DL_RXBIT_CNTR_PMA_DISABLE",
		parameter[17:0] ch0_rx_dl_rxbit_rollover_atom                       = 18'b111110100100001111,
		parameter[17:0] ch1_rx_dl_rx_lat_bit_for_async_atom                 = 18'b111110100110100101,
		parameter       ch1_rx_dl_rxbit_cntr_pma_atom                       = "CH1_RX_DL_RXBIT_CNTR_PMA_ENABLE",
		parameter[17:0] ch1_rx_dl_rxbit_rollover_atom                       = 18'b001001111001000101,
		parameter[17:0] ch2_rx_dl_rx_lat_bit_for_async_atom                 = 18'b111010100000111101,
		parameter       ch2_rx_dl_rxbit_cntr_pma_atom                       = "CH2_RX_DL_RXBIT_CNTR_PMA_DISABLE",
		parameter[17:0] ch2_rx_dl_rxbit_rollover_atom                       = 18'b111000111110011110,
		parameter[17:0] ch3_rx_dl_rx_lat_bit_for_async_atom                 = 18'b100000100111100001,
		parameter       ch3_rx_dl_rxbit_cntr_pma_atom                       = "CH3_RX_DL_RXBIT_CNTR_PMA_DISABLE",
		parameter[17:0] ch3_rx_dl_rxbit_rollover_atom                       = 18'b001101111001101011,
		parameter       ch0_tx_bond_size_atom                               = "CH0_TX_BOND_SIZE_X4",
		parameter       ch1_tx_bond_size_atom                               = "CH1_TX_BOND_SIZE_X4",
		parameter       ch2_tx_bond_size_atom                               = "CH2_TX_BOND_SIZE_X4",
		parameter       ch3_tx_bond_size_atom                               = "CH3_TX_BOND_SIZE_X4",
		parameter       pcie_parity_bypass                                  = "true",
		parameter       rxbuf_limit_bypass                                  = 7,
		parameter       maxpayload_size                                     = "MAXPAYLOAD_SIZE_MAX_PAYLOAD_512",
		parameter       pldclk_rate                                         = "PLDCLK_RATE_FAST",
		parameter       port_type                                           = "PORT_TYPE_NATIVE_EP",
		parameter       sris_enable                                         = "SRIS_ENABLE_DISABLED",
		parameter       sris_mode                                           = "false",
		parameter       sim_mode                                            = "SIM_MODE_DISABLE_VSIM_MODE",
		parameter       sup_mode                                            = "SUP_MODE_USER_MODE",
		parameter       cvp_enable                                          = "CVP_ENABLE_DISABLED",
		parameter       cii_monitor_en                                      = "CII_MONITOR_EN_DISABLE",
		parameter[31:0] pclk_clk_hz                                         = 32'b00111011100110101100101000000000,
		parameter       pf0_cap_link_surprise_down_err_cap                  = "PF0_CAP_LINK_SURPRISE_DOWN_ERR_CAP_DISABLE",
		parameter[31:0] sys_clk_hz                                          = 32'b00010100110111001001001110000000,
		parameter       link_rate                                           = "LINK_RATE_GEN4",
		parameter       link_width                                          = "LINK_WIDTH_X4",
		parameter       num_of_lanes                                        = "NUM_OF_LANES_NUM_4",
		parameter       pf0_dsp_16g_tx_preset0                              = 7,
		parameter       pf0_dsp_16g_tx_preset1                              = 7,
		parameter       pf0_dsp_16g_tx_preset2                              = 7,
		parameter       pf0_dsp_16g_tx_preset3                              = 7,
		parameter       pf0_dsp_16g_tx_preset4                              = 0,
		parameter       pf0_dsp_16g_tx_preset5                              = 0,
		parameter       pf0_dsp_16g_tx_preset6                              = 0,
		parameter       pf0_dsp_16g_tx_preset7                              = 0,
		parameter       pf0_dsp_16g_tx_preset8                              = 0,
		parameter       pf0_dsp_16g_tx_preset9                              = 0,
		parameter       pf0_dsp_16g_tx_preset10                             = 0,
		parameter       pf0_dsp_16g_tx_preset11                             = 0,
		parameter       pf0_dsp_16g_tx_preset12                             = 0,
		parameter       pf0_dsp_16g_tx_preset13                             = 0,
		parameter       pf0_dsp_16g_tx_preset14                             = 0,
		parameter       pf0_dsp_16g_tx_preset15                             = 0,
		parameter       pf0_dsp_tx_preset0                                  = 9,
		parameter       pf0_dsp_tx_preset1                                  = 9,
		parameter       pf0_dsp_tx_preset2                                  = 9,
		parameter       pf0_dsp_tx_preset3                                  = 9,
		parameter       pf0_dsp_tx_preset4                                  = 0,
		parameter       pf0_dsp_tx_preset5                                  = 0,
		parameter       pf0_dsp_tx_preset6                                  = 0,
		parameter       pf0_dsp_tx_preset7                                  = 0,
		parameter       pf0_dsp_tx_preset8                                  = 0,
		parameter       pf0_dsp_tx_preset9                                  = 0,
		parameter       pf0_dsp_tx_preset10                                 = 0,
		parameter       pf0_dsp_tx_preset11                                 = 0,
		parameter       pf0_dsp_tx_preset12                                 = 0,
		parameter       pf0_dsp_tx_preset13                                 = 0,
		parameter       pf0_dsp_tx_preset14                                 = 0,
		parameter       pf0_dsp_tx_preset15                                 = 0,
		parameter       pf0_usp_16g_tx_preset0                              = 7,
		parameter       pf0_usp_16g_tx_preset1                              = 7,
		parameter       pf0_usp_16g_tx_preset2                              = 7,
		parameter       pf0_usp_16g_tx_preset3                              = 7,
		parameter       pf0_usp_16g_tx_preset4                              = 0,
		parameter       pf0_usp_16g_tx_preset5                              = 0,
		parameter       pf0_usp_16g_tx_preset6                              = 0,
		parameter       pf0_usp_16g_tx_preset7                              = 0,
		parameter       pf0_usp_16g_tx_preset8                              = 0,
		parameter       pf0_usp_16g_tx_preset9                              = 0,
		parameter       pf0_usp_16g_tx_preset10                             = 0,
		parameter       pf0_usp_16g_tx_preset11                             = 0,
		parameter       pf0_usp_16g_tx_preset12                             = 0,
		parameter       pf0_usp_16g_tx_preset13                             = 0,
		parameter       pf0_usp_16g_tx_preset14                             = 0,
		parameter       pf0_usp_16g_tx_preset15                             = 0,
		parameter       pf0_usp_tx_preset0                                  = 9,
		parameter       pf0_usp_tx_preset1                                  = 9,
		parameter       pf0_usp_tx_preset2                                  = 9,
		parameter       pf0_usp_tx_preset3                                  = 9,
		parameter       pf0_usp_tx_preset4                                  = 0,
		parameter       pf0_usp_tx_preset5                                  = 0,
		parameter       pf0_usp_tx_preset6                                  = 0,
		parameter       pf0_usp_tx_preset7                                  = 0,
		parameter       pf0_usp_tx_preset8                                  = 0,
		parameter       pf0_usp_tx_preset9                                  = 0,
		parameter       pf0_usp_tx_preset10                                 = 0,
		parameter       pf0_usp_tx_preset11                                 = 0,
		parameter       pf0_usp_tx_preset12                                 = 0,
		parameter       pf0_usp_tx_preset13                                 = 0,
		parameter       pf0_usp_tx_preset14                                 = 0,
		parameter       pf0_usp_tx_preset15                                 = 0,
		parameter       pf0_pci_type0_bar0_enabled                          = "PF0_PCI_TYPE0_BAR0_ENABLED_ENABLED",
		parameter[31:0] pf0_pci_type0_bar0_mask_31_1                        = 32'b00000000000000000111111111111111,
		parameter       pf0_bar0_prefetch                                   = "true",
		parameter       pf0_bar0_type                                       = "PF0_BAR0_TYPE_BAR_MEM64",
		parameter       pf0_pci_type0_bar1_enabled                          = "PF0_PCI_TYPE0_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf0_pci_type0_bar1_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf0_bar1_prefetch                                   = "false",
		parameter       pf0_pci_type0_bar2_enabled                          = "PF0_PCI_TYPE0_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf0_pci_type0_bar2_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf0_bar2_prefetch                                   = "false",
		parameter       pf0_bar2_type                                       = "PF0_BAR2_TYPE_BAR_MEM32",
		parameter       pf0_pci_type0_bar3_enabled                          = "PF0_PCI_TYPE0_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf0_pci_type0_bar3_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf0_bar3_prefetch                                   = "false",
		parameter       pf0_pci_type0_bar4_enabled                          = "PF0_PCI_TYPE0_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf0_pci_type0_bar4_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf0_bar4_prefetch                                   = "false",
		parameter       pf0_bar4_type                                       = "PF0_BAR4_TYPE_BAR_MEM32",
		parameter       pf0_pci_type0_bar5_enabled                          = "PF0_PCI_TYPE0_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf0_pci_type0_bar5_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf0_bar5_prefetch                                   = "false",
		parameter       pf0_rom_bar_enable                                  = "PF0_ROM_BAR_ENABLE_DISABLED",
		parameter       pf0_rom_mask                                        = 0,
		parameter       pf0_rom_bar_enabled                                 = "PF0_ROM_BAR_ENABLED_DISABLED",
		parameter       pf0_rp_rom_bar_enabled                              = "PF0_RP_ROM_BAR_ENABLED_DISABLED",
		parameter       pf0_rp_rom_mask                                     = 0,
		parameter       pf0_sriov_vf_bar0_enabled                           = "PF0_SRIOV_VF_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf0_sriov_vf_bar0_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf0_sriov_vf_bar0_prefetch                          = "false",
		parameter       pf0_sriov_vf_bar0_type                              = "PF0_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf0_sriov_vf_bar1_enabled                           = "PF0_SRIOV_VF_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf0_sriov_vf_bar1_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf0_sriov_vf_bar1_prefetch                          = "false",
		parameter       pf0_sriov_vf_bar2_enabled                           = "PF0_SRIOV_VF_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf0_sriov_vf_bar2_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf0_sriov_vf_bar2_prefetch                          = "false",
		parameter       pf0_sriov_vf_bar2_type                              = "PF0_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf0_sriov_vf_bar3_enabled                           = "PF0_SRIOV_VF_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf0_sriov_vf_bar3_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf0_sriov_vf_bar3_prefetch                          = "false",
		parameter       pf0_sriov_vf_bar4_enabled                           = "PF0_SRIOV_VF_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf0_sriov_vf_bar4_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf0_sriov_vf_bar4_prefetch                          = "false",
		parameter       pf0_sriov_vf_bar4_type                              = "PF0_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf0_sriov_vf_bar5_enabled                           = "PF0_SRIOV_VF_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf0_sriov_vf_bar5_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf0_sriov_vf_bar5_prefetch                          = "false",
		parameter       pf1_pci_type0_bar0_enabled                          = "PF1_PCI_TYPE0_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf1_pci_type0_bar0_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf1_bar0_prefetch                                   = "false",
		parameter       pf1_bar0_type                                       = "PF1_BAR0_TYPE_BAR_MEM32",
		parameter       pf1_pci_type0_bar1_enabled                          = "PF1_PCI_TYPE0_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf1_pci_type0_bar1_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf1_bar1_prefetch                                   = "false",
		parameter       pf1_pci_type0_bar2_enabled                          = "PF1_PCI_TYPE0_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf1_pci_type0_bar2_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf1_bar2_prefetch                                   = "false",
		parameter       pf1_bar2_type                                       = "PF1_BAR2_TYPE_BAR_MEM32",
		parameter       pf1_pci_type0_bar3_enabled                          = "PF1_PCI_TYPE0_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf1_pci_type0_bar3_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf1_bar3_prefetch                                   = "false",
		parameter       pf1_pci_type0_bar4_enabled                          = "PF1_PCI_TYPE0_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf1_pci_type0_bar4_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf1_bar4_prefetch                                   = "false",
		parameter       pf1_bar4_type                                       = "PF1_BAR4_TYPE_BAR_MEM32",
		parameter       pf1_pci_type0_bar5_enabled                          = "PF1_PCI_TYPE0_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf1_pci_type0_bar5_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf1_bar5_prefetch                                   = "false",
		parameter       pf1_rom_bar_enable                                  = "PF1_ROM_BAR_ENABLE_DISABLED",
		parameter       pf1_rom_mask                                        = 0,
		parameter       pf1_rom_bar_enabled                                 = "PF1_ROM_BAR_ENABLED_DISABLED",
		parameter       pf1_sriov_vf_bar0_enabled                           = "PF1_SRIOV_VF_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf1_sriov_vf_bar0_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf1_sriov_vf_bar0_prefetch                          = "false",
		parameter       pf1_sriov_vf_bar0_type                              = "PF1_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf1_sriov_vf_bar1_enabled                           = "PF1_SRIOV_VF_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf1_sriov_vf_bar1_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf1_sriov_vf_bar1_prefetch                          = "false",
		parameter       pf1_sriov_vf_bar2_enabled                           = "PF1_SRIOV_VF_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf1_sriov_vf_bar2_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf1_sriov_vf_bar2_prefetch                          = "false",
		parameter       pf1_sriov_vf_bar2_type                              = "PF1_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf1_sriov_vf_bar3_enabled                           = "PF1_SRIOV_VF_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf1_sriov_vf_bar3_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf1_sriov_vf_bar3_prefetch                          = "false",
		parameter       pf1_sriov_vf_bar4_enabled                           = "PF1_SRIOV_VF_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf1_sriov_vf_bar4_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf1_sriov_vf_bar4_prefetch                          = "false",
		parameter       pf1_sriov_vf_bar4_type                              = "PF1_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf1_sriov_vf_bar5_enabled                           = "PF1_SRIOV_VF_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf1_sriov_vf_bar5_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf1_sriov_vf_bar5_prefetch                          = "false",
		parameter       pf2_pci_type0_bar0_enabled                          = "PF2_PCI_TYPE0_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf2_pci_type0_bar0_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf2_bar0_prefetch                                   = "false",
		parameter       pf2_bar0_type                                       = "PF2_BAR0_TYPE_BAR_MEM32",
		parameter       pf2_pci_type0_bar1_enabled                          = "PF2_PCI_TYPE0_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf2_pci_type0_bar1_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf2_bar1_prefetch                                   = "false",
		parameter       pf2_pci_type0_bar2_enabled                          = "PF2_PCI_TYPE0_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf2_pci_type0_bar2_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf2_bar2_prefetch                                   = "false",
		parameter       pf2_bar2_type                                       = "PF2_BAR2_TYPE_BAR_MEM32",
		parameter       pf2_pci_type0_bar3_enabled                          = "PF2_PCI_TYPE0_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf2_pci_type0_bar3_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf2_bar3_prefetch                                   = "false",
		parameter       pf2_pci_type0_bar4_enabled                          = "PF2_PCI_TYPE0_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf2_pci_type0_bar4_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf2_bar4_prefetch                                   = "false",
		parameter       pf2_bar4_type                                       = "PF2_BAR4_TYPE_BAR_MEM32",
		parameter       pf2_pci_type0_bar5_enabled                          = "PF2_PCI_TYPE0_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf2_pci_type0_bar5_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf2_bar5_prefetch                                   = "false",
		parameter       pf2_rom_bar_enable                                  = "PF2_ROM_BAR_ENABLE_DISABLED",
		parameter       pf2_rom_mask                                        = 0,
		parameter       pf2_rom_bar_enabled                                 = "PF2_ROM_BAR_ENABLED_DISABLED",
		parameter       pf2_sriov_vf_bar0_enabled                           = "PF2_SRIOV_VF_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf2_sriov_vf_bar0_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf2_sriov_vf_bar0_prefetch                          = "false",
		parameter       pf2_sriov_vf_bar0_type                              = "PF2_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf2_sriov_vf_bar1_enabled                           = "PF2_SRIOV_VF_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf2_sriov_vf_bar1_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf2_sriov_vf_bar1_prefetch                          = "false",
		parameter       pf2_sriov_vf_bar2_enabled                           = "PF2_SRIOV_VF_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf2_sriov_vf_bar2_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf2_sriov_vf_bar2_prefetch                          = "false",
		parameter       pf2_sriov_vf_bar2_type                              = "PF2_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf2_sriov_vf_bar3_enabled                           = "PF2_SRIOV_VF_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf2_sriov_vf_bar3_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf2_sriov_vf_bar3_prefetch                          = "false",
		parameter       pf2_sriov_vf_bar4_enabled                           = "PF2_SRIOV_VF_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf2_sriov_vf_bar4_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf2_sriov_vf_bar4_prefetch                          = "false",
		parameter       pf2_sriov_vf_bar4_type                              = "PF2_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf2_sriov_vf_bar5_enabled                           = "PF2_SRIOV_VF_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf2_sriov_vf_bar5_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf2_sriov_vf_bar5_prefetch                          = "false",
		parameter       pf3_pci_type0_bar0_enabled                          = "PF3_PCI_TYPE0_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf3_pci_type0_bar0_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf3_bar0_prefetch                                   = "false",
		parameter       pf3_bar0_type                                       = "PF3_BAR0_TYPE_BAR_MEM32",
		parameter       pf3_pci_type0_bar1_enabled                          = "PF3_PCI_TYPE0_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf3_pci_type0_bar1_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf3_bar1_prefetch                                   = "false",
		parameter       pf3_pci_type0_bar2_enabled                          = "PF3_PCI_TYPE0_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf3_pci_type0_bar2_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf3_bar2_prefetch                                   = "false",
		parameter       pf3_bar2_type                                       = "PF3_BAR2_TYPE_BAR_MEM32",
		parameter       pf3_pci_type0_bar3_enabled                          = "PF3_PCI_TYPE0_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf3_pci_type0_bar3_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf3_bar3_prefetch                                   = "false",
		parameter       pf3_pci_type0_bar4_enabled                          = "PF3_PCI_TYPE0_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf3_pci_type0_bar4_mask_31_1                        = 32'b00000000000000000000000000000000,
		parameter       pf3_bar4_prefetch                                   = "false",
		parameter       pf3_bar4_type                                       = "PF3_BAR4_TYPE_BAR_MEM32",
		parameter       pf3_pci_type0_bar5_enabled                          = "PF3_PCI_TYPE0_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf3_pci_type0_bar5_mask_31_0                        = 32'b00000000000000000000000000000000,
		parameter       pf3_bar5_prefetch                                   = "false",
		parameter       pf3_rom_bar_enable                                  = "PF3_ROM_BAR_ENABLE_DISABLED",
		parameter       pf3_rom_mask                                        = 0,
		parameter       pf3_rom_bar_enabled                                 = "PF3_ROM_BAR_ENABLED_DISABLED",
		parameter       pf3_sriov_vf_bar0_enabled                           = "PF3_SRIOV_VF_BAR0_ENABLED_DISABLED",
		parameter[31:0] pf3_sriov_vf_bar0_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf3_sriov_vf_bar0_prefetch                          = "false",
		parameter       pf3_sriov_vf_bar0_type                              = "PF3_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf3_sriov_vf_bar1_enabled                           = "PF3_SRIOV_VF_BAR1_ENABLED_DISABLED",
		parameter[31:0] pf3_sriov_vf_bar1_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf3_sriov_vf_bar1_prefetch                          = "false",
		parameter       pf3_sriov_vf_bar2_enabled                           = "PF3_SRIOV_VF_BAR2_ENABLED_DISABLED",
		parameter[31:0] pf3_sriov_vf_bar2_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf3_sriov_vf_bar2_prefetch                          = "false",
		parameter       pf3_sriov_vf_bar2_type                              = "PF3_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf3_sriov_vf_bar3_enabled                           = "PF3_SRIOV_VF_BAR3_ENABLED_DISABLED",
		parameter[31:0] pf3_sriov_vf_bar3_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf3_sriov_vf_bar3_prefetch                          = "false",
		parameter       pf3_sriov_vf_bar4_enabled                           = "PF3_SRIOV_VF_BAR4_ENABLED_DISABLED",
		parameter[31:0] pf3_sriov_vf_bar4_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf3_sriov_vf_bar4_prefetch                          = "false",
		parameter       pf3_sriov_vf_bar4_type                              = "PF3_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32",
		parameter       pf3_sriov_vf_bar5_enabled                           = "PF3_SRIOV_VF_BAR5_ENABLED_DISABLED",
		parameter[31:0] pf3_sriov_vf_bar5_mask                              = 32'b00000000000000000000000000000000,
		parameter       pf3_sriov_vf_bar5_prefetch                          = "false",
		parameter       pf1_enable                                          = "PF1_ENABLE_DISABLED",
		parameter       pf2_enable                                          = "PF2_ENABLE_DISABLED",
		parameter       pf3_enable                                          = "PF3_ENABLE_DISABLED",
		parameter       pf0_sriov_enable                                    = "PF0_SRIOV_ENABLE_DISABLED",
		parameter       pf1_sriov_enable                                    = "PF1_SRIOV_ENABLE_DISABLED",
		parameter       pf2_sriov_enable                                    = "PF2_SRIOV_ENABLE_DISABLED",
		parameter       pf3_sriov_enable                                    = "PF3_SRIOV_ENABLE_DISABLED",
		parameter       pf0_sriov_cap_sup_page_size                         = 0,
		parameter       pf1_sriov_cap_sup_page_size                         = 0,
		parameter       pf2_sriov_cap_sup_page_size                         = 0,
		parameter       pf3_sriov_cap_sup_page_size                         = 0,
		parameter       pf0_sriov_num_vf                                    = 0,
		parameter       pf1_sriov_num_vf                                    = 0,
		parameter       pf2_sriov_num_vf                                    = 0,
		parameter       pf3_sriov_num_vf                                    = 0,
		parameter       pf0_msi_enable                                      = "PF0_MSI_ENABLE_ENABLED",
		parameter       pf0_pci_msi_ext_data_cap                            = "false",
		parameter       pf0_pci_msi_ext_data_en                             = "false",
		parameter       pf0_pci_msi_64_bit_addr_cap                         = "false",
		parameter       pf0_pci_msi_multiple_msg_cap                        = "PF0_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1",
		parameter       pf0_msix_enable                                     = "PF0_MSIX_ENABLE_DISABLED",
		parameter       pf0_pci_msix_table_size                             = 0,
		parameter       pf0_pci_msix_table_offset                           = 0,
		parameter       pf0_pci_msix_bir                                    = 0,
		parameter       pf0_pci_msix_pba                                    = 0,
		parameter       pf0_pci_msix_pba_offset                             = 0,
		parameter       pf0_pci_msix_table_size_vfcomm_cs2                  = 0,
		parameter       pf0_exvf_msix_cap_enable                            = "PF0_EXVF_MSIX_CAP_ENABLE_DISABLED",
		parameter       exvf_msix_tablesize_pf0                             = 0,
		parameter       exvf_msixtable_offset_pf0                           = 0,
		parameter       exvf_msixtable_bir_pf0                              = 0,
		parameter       exvf_msixpba_offset_pf0                             = 0,
		parameter       exvf_msixpba_bir_pf0                                = 0,
		parameter       pf1_msi_enable                                      = "PF1_MSI_ENABLE_DISABLED",
		parameter       pf1_pci_msi_ext_data_cap                            = "false",
		parameter       pf1_pci_msi_ext_data_en                             = "false",
		parameter       pf1_pci_msi_64_bit_addr_cap                         = "false",
		parameter       pf1_pci_msi_multiple_msg_cap                        = "PF1_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1",
		parameter       pf1_msix_enable                                     = "PF1_MSIX_ENABLE_DISABLED",
		parameter       pf1_pci_msix_table_size                             = 0,
		parameter       pf1_pci_msix_table_offset                           = 0,
		parameter       pf1_pci_msix_bir                                    = 0,
		parameter       pf1_pci_msix_pba                                    = 0,
		parameter       pf1_pci_msix_pba_offset                             = 0,
		parameter       pf1_pci_msix_table_size_vfcomm_cs2                  = 0,
		parameter       pf1_exvf_msix_cap_enable                            = "PF1_EXVF_MSIX_CAP_ENABLE_DISABLED",
		parameter       exvf_msix_tablesize_pf1                             = 0,
		parameter       exvf_msixtable_offset_pf1                           = 0,
		parameter       exvf_msixtable_bir_pf1                              = 0,
		parameter       exvf_msixpba_offset_pf1                             = 0,
		parameter       exvf_msixpba_bir_pf1                                = 0,
		parameter       pf2_msi_enable                                      = "PF2_MSI_ENABLE_DISABLED",
		parameter       pf2_pci_msi_ext_data_cap                            = "false",
		parameter       pf2_pci_msi_ext_data_en                             = "false",
		parameter       pf2_pci_msi_64_bit_addr_cap                         = "false",
		parameter       pf2_pci_msi_multiple_msg_cap                        = "PF2_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1",
		parameter       pf2_msix_enable                                     = "PF2_MSIX_ENABLE_DISABLED",
		parameter       pf2_pci_msix_bir                                    = 0,
		parameter       pf2_pci_msix_pba                                    = 0,
		parameter       pf2_pci_msix_pba_offset                             = 0,
		parameter       pf2_pci_msix_table_offset                           = 0,
		parameter       pf2_pci_msix_table_size                             = 0,
		parameter       pf2_pci_msix_table_size_vfcomm_cs2                  = 0,
		parameter       pf2_exvf_msix_cap_enable                            = "PF2_EXVF_MSIX_CAP_ENABLE_DISABLED",
		parameter       exvf_msix_tablesize_pf2                             = 0,
		parameter       exvf_msixtable_offset_pf2                           = 0,
		parameter       exvf_msixtable_bir_pf2                              = 0,
		parameter       exvf_msixpba_offset_pf2                             = 0,
		parameter       exvf_msixpba_bir_pf2                                = 0,
		parameter       pf3_msi_enable                                      = "PF3_MSI_ENABLE_DISABLED",
		parameter       pf3_pci_msi_ext_data_cap                            = "false",
		parameter       pf3_pci_msi_ext_data_en                             = "false",
		parameter       pf3_pci_msi_64_bit_addr_cap                         = "false",
		parameter       pf3_pci_msi_multiple_msg_cap                        = "PF3_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1",
		parameter       pf3_msix_enable                                     = "PF3_MSIX_ENABLE_DISABLED",
		parameter       pf3_pci_msix_bir                                    = 0,
		parameter       pf3_pci_msix_pba                                    = 0,
		parameter       pf3_pci_msix_pba_offset                             = 0,
		parameter       pf3_pci_msix_table_offset                           = 0,
		parameter       pf3_pci_msix_table_size                             = 0,
		parameter       pf3_pci_msix_table_size_vfcomm_cs2                  = 0,
		parameter       pf3_exvf_msix_cap_enable                            = "PF3_EXVF_MSIX_CAP_ENABLE_DISABLED",
		parameter       exvf_msix_tablesize_pf3                             = 0,
		parameter       exvf_msixtable_offset_pf3                           = 0,
		parameter       exvf_msixtable_bir_pf3                              = 0,
		parameter       exvf_msixpba_offset_pf3                             = 0,
		parameter       exvf_msixpba_bir_pf3                                = 0,
		parameter       pf0_prs_ext_cap_enable                              = "PF0_PRS_EXT_CAP_ENABLE_DISABLED",
		parameter       pf0_prs_ext_cap_outstanding_capacity                = 0,
		parameter       pf1_prs_ext_cap_enable                              = "PF1_PRS_EXT_CAP_ENABLE_DISABLED",
		parameter       pf1_prs_ext_cap_outstanding_capacity                = 0,
		parameter       pf2_prs_ext_cap_enable                              = "PF2_PRS_EXT_CAP_ENABLE_DISABLED",
		parameter       pf2_prs_ext_cap_outstanding_capacity                = 0,
		parameter       pf3_prs_ext_cap_enable                              = "PF3_PRS_EXT_CAP_ENABLE_DISABLED",
		parameter       pf3_prs_ext_cap_outstanding_capacity                = 0,
		parameter       pf0_pasid_cap_enable                                = "PF0_PASID_CAP_ENABLE_DISABLED",
		parameter       pf0_pasid_cap_execute_permission_supported          = "PF0_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED",
		parameter       pf0_pasid_cap_max_pasid_width                       = 0,
		parameter       pf0_pasid_cap_privileged_mode_supported             = "PF0_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED",
		parameter       pf1_pasid_cap_enable                                = "PF1_PASID_CAP_ENABLE_DISABLED",
		parameter       pf1_pasid_cap_execute_permission_supported          = "PF1_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED",
		parameter       pf1_pasid_cap_max_pasid_width                       = 0,
		parameter       pf1_pasid_cap_privileged_mode_supported             = "PF1_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED",
		parameter       pf2_pasid_cap_enable                                = "PF2_PASID_CAP_ENABLE_DISABLED",
		parameter       pf2_pasid_cap_execute_permission_supported          = "PF2_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED",
		parameter       pf2_pasid_cap_max_pasid_width                       = 0,
		parameter       pf2_pasid_cap_privileged_mode_supported             = "PF2_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED",
		parameter       pf3_pasid_cap_enable                                = "PF3_PASID_CAP_ENABLE_DISABLED",
		parameter       pf3_pasid_cap_execute_permission_supported          = "PF3_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED",
		parameter       pf3_pasid_cap_max_pasid_width                       = 0,
		parameter       pf3_pasid_cap_privileged_mode_supported             = "PF3_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED",
		parameter       pf0_sn_cap_enable                                   = "PF0_SN_CAP_ENABLE_DISABLED",
		parameter[31:0] pf0_sn_ser_num_reg_1_dw                             = 32'b00000000000000000000000000000000,
		parameter[31:0] pf0_sn_ser_num_reg_2_dw                             = 32'b00000000000000000000000000000000,
		parameter       pf1_sn_cap_enable                                   = "PF1_SN_CAP_ENABLE_DISABLED",
		parameter[31:0] pf1_sn_ser_num_reg_1_dw                             = 32'b00000000000000000000000000000000,
		parameter[31:0] pf1_sn_ser_num_reg_2_dw                             = 32'b00000000000000000000000000000000,
		parameter       pf2_sn_cap_enable                                   = "PF2_SN_CAP_ENABLE_DISABLED",
		parameter[31:0] pf2_sn_ser_num_reg_1_dw                             = 32'b00000000000000000000000000000000,
		parameter[31:0] pf2_sn_ser_num_reg_2_dw                             = 32'b00000000000000000000000000000000,
		parameter       pf3_sn_cap_enable                                   = "PF3_SN_CAP_ENABLE_DISABLED",
		parameter[31:0] pf3_sn_ser_num_reg_1_dw                             = 32'b00000000000000000000000000000000,
		parameter[31:0] pf3_sn_ser_num_reg_2_dw                             = 32'b00000000000000000000000000000000,
		parameter       pf0_pcie_cap_ep_l0s_accpt_latency                   = 0,
		parameter       pf0_pcie_cap_ep_l1_accpt_latency                    = 0,
		parameter       pf0_pcie_cap_l0s_exit_latency_commclk_dis           = 0,
		parameter       pf0_pcie_cap_l1_exit_latency_commclk_dis            = 0,
		parameter       pf1_pcie_cap_ep_l0s_accpt_latency                   = 0,
		parameter       pf1_pcie_cap_ep_l1_accpt_latency                    = 0,
		parameter       pf1_pcie_cap_l0s_exit_latency_commclk_dis           = 0,
		parameter       pf1_pcie_cap_l1_exit_latency_commclk_dis            = 0,
		parameter       pf2_pcie_cap_ep_l0s_accpt_latency                   = 0,
		parameter       pf2_pcie_cap_ep_l1_accpt_latency                    = 0,
		parameter       pf2_pcie_cap_l0s_exit_latency_commclk_dis           = 0,
		parameter       pf2_pcie_cap_l1_exit_latency_commclk_dis            = 0,
		parameter       pf3_pcie_cap_ep_l0s_accpt_latency                   = 0,
		parameter       pf3_pcie_cap_ep_l1_accpt_latency                    = 0,
		parameter       pf3_pcie_cap_l0s_exit_latency_commclk_dis           = 0,
		parameter       pf3_pcie_cap_l1_exit_latency_commclk_dis            = 0,
		parameter       pf0_pcie_cap_flr_cap                                = "PF0_PCIE_CAP_FLR_CAP_NOT_CAPABLE",
		parameter       pf1_pcie_cap_flr_cap                                = "PF1_PCIE_CAP_FLR_CAP_NOT_CAPABLE",
		parameter       pf2_pcie_cap_flr_cap                                = "PF2_PCIE_CAP_FLR_CAP_NOT_CAPABLE",
		parameter       pf3_pcie_cap_flr_cap                                = "PF3_PCIE_CAP_FLR_CAP_NOT_CAPABLE",
		parameter       pf0_pcie_cap_port_num                               = 1,
		parameter       pf1_pcie_cap_port_num                               = 0,
		parameter       pf2_pcie_cap_port_num                               = 0,
		parameter       pf3_pcie_cap_port_num                               = 0,
		parameter       pf0_pcie_cap_slot_clk_config                        = "true",
		parameter       pf1_pcie_cap_slot_clk_config                        = "false",
		parameter       pf2_pcie_cap_slot_clk_config                        = "false",
		parameter       pf3_pcie_cap_slot_clk_config                        = "false",
		parameter       pf0_ltr_cap_enable                                  = "PF0_LTR_CAP_ENABLE_DISABLED",
		parameter       pf0_pcie_slot_imp                                   = "PF0_PCIE_SLOT_IMP_NOT_IMPLEMENTED",
		parameter       pf0_pcie_cap_slot_power_limit_scale                 = 0,
		parameter       pf0_pcie_cap_slot_power_limit_value                 = 0,
		parameter       pf0_pcie_cap_phy_slot_num                           = 0,
		parameter       pf0_pcie_cap_hot_plug_capable                       = "false",
		parameter       pf0_pcie_cap_ext_tag_en                             = "true",
		parameter       pf1_pcie_cap_ext_tag_en                             = "false",
		parameter       pf2_pcie_cap_ext_tag_en                             = "false",
		parameter       pf3_pcie_cap_ext_tag_en                             = "false",
		parameter       cfg_ptm_auto_update_signal                          = "false",
		parameter       ptm_autoupdate                                      = "PTM_AUTOUPDATE_AUTOUPDATE_DISABLE",
		parameter       ptm_enable                                          = "PTM_ENABLE_DISABLE",
		parameter       pf0_ats_cap_enable                                  = "PF0_ATS_CAP_ENABLE_DISABLED",
		parameter       pf0_exvf_ats_cap_enable                             = "PF0_EXVF_ATS_CAP_ENABLE_DISABLED",
		parameter       pf0_ats_cap_invalidate_q_depth                      = 0,
		parameter       pf0_ats_exvf_align_request                          = "PF0_ATS_EXVF_ALIGN_REQUEST_DISABLE",
		parameter       pf1_ats_cap_enable                                  = "PF1_ATS_CAP_ENABLE_DISABLED",
		parameter       pf1_exvf_ats_cap_enable                             = "PF1_EXVF_ATS_CAP_ENABLE_DISABLED",
		parameter       pf1_ats_cap_invalidate_q_depth                      = 0,
		parameter       pf1_ats_exvf_align_request                          = "PF1_ATS_EXVF_ALIGN_REQUEST_DISABLE",
		parameter       pf2_ats_cap_enable                                  = "PF2_ATS_CAP_ENABLE_DISABLED",
		parameter       pf2_exvf_ats_cap_enable                             = "PF2_EXVF_ATS_CAP_ENABLE_DISABLED",
		parameter       pf2_ats_cap_invalidate_q_depth                      = 0,
		parameter       pf2_ats_exvf_align_request                          = "PF2_ATS_EXVF_ALIGN_REQUEST_DISABLE",
		parameter       pf3_ats_cap_enable                                  = "PF3_ATS_CAP_ENABLE_DISABLED",
		parameter       pf3_exvf_ats_cap_enable                             = "PF3_EXVF_ATS_CAP_ENABLE_DISABLED",
		parameter       pf3_ats_cap_invalidate_q_depth                      = 0,
		parameter       pf3_ats_exvf_align_request                          = "PF3_ATS_EXVF_ALIGN_REQUEST_DISABLE",
		parameter       pf0_tph_cap_enable                                  = "PF0_TPH_CAP_ENABLE_DISABLED",
		parameter       pf0_tph_req_cap_int_vec                             = "PF0_TPH_REQ_CAP_INT_VEC_DISABLED",
		parameter       pf0_tph_req_cap_int_vec_vfcomm_cs2                  = "PF0_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED",
		parameter       pf0_tph_req_cap_st_table_loc_0_vfcomm_cs2           = "PF0_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF",
		parameter       pf0_tph_req_cap_st_table_loc_1                      = "PF0_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE",
		parameter       pf0_tph_req_cap_st_table_loc_1_vfcomm_cs2           = "PF0_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF",
		parameter       pf0_tph_req_cap_st_table_size                       = 0,
		parameter       pf0_tph_req_cap_st_table_size_vfcomm_cs2            = 0,
		parameter       pf0_tph_req_device_spec                             = "PF0_TPH_REQ_DEVICE_SPEC_DISABLED",
		parameter       pf0_tph_req_device_spec_vfcomm_cs2                  = "PF0_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED",
		parameter       pf0_exvf_tph_cap_enable                             = "PF0_EXVF_TPH_CAP_ENABLE_DISABLED",
		parameter       exvf_tph_sttablelocation_pf0                        = 0,
		parameter       exvf_tph_sttablesize_pf0                            = 0,
		parameter       pf1_tph_cap_enable                                  = "PF1_TPH_CAP_ENABLE_DISABLED",
		parameter       pf1_tph_req_cap_int_vec                             = "PF1_TPH_REQ_CAP_INT_VEC_DISABLED",
		parameter       pf1_tph_req_cap_int_vec_vfcomm_cs2                  = "PF1_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED",
		parameter       pf1_tph_req_cap_st_table_loc_0_vfcomm_cs2           = "PF1_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF",
		parameter       pf1_tph_req_cap_st_table_loc_1                      = "PF1_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE",
		parameter       pf1_tph_req_cap_st_table_loc_1_vfcomm_cs2           = "PF1_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF",
		parameter       pf1_tph_req_cap_st_table_size                       = 0,
		parameter       pf1_tph_req_cap_st_table_size_vfcomm_cs2            = 0,
		parameter       pf1_tph_req_device_spec                             = "PF1_TPH_REQ_DEVICE_SPEC_DISABLED",
		parameter       pf1_tph_req_device_spec_vfcomm_cs2                  = "PF1_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED",
		parameter       pf1_exvf_tph_cap_enable                             = "PF1_EXVF_TPH_CAP_ENABLE_DISABLED",
		parameter       exvf_tph_sttablelocation_pf1                        = 0,
		parameter       exvf_tph_sttablesize_pf1                            = 0,
		parameter       pf2_tph_cap_enable                                  = "PF2_TPH_CAP_ENABLE_DISABLED",
		parameter       pf2_tph_req_cap_int_vec                             = "PF2_TPH_REQ_CAP_INT_VEC_DISABLED",
		parameter       pf2_tph_req_cap_int_vec_vfcomm_cs2                  = "PF2_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED",
		parameter       pf2_tph_req_cap_st_table_loc_0_vfcomm_cs2           = "PF2_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF",
		parameter       pf2_tph_req_cap_st_table_loc_1                      = "PF2_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE",
		parameter       pf2_tph_req_cap_st_table_loc_1_vfcomm_cs2           = "PF2_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF",
		parameter       pf2_tph_req_cap_st_table_size                       = 0,
		parameter       pf2_tph_req_cap_st_table_size_vfcomm_cs2            = 0,
		parameter       pf2_tph_req_device_spec                             = "PF2_TPH_REQ_DEVICE_SPEC_DISABLED",
		parameter       pf2_tph_req_device_spec_vfcomm_cs2                  = "PF2_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED",
		parameter       pf2_exvf_tph_cap_enable                             = "PF2_EXVF_TPH_CAP_ENABLE_DISABLED",
		parameter       exvf_tph_sttablelocation_pf2                        = 0,
		parameter       exvf_tph_sttablesize_pf2                            = 0,
		parameter       pf3_tph_cap_enable                                  = "PF3_TPH_CAP_ENABLE_DISABLED",
		parameter       pf3_tph_req_cap_int_vec                             = "PF3_TPH_REQ_CAP_INT_VEC_DISABLED",
		parameter       pf3_tph_req_cap_int_vec_vfcomm_cs2                  = "PF3_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED",
		parameter       pf3_tph_req_cap_st_table_loc_0_vfcomm_cs2           = "PF3_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF",
		parameter       pf3_tph_req_cap_st_table_loc_1                      = "PF3_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE",
		parameter       pf3_tph_req_cap_st_table_loc_1_vfcomm_cs2           = "PF3_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF",
		parameter       pf3_tph_req_cap_st_table_size                       = 0,
		parameter       pf3_tph_req_cap_st_table_size_vfcomm_cs2            = 0,
		parameter       pf3_tph_req_device_spec                             = "PF3_TPH_REQ_DEVICE_SPEC_DISABLED",
		parameter       pf3_tph_req_device_spec_vfcomm_cs2                  = "PF3_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED",
		parameter       pf3_exvf_tph_cap_enable                             = "PF3_EXVF_TPH_CAP_ENABLE_DISABLED",
		parameter       exvf_tph_sttablelocation_pf3                        = 0,
		parameter       exvf_tph_sttablesize_pf3                            = 0,
		parameter       pf0_acs_cap_enable                                  = "PF0_ACS_CAP_ENABLE_DISABLED",
		parameter       pf0_exvf_acs_cap_enable                             = "PF0_EXVF_ACS_CAP_ENABLE_DISABLED",
		parameter       pf0_acs_cap_acs_src_valid                           = "PF0_ACS_CAP_ACS_SRC_VALID_DISABLED",
		parameter       pf0_acs_cap_acs_at_block                            = "PF0_ACS_CAP_ACS_AT_BLOCK_DISABLED",
		parameter       pf0_acs_cap_acs_p2p_req_redirect                    = "PF0_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED",
		parameter       pf0_acs_cap_acs_p2p_cpl_redirect                    = "PF0_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED",
		parameter       pf0_acs_cap_acs_usp_forwarding                      = "PF0_ACS_CAP_ACS_USP_FORWARDING_DISABLED",
		parameter       pf0_acs_cap_acs_p2p_egress_control                  = "PF0_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED",
		parameter       pf0_acs_cap_acs_egress_ctrl_size                    = 8,
		parameter       pf0_acs_cap_acs_direct_translated_p2p               = "PF0_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED",
		parameter       pf1_acs_cap_enable                                  = "PF1_ACS_CAP_ENABLE_DISABLED",
		parameter       pf1_exvf_acs_cap_enable                             = "PF1_EXVF_ACS_CAP_ENABLE_DISABLED",
		parameter       pf1_acs_cap_acs_src_valid                           = "PF1_ACS_CAP_ACS_SRC_VALID_DISABLED",
		parameter       pf1_acs_cap_acs_at_block                            = "PF1_ACS_CAP_ACS_AT_BLOCK_DISABLED",
		parameter       pf1_acs_cap_acs_p2p_req_redirect                    = "PF1_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED",
		parameter       pf1_acs_cap_acs_p2p_cpl_redirect                    = "PF1_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED",
		parameter       pf1_acs_cap_acs_usp_forwarding                      = "PF1_ACS_CAP_ACS_USP_FORWARDING_DISABLED",
		parameter       pf1_acs_cap_acs_p2p_egress_control                  = "PF1_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED",
		parameter       pf1_acs_cap_acs_egress_ctrl_size                    = 8,
		parameter       pf1_acs_cap_acs_direct_translated_p2p               = "PF1_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED",
		parameter       pf2_acs_cap_enable                                  = "PF2_ACS_CAP_ENABLE_DISABLED",
		parameter       pf2_exvf_acs_cap_enable                             = "PF2_EXVF_ACS_CAP_ENABLE_DISABLED",
		parameter       pf2_acs_cap_acs_src_valid                           = "PF2_ACS_CAP_ACS_SRC_VALID_DISABLED",
		parameter       pf2_acs_cap_acs_at_block                            = "PF2_ACS_CAP_ACS_AT_BLOCK_DISABLED",
		parameter       pf2_acs_cap_acs_p2p_req_redirect                    = "PF2_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED",
		parameter       pf2_acs_cap_acs_p2p_cpl_redirect                    = "PF2_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED",
		parameter       pf2_acs_cap_acs_usp_forwarding                      = "PF2_ACS_CAP_ACS_USP_FORWARDING_DISABLED",
		parameter       pf2_acs_cap_acs_p2p_egress_control                  = "PF2_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED",
		parameter       pf2_acs_cap_acs_egress_ctrl_size                    = 8,
		parameter       pf2_acs_cap_acs_direct_translated_p2p               = "PF2_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED",
		parameter       pf3_acs_cap_enable                                  = "PF3_ACS_CAP_ENABLE_DISABLED",
		parameter       pf3_exvf_acs_cap_enable                             = "PF3_EXVF_ACS_CAP_ENABLE_DISABLED",
		parameter       pf3_acs_cap_acs_src_valid                           = "PF3_ACS_CAP_ACS_SRC_VALID_DISABLED",
		parameter       pf3_acs_cap_acs_at_block                            = "PF3_ACS_CAP_ACS_AT_BLOCK_DISABLED",
		parameter       pf3_acs_cap_acs_p2p_req_redirect                    = "PF3_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED",
		parameter       pf3_acs_cap_acs_p2p_cpl_redirect                    = "PF3_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED",
		parameter       pf3_acs_cap_acs_usp_forwarding                      = "PF3_ACS_CAP_ACS_USP_FORWARDING_DISABLED",
		parameter       pf3_acs_cap_acs_p2p_egress_control                  = "PF3_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED",
		parameter       pf3_acs_cap_acs_egress_ctrl_size                    = 8,
		parameter       pf3_acs_cap_acs_direct_translated_p2p               = "PF3_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED",
		parameter       pf0_virtio_en                                       = "PF0_VIRTIO_EN_DISABLED",
		parameter       pf1_virtio_en                                       = "PF1_VIRTIO_EN_DISABLED",
		parameter       pf2_virtio_en                                       = "PF2_VIRTIO_EN_DISABLED",
		parameter       pf3_virtio_en                                       = "PF3_VIRTIO_EN_DISABLED",
		parameter       pf0_exvf_virtio_en                                  = "PF0_EXVF_VIRTIO_EN_DISABLED",
		parameter       pf1_exvf_virtio_en                                  = "PF1_EXVF_VIRTIO_EN_DISABLED",
		parameter       pf2_exvf_virtio_en                                  = "PF2_EXVF_VIRTIO_EN_DISABLED",
		parameter       pf3_exvf_virtio_en                                  = "PF3_EXVF_VIRTIO_EN_DISABLED",
		parameter       pf0_pci_type0_device_id                             = 0,
		parameter       pf0_pci_type0_vendor_id                             = 4466,
		parameter       pf0_revision_id                                     = 1,
		parameter       pf0_base_class_code                                 = 255,
		parameter       pf0_subclass_code                                   = 0,
		parameter       pf0_program_interface                               = 0,
		parameter       pf0_subsys_vendor_id                                = 0,
		parameter       pf0_subsys_dev_id                                   = 0,
		parameter       pf0_sriov_vf_device_id                              = 0,
		parameter       exvf_subsysid_pf0                                   = 0,
		parameter       pf1_pci_type0_vendor_id                             = 0,
		parameter       pf1_pci_type0_device_id                             = 0,
		parameter       pf1_revision_id                                     = 0,
		parameter       pf1_base_class_code                                 = 0,
		parameter       pf1_subclass_code                                   = 0,
		parameter       pf1_program_interface                               = 0,
		parameter       pf1_subsys_vendor_id                                = 0,
		parameter       pf1_subsys_dev_id                                   = 0,
		parameter       pf1_sriov_vf_device_id                              = 0,
		parameter       exvf_subsysid_pf1                                   = 0,
		parameter       pf2_pci_type0_vendor_id                             = 0,
		parameter       pf2_pci_type0_device_id                             = 0,
		parameter       pf2_revision_id                                     = 0,
		parameter       pf2_base_class_code                                 = 0,
		parameter       pf2_subclass_code                                   = 0,
		parameter       pf2_program_interface                               = 0,
		parameter       pf2_subsys_vendor_id                                = 0,
		parameter       pf2_subsys_dev_id                                   = 0,
		parameter       pf2_sriov_vf_device_id                              = 0,
		parameter       exvf_subsysid_pf2                                   = 0,
		parameter       pf3_pci_type0_vendor_id                             = 0,
		parameter       pf3_pci_type0_device_id                             = 0,
		parameter       pf3_revision_id                                     = 0,
		parameter       pf3_base_class_code                                 = 0,
		parameter       pf3_subclass_code                                   = 0,
		parameter       pf3_program_interface                               = 0,
		parameter       pf3_subsys_vendor_id                                = 0,
		parameter       pf3_subsys_dev_id                                   = 0,
		parameter       pf3_sriov_vf_device_id                              = 0,
		parameter       exvf_subsysid_pf3                                   = 0,
		parameter       vsec_select                                         = "false",
		parameter       pf0_user_vsec_cap_enable                            = "PF0_USER_VSEC_CAP_ENABLE_DISABLED",
		parameter       pf1_user_vsec_cap_enable                            = "PF1_USER_VSEC_CAP_ENABLE_DISABLED",
		parameter       pf2_user_vsec_cap_enable                            = "PF2_USER_VSEC_CAP_ENABLE_DISABLED",
		parameter       pf3_user_vsec_cap_enable                            = "PF3_USER_VSEC_CAP_ENABLE_DISABLED",
		parameter       vsec_next_offset                                    = 0,
		parameter       pf1_user_vsec_offset                                = 0,
		parameter       pf2_user_vsec_offset                                = 0,
		parameter       pf3_user_vsec_offset                                = 0,
		parameter       cvp_vendor_specific_header_id                       = 0,
		parameter       drop_vendor0_msg                                    = "FALSE",
		parameter       drop_vendor1_msg                                    = "FALSE",
		parameter       pf0_int_pin                                         = "PF0_INT_PIN_NO_INT",
		parameter       pf1_int_pin                                         = "PF1_INT_PIN_NO_INT",
		parameter       pf2_int_pin                                         = "PF2_INT_PIN_NO_INT",
		parameter       pf3_int_pin                                         = "PF3_INT_PIN_NO_INT",
		parameter       dtk_mode_en                                         = "DTK_MODE_EN_ENABLE",
		parameter       hrc_arb_sel                                         = "HRC_ARB_SEL_LOCAL_QUAD_ARB",
		parameter       num_arb_ip                                          = 1,
		parameter       pcie_hrc_pulse_sel                                  = 0,
		parameter       pf0_port_logic_fast_link_mode                       = "PF0_PORT_LOGIC_FAST_LINK_MODE_DISABLE",
		parameter       pf0_prefetch_decode                                 = "PF0_PREFETCH_DECODE_PREF64",
		parameter       usb_hrc_pulse_sel                                   = 0,
		parameter       pcie_pcs_mode                                       = "PCIE_PCS_MODE_PCIE",
		parameter       sm_hssi_pcie_pcs_clk_mux_0_sel                      = "SEL_SAME_QUAD_PCLK0",
		parameter       sm_hssi_pcie_pcs_clk_mux_1_sel                      = "SEL_SAME_QUAD_PCLK0",
		parameter       sm_hssi_pcie_pcs_clk_mux_2_sel                      = "SEL_SAME_QUAD_PCLK0",
		parameter       sm_hssi_pcie_pcs_clk_mux_3_sel                      = "SEL_SAME_QUAD_PCLK0",
		parameter       sm_hssi_pcie_pcs_hps_clkmux_0_sel                   = "SEL_HPS_PCS1_ENABLED",
		parameter       sm_hssi_pcie_pcs_rst_mux_0_sel                      = "SEL_SAME_QUAD_PCS_RST",
		parameter       sm_hssi_pcie_pcs_rst_mux_1_sel                      = "SEL_SAME_QUAD_PCS_RST",
		parameter       sm_hssi_pcie_pcs_rst_mux_2_sel                      = "SEL_SAME_QUAD_PCS_RST",
		parameter       sm_hssi_pcie_pcs_rst_mux_3_sel                      = "SEL_SAME_QUAD_PCS_RST",
		parameter       sm_hssi_pcie_pcs_tx_mux_0_sel                       = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_tx_mux_1_sel                       = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_tx_mux_2_sel                       = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_tx_mux_3_sel                       = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_hps_demux_0_sel                    = "SEL_HPS_PCS1_ENABLED",
		parameter       sm_hssi_pcie_pcs_hps_mux_0_sel                      = "SEL_HPS_PCS1_ENABLED",
		parameter       sm_hssi_pcie_pcs_rx_demux_0_sel                     = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_rx_demux_1_sel                     = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_rx_demux_2_sel                     = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_pcs_rx_demux_3_sel                     = "SEL_SAME_QUAD_PCIE_CTRL",
		parameter       sm_hssi_pcie_clk_mux_0_sel                          = "SEL_MIDDLE",
		parameter       sm_hssi_pcie_data_mux_0_sel                         = "SEL_MIDDLE",
		parameter       sm_hssi_pld_chnl_dp_0_dr_enabled                    = "DR_ENABLED_DR_DISABLED",
		parameter       sm_hssi_pld_chnl_dp_0_duplex_mode                   = "DUPLEX_MODE_DUPLEX",
		parameter       sm_hssi_pld_chnl_dp_0_pld_channel_identifier        = "PLD_CHANNEL_IDENTIFIER_PHIP",
		parameter       sm_hssi_pld_chnl_dp_0_rx_clkout1_divider            = "RX_CLKOUT1_DIVIDER_DIV1",
		parameter       sm_hssi_pld_chnl_dp_0_rx_clkout2_divider            = "RX_CLKOUT2_DIVIDER_DIV1",
		parameter       sm_hssi_pld_chnl_dp_0_rx_en                         = "TRUE",
		parameter       sm_hssi_pld_chnl_dp_0_rx_fifo_mode                  = "RX_FIFO_MODE_PHASE_COMP",
		parameter       sm_hssi_pld_chnl_dp_0_rx_fifo_width                 = "RX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH",
		parameter[35:0] sm_hssi_pld_chnl_dp_0_rx_fifo_wr_clk_hz             = 36'b000000010001111000011010001100000000,
		parameter       sm_hssi_pld_chnl_dp_0_rx_user1_clk_dynamic_mux      = "RX_USER1_CLK_DYNAMIC_MUX_C2",
		parameter       sm_hssi_pld_chnl_dp_0_rx_user2_clk_dynamic_mux      = "RX_USER2_CLK_DYNAMIC_MUX_UX",
		parameter       sm_hssi_pld_chnl_dp_0_sup_mode                      = "SUP_MODE_USER_MODE",
		parameter       sm_hssi_pld_chnl_dp_0_tx_clkout1_divider            = "TX_CLKOUT1_DIVIDER_DIV1",
		parameter       sm_hssi_pld_chnl_dp_0_tx_clkout2_divider            = "TX_CLKOUT2_DIVIDER_DIV1",
		parameter       sm_hssi_pld_chnl_dp_0_tx_en                         = "TRUE",
		parameter       sm_hssi_pld_chnl_dp_0_tx_fifo_mode                  = "TX_FIFO_MODE_PHASE_COMP",
		parameter[35:0] sm_hssi_pld_chnl_dp_0_tx_fifo_rd_clk_hz             = 36'b000000010001111000011010001100000000,
		parameter       sm_hssi_pld_chnl_dp_0_tx_fifo_width                 = "TX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH",
		parameter       sm_hssi_pld_chnl_dp_0_tx_user1_clk_dynamic_mux      = "TX_USER1_CLK_DYNAMIC_MUX_C1",
		parameter       sm_hssi_pld_chnl_dp_0_tx_user2_clk_dynamic_mux      = "TX_USER2_CLK_DYNAMIC_MUX_UNUSED",
		parameter       sm_hssi_pld_chnl_dp_0_vc_rx_pldif_wm_en             = "VC_RX_PLDIF_WM_EN_DISABLE",
		parameter       sm_pld_rx_mux_0_sel                                 = "SEL_PCIE",
		parameter       sm_pld_tx_demux_0_sel                               = "SEL_PCIE",
		parameter       sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_sel           = "SEL_PCIE",
		parameter       sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_sel           = "SEL_PCIE"
	) (
		input  wire [((hal_num_of_lanes_hwtcl+1)*80)-1:0]  i_hio_txdata,                                //                           i_hio_txdata.data,                                        Stats Snapshot
		input  wire [((hal_num_of_lanes_hwtcl+1)*10)-1:0]  i_hio_txdata_extra,                          //                     i_hio_txdata_extra.data,                                        RX PFC
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_txdata_fifo_wr_en,                     //                i_hio_txdata_fifo_wr_en.data,                                        CSR access address
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rxdata_fifo_rd_en,                     //                i_hio_rxdata_fifo_rd_en.data,                                        RX error bits asserted on the EOP cycle
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_ptp_rst_n,                             //                        i_hio_ptp_rst_n.reset,                                       Stats Snapshot
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_ehip_rx_rst_n,                         //                    i_hio_ehip_rx_rst_n.reset,                                       RX PFC
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_ehip_tx_rst_n,                         //                    i_hio_ehip_tx_rst_n.reset,                                       CSR access address
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_ehip_signal_ok,                        //                   i_hio_ehip_signal_ok.reset,                                       RX error bits asserted on the EOP cycle
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_sfreeze_2_r03f_rx_mac_srfz_n,          //     i_hio_sfreeze_2_r03f_rx_mac_srfz_n.reset,                                       Stats Snapshot
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_sfreeze_3_c2f_tx_deskew_srfz_n,        //   i_hio_sfreeze_3_c2f_tx_deskew_srfz_n.reset,                                       RX PFC
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n,          //     i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n.reset,                                       CSR access address
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstfec_fec_rx_rst_n,                   //              i_hio_rstfec_fec_rx_rst_n.reset,                                       RX error bits asserted on the EOP cycle
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstfec_fec_tx_rst_n,                   //              i_hio_rstfec_fec_tx_rst_n.reset,                                       RX error bits asserted on the EOP cycle
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstfec_fec_csr_ret,                    //               i_hio_rstfec_fec_csr_ret.reset,                                       Stats Snapshot
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstfec_rx_fec_sfrz_n,                  //             i_hio_rstfec_rx_fec_sfrz_n.reset,                                       RX PFC
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstfec_tx_fec_sfrz_n,                  //             i_hio_rstfec_tx_fec_sfrz_n.reset,                                       CSR access address
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstxcvrif_xcvrif_rx_rst_n,             //        i_hio_rstxcvrif_xcvrif_rx_rst_n.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstxcvrif_xcvrif_tx_rst_n,             //        i_hio_rstxcvrif_xcvrif_tx_rst_n.reset,                                       Stats Snapshot
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstxcvrif_xcvrif_signal_ok,            //       i_hio_rstxcvrif_xcvrif_signal_ok.reset,                                       RX PFC
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstxcvrif_rx_xcvrif_sfrz_n,            //       i_hio_rstxcvrif_rx_xcvrif_sfrz_n.reset,                                       CSR access address
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rstxcvrif_tx_xcvrif_sfrz_n,            //       i_hio_rstxcvrif_tx_xcvrif_sfrz_n.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_pld_clrhip,                        //                   i_hio_rst_pld_clrhip.reset,                                       Stats Snapshot
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_pld_clrpcs,                        //                   i_hio_rst_pld_clrpcs.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_pld_perstn,                        //                   i_hio_rst_pld_perstn.reset,                                       CSR access address
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_pld_ready,                         //                    i_hio_rst_pld_ready.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_pld_adapter_rx_pld_rst_n,          //     i_hio_rst_pld_adapter_rx_pld_rst_n.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_pld_adapter_tx_pld_rst_n,          //     i_hio_rst_pld_adapter_tx_pld_rst_n.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_ux_rx_pma_rst_n,                   //              i_hio_rst_ux_rx_pma_rst_n.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_ux_rx_sfrz,                        //                   i_hio_rst_ux_rx_sfrz.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_rst_ux_tx_pma_rst_n,                   //              i_hio_rst_ux_tx_pma_rst_n.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   i_hio_pld_reset_clk_row,                     //                i_hio_pld_reset_clk_row.reset
		input  wire [((hal_num_of_lanes_hwtcl+1)*80)-1:0]  i_hio_uxquad_async,                          //                     i_hio_uxquad_async.data
		input  wire [((hal_num_of_lanes_hwtcl+1)*80)-1:0]  i_hio_uxquad_async_pcie_mux,                 //            i_hio_uxquad_async_pcie_mux.data
		input  wire [(hal_num_of_lanes_hwtcl*1)-1:0]       rx_serial_n,                                 //                            rx_serial_n.data
		input  wire [(hal_num_of_lanes_hwtcl*1)-1:0]       rx_serial_p,                                 //                            rx_serial_p.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_txdata_fifo_wr_empty,                  //             o_hio_txdata_fifo_wr_empty.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_txdata_fifo_wr_pempty,                 //            o_hio_txdata_fifo_wr_pempty.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_txdata_fifo_wr_full,                   //              o_hio_txdata_fifo_wr_full.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_txdata_fifo_wr_pfull,                  //             o_hio_txdata_fifo_wr_pfull.data
		output wire [((hal_num_of_lanes_hwtcl+1)*80)-1:0]  o_hio_rxdata,                                //                           o_hio_rxdata.data
		output wire [((hal_num_of_lanes_hwtcl+1)*10)-1:0]  o_hio_rxdata_extra,                          //                     o_hio_rxdata_extra.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rxdata_fifo_rd_empty,                  //             o_hio_rxdata_fifo_rd_empty.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rxdata_fifo_rd_pempty,                 //            o_hio_rxdata_fifo_rd_pempty.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rxdata_fifo_rd_full,                   //              o_hio_rxdata_fifo_rd_full.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rxdata_fifo_rd_pfull,                  //             o_hio_rxdata_fifo_rd_pfull.data
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rstepcs_rx_pcs_fully_aligned,          //     o_hio_rstepcs_rx_pcs_fully_aligned.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rstfec_fec_rx_rdy_n,                   //              o_hio_rstfec_fec_rx_rdy_n.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_flux0_cpi_cmn_busy,                //           o_hio_rst_flux0_cpi_cmn_busy.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_oflux_rx_srds_rdy,                 //            o_hio_rst_oflux_rx_srds_rdy.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_ux_all_synthlockstatus,            //       o_hio_rst_ux_all_synthlockstatus.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_ux_octl_pcs_rxstatus,              //         o_hio_rst_ux_octl_pcs_rxstatus.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_ux_octl_pcs_txstatus,              //         o_hio_rst_ux_octl_pcs_txstatus.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_ux_rxcdrlock2data,                 //            o_hio_rst_ux_rxcdrlock2data.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*1)-1:0]   o_hio_rst_ux_rxcdrlockstatus,                //           o_hio_rst_ux_rxcdrlockstatus.reset
		output wire [((hal_num_of_lanes_hwtcl+1)*50)-1:0]  o_hio_uxquad_async,                          //                     o_hio_uxquad_async.data
		output wire [(hal_num_of_lanes_hwtcl*1)-1:0]       tx_serial_p,                                 //                            tx_serial_p.data
		output wire [(hal_num_of_lanes_hwtcl*1)-1:0]       tx_serial_n,                                 //                            tx_serial_n.data
		input  wire [((hal_num_of_lanes_hwtcl+1)*100)-1:0] i_hio_txdata_async,                          //                     i_hio_txdata_async.data
		input  wire [((hal_num_of_lanes_hwtcl+1)*10)-1:0]  i_hio_txdata_direct,                         //                    i_hio_txdata_direct.data
		output wire [((hal_num_of_lanes_hwtcl+1)*100)-1:0] o_hio_rxdata_async,                          //                     o_hio_rxdata_async.data
		output wire [((hal_num_of_lanes_hwtcl+1)*10)-1:0]  o_hio_rxdata_direct,                         //                    o_hio_rxdata_direct.data
		output wire [(hal_num_of_lanes_hwtcl*1)-1:0]       ioack_cdrdiv_left_ux_bidir_out,              //         ioack_cdrdiv_left_ux_bidir_out.data
		input  wire                                        i_refclk_tx_p,                               //                          i_refclk_tx_p.clk
		input  wire                                        i_syspll_c0_clk,                             //                        i_syspll_c0_clk.clk
		input  wire                                        i_syspll_c1_clk,                             //                        i_syspll_c1_clk.clk
		input  wire                                        i_syspll_c2_clk,                             //                        i_syspll_c2_clk.clk
		input  wire                                        i_flux_clk,                                  //                             i_flux_clk.clk
		input  wire                                        i_flux_clk_1,                                //                           i_flux_clk_1.clk
		input  wire                                        i_refclk_rx_p,                               //                          i_refclk_rx_p.clk
		input  wire                                        i_ss_vccl_syspll_locked,                     //                i_ss_vccl_syspll_locked.clk
		output wire                                        o_hio_pcie_user_rx_clk1_clk,                 //            o_hio_pcie_user_rx_clk1_clk.clk
		output wire                                        o_hio_pcie_user_rx_clk2_clk,                 //            o_hio_pcie_user_rx_clk2_clk.clk
		output wire                                        o_hio_pcie_user_tx_clk1_clk,                 //            o_hio_pcie_user_tx_clk1_clk.clk
		output wire                                        o_hio_pcie_user_tx_clk2_clk,                 //            o_hio_pcie_user_tx_clk2_clk.clk
		output wire                                        o_pcs4_pipe_rst_n,                           //                               phip_hal.o_pcs4_pipe_rst_n,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe4_dirfeedback,                       //                                       .i_rxpipe4_dirfeedback,                       Check User Guide for details
		input  wire [7:0]                                  i_rxpipe4_linkevaluationfeedbackfiguremerit, //                                       .i_rxpipe4_linkevaluationfeedbackfiguremerit, Check User Guide for details
		input  wire [5:0]                                  i_rxpipe4_localfs,                           //                                       .i_rxpipe4_localfs,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe4_locallf,                           //                                       .i_rxpipe4_locallf,                           Check User Guide for details
		input  wire                                        i_rxpipe4_localtxcoefficientsvalid,          //                                       .i_rxpipe4_localtxcoefficientsvalid,          Check User Guide for details
		input  wire [17:0]                                 i_rxpipe4_localtxpresetcoefficients,         //                                       .i_rxpipe4_localtxpresetcoefficients,         Check User Guide for details
		input  wire [7:0]                                  i_rxpipe4_p2m_bus,                           //                                       .i_rxpipe4_p2m_bus,                           Check User Guide for details
		input  wire                                        i_rxpipe4_pclkchangeok,                      //                                       .i_rxpipe4_pclkchangeok,                      Check User Guide for details
		input  wire                                        i_rxpipe4_phystatus,                         //                                       .i_rxpipe4_phystatus,                         Check User Guide for details
		input  wire [39:0]                                 i_rxpipe4_rxdata,                            //                                       .i_rxpipe4_rxdata,                            Check User Guide for details
		input  wire [3:0]                                  i_rxpipe4_rxdatak,                           //                                       .i_rxpipe4_rxdatak,                           Check User Guide for details
		input  wire                                        i_rxpipe4_rxdatavalid,                       //                                       .i_rxpipe4_rxdatavalid,                       Check User Guide for details
		input  wire                                        i_rxpipe4_rxelecidlea,                       //                                       .i_rxpipe4_rxelecidlea,                       Check User Guide for details
		input  wire                                        i_rxpipe4_rxstandbystatus,                   //                                       .i_rxpipe4_rxstandbystatus,                   Check User Guide for details
		input  wire                                        i_rxpipe4_rxstartblock,                      //                                       .i_rxpipe4_rxstartblock,                      Check User Guide for details
		input  wire [2:0]                                  i_rxpipe4_rxstatus,                          //                                       .i_rxpipe4_rxstatus,                          Check User Guide for details
		input  wire [3:0]                                  i_rxpipe4_rxsyncheader,                      //                                       .i_rxpipe4_rxsyncheader,                      Check User Guide for details
		input  wire                                        i_rxpipe4_rxvalid,                           //                                       .i_rxpipe4_rxvalid,                           Check User Guide for details
		output wire                                        o_txpipe4_asyncpowerchangeack,               //                                       .o_txpipe4_asyncpowerchangeack,               Check User Guide for details
		output wire                                        o_txpipe4_blockaligncontrol,                 //                                       .o_txpipe4_blockaligncontrol,                 Check User Guide for details
		output wire                                        o_txpipe4_cfg_hw_auto_sp_dis,                //                                       .o_txpipe4_cfg_hw_auto_sp_dis,                Check User Guide for details
		output wire                                        o_txpipe4_dirchange,                         //                                       .o_txpipe4_dirchange,                         Check User Guide for details
		output wire                                        o_txpipe4_ebuf_mode,                         //                                       .o_txpipe4_ebuf_mode,                         Check User Guide for details
		output wire                                        o_txpipe4_encodedecodebypass,                //                                       .o_txpipe4_encodedecodebypass,                Check User Guide for details
		output wire [5:0]                                  o_txpipe4_fs,                                //                                       .o_txpipe4_fs,                                Check User Guide for details
		output wire                                        o_txpipe4_getlocalpresetcoefficients,        //                                       .o_txpipe4_getlocalpresetcoefficients,        Check User Guide for details
		output wire                                        o_txpipe4_invalidrequest,                    //                                       .o_txpipe4_invalidrequest,                    Check User Guide for details
		output wire [5:0]                                  o_txpipe4_lf,                                //                                       .o_txpipe4_lf,                                Check User Guide for details
		output wire [4:0]                                  o_txpipe4_localpresetindex,                  //                                       .o_txpipe4_localpresetindex,                  Check User Guide for details
		output wire                                        o_txpipe4_lowpin_nt,                         //                                       .o_txpipe4_lowpin_nt,                         Check User Guide for details
		output wire [7:0]                                  o_txpipe4_m2p_bus,                           //                                       .o_txpipe4_m2p_bus,                           Check User Guide for details
		output wire [2:0]                                  o_txpipe4_pclk_rate,                         //                                       .o_txpipe4_pclk_rate,                         Check User Guide for details
		output wire                                        o_txpipe4_pclkchangeack,                     //                                       .o_txpipe4_pclkchangeack,                     Check User Guide for details
		output wire [3:0]                                  o_txpipe4_phy_mode_nt,                       //                                       .o_txpipe4_phy_mode_nt,                       Check User Guide for details
		output wire [3:0]                                  o_txpipe4_powerdown,                         //                                       .o_txpipe4_powerdown,                         Check User Guide for details
		output wire [2:0]                                  o_txpipe4_rate,                              //                                       .o_txpipe4_rate,                              Check User Guide for details
		output wire                                        o_txpipe4_rxelecidle_disable_a,              //                                       .o_txpipe4_rxelecidle_disable_a,              Check User Guide for details
		output wire                                        o_txpipe4_rxeqclr,                           //                                       .o_txpipe4_rxeqclr,                           Check User Guide for details
		output wire                                        o_txpipe4_rxeqeval,                          //                                       .o_txpipe4_rxeqeval,                          Check User Guide for details
		output wire                                        o_txpipe4_rxeqinprogress,                    //                                       .o_txpipe4_rxeqinprogress,                    Check User Guide for details
		output wire                                        o_txpipe4_rxeqtraining,                      //                                       .o_txpipe4_rxeqtraining,                      Check User Guide for details
		output wire                                        o_txpipe4_rxpolarity,                        //                                       .o_txpipe4_rxpolarity,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe4_rxpresethint,                      //                                       .o_txpipe4_rxpresethint,                      Check User Guide for details
		output wire                                        o_txpipe4_rxstandby,                         //                                       .o_txpipe4_rxstandby,                         Check User Guide for details
		output wire                                        o_txpipe4_rxtermination,                     //                                       .o_txpipe4_rxtermination,                     Check User Guide for details
		output wire                                        o_txpipe4_srisenable,                        //                                       .o_txpipe4_srisenable,                        Check User Guide for details
		output wire                                        o_txpipe4_txcmnmode_disable_a,               //                                       .o_txpipe4_txcmnmode_disable_a,               Check User Guide for details
		output wire                                        o_txpipe4_txcompliance,                      //                                       .o_txpipe4_txcompliance,                      Check User Guide for details
		output wire [39:0]                                 o_txpipe4_txdata,                            //                                       .o_txpipe4_txdata,                            Check User Guide for details
		output wire [3:0]                                  o_txpipe4_txdatak,                           //                                       .o_txpipe4_txdatak,                           Check User Guide for details
		output wire                                        o_txpipe4_txdatavalid,                       //                                       .o_txpipe4_txdatavalid,                       Check User Guide for details
		output wire [17:0]                                 o_txpipe4_txdeemph,                          //                                       .o_txpipe4_txdeemph,                          Check User Guide for details
		output wire                                        o_txpipe4_txdtctrx_lb,                       //                                       .o_txpipe4_txdtctrx_lb,                       Check User Guide for details
		output wire                                        o_txpipe4_txelecidle,                        //                                       .o_txpipe4_txelecidle,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe4_txmargin,                          //                                       .o_txpipe4_txmargin,                          Check User Guide for details
		output wire                                        o_txpipe4_txoneszeros,                       //                                       .o_txpipe4_txoneszeros,                       Check User Guide for details
		output wire                                        o_txpipe4_txstartblock,                      //                                       .o_txpipe4_txstartblock,                      Check User Guide for details
		output wire                                        o_txpipe4_txswing,                           //                                       .o_txpipe4_txswing,                           Check User Guide for details
		output wire [3:0]                                  o_txpipe4_txsyncheader,                      //                                       .o_txpipe4_txsyncheader,                      Check User Guide for details
		output wire [2:0]                                  o_txpipe4_width,                             //                                       .o_txpipe4_width,                             Check User Guide for details
		output wire                                        o_pcs5_pipe_rst_n,                           //                                       .o_pcs5_pipe_rst_n,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe5_dirfeedback,                       //                                       .i_rxpipe5_dirfeedback,                       Check User Guide for details
		input  wire [7:0]                                  i_rxpipe5_linkevaluationfeedbackfiguremerit, //                                       .i_rxpipe5_linkevaluationfeedbackfiguremerit, Check User Guide for details
		input  wire [5:0]                                  i_rxpipe5_localfs,                           //                                       .i_rxpipe5_localfs,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe5_locallf,                           //                                       .i_rxpipe5_locallf,                           Check User Guide for details
		input  wire                                        i_rxpipe5_localtxcoefficientsvalid,          //                                       .i_rxpipe5_localtxcoefficientsvalid,          Check User Guide for details
		input  wire [17:0]                                 i_rxpipe5_localtxpresetcoefficients,         //                                       .i_rxpipe5_localtxpresetcoefficients,         Check User Guide for details
		input  wire [7:0]                                  i_rxpipe5_p2m_bus,                           //                                       .i_rxpipe5_p2m_bus,                           Check User Guide for details
		input  wire                                        i_rxpipe5_pclkchangeok,                      //                                       .i_rxpipe5_pclkchangeok,                      Check User Guide for details
		input  wire                                        i_rxpipe5_phystatus,                         //                                       .i_rxpipe5_phystatus,                         Check User Guide for details
		input  wire [39:0]                                 i_rxpipe5_rxdata,                            //                                       .i_rxpipe5_rxdata,                            Check User Guide for details
		input  wire [3:0]                                  i_rxpipe5_rxdatak,                           //                                       .i_rxpipe5_rxdatak,                           Check User Guide for details
		input  wire                                        i_rxpipe5_rxdatavalid,                       //                                       .i_rxpipe5_rxdatavalid,                       Check User Guide for details
		input  wire                                        i_rxpipe5_rxelecidlea,                       //                                       .i_rxpipe5_rxelecidlea,                       Check User Guide for details
		input  wire                                        i_rxpipe5_rxstandbystatus,                   //                                       .i_rxpipe5_rxstandbystatus,                   Check User Guide for details
		input  wire                                        i_rxpipe5_rxstartblock,                      //                                       .i_rxpipe5_rxstartblock,                      Check User Guide for details
		input  wire [2:0]                                  i_rxpipe5_rxstatus,                          //                                       .i_rxpipe5_rxstatus,                          Check User Guide for details
		input  wire [3:0]                                  i_rxpipe5_rxsyncheader,                      //                                       .i_rxpipe5_rxsyncheader,                      Check User Guide for details
		input  wire                                        i_rxpipe5_rxvalid,                           //                                       .i_rxpipe5_rxvalid,                           Check User Guide for details
		output wire                                        o_txpipe5_asyncpowerchangeack,               //                                       .o_txpipe5_asyncpowerchangeack,               Check User Guide for details
		output wire                                        o_txpipe5_blockaligncontrol,                 //                                       .o_txpipe5_blockaligncontrol,                 Check User Guide for details
		output wire                                        o_txpipe5_cfg_hw_auto_sp_dis,                //                                       .o_txpipe5_cfg_hw_auto_sp_dis,                Check User Guide for details
		output wire                                        o_txpipe5_dirchange,                         //                                       .o_txpipe5_dirchange,                         Check User Guide for details
		output wire                                        o_txpipe5_ebuf_mode,                         //                                       .o_txpipe5_ebuf_mode,                         Check User Guide for details
		output wire                                        o_txpipe5_encodedecodebypass,                //                                       .o_txpipe5_encodedecodebypass,                Check User Guide for details
		output wire [5:0]                                  o_txpipe5_fs,                                //                                       .o_txpipe5_fs,                                Check User Guide for details
		output wire                                        o_txpipe5_getlocalpresetcoefficients,        //                                       .o_txpipe5_getlocalpresetcoefficients,        Check User Guide for details
		output wire                                        o_txpipe5_invalidrequest,                    //                                       .o_txpipe5_invalidrequest,                    Check User Guide for details
		output wire [5:0]                                  o_txpipe5_lf,                                //                                       .o_txpipe5_lf,                                Check User Guide for details
		output wire [4:0]                                  o_txpipe5_localpresetindex,                  //                                       .o_txpipe5_localpresetindex,                  Check User Guide for details
		output wire                                        o_txpipe5_lowpin_nt,                         //                                       .o_txpipe5_lowpin_nt,                         Check User Guide for details
		output wire [7:0]                                  o_txpipe5_m2p_bus,                           //                                       .o_txpipe5_m2p_bus,                           Check User Guide for details
		output wire [2:0]                                  o_txpipe5_pclk_rate,                         //                                       .o_txpipe5_pclk_rate,                         Check User Guide for details
		output wire                                        o_txpipe5_pclkchangeack,                     //                                       .o_txpipe5_pclkchangeack,                     Check User Guide for details
		output wire [3:0]                                  o_txpipe5_phy_mode_nt,                       //                                       .o_txpipe5_phy_mode_nt,                       Check User Guide for details
		output wire [3:0]                                  o_txpipe5_powerdown,                         //                                       .o_txpipe5_powerdown,                         Check User Guide for details
		output wire [2:0]                                  o_txpipe5_rate,                              //                                       .o_txpipe5_rate,                              Check User Guide for details
		output wire                                        o_txpipe5_rxelecidle_disable_a,              //                                       .o_txpipe5_rxelecidle_disable_a,              Check User Guide for details
		output wire                                        o_txpipe5_rxeqclr,                           //                                       .o_txpipe5_rxeqclr,                           Check User Guide for details
		output wire                                        o_txpipe5_rxeqeval,                          //                                       .o_txpipe5_rxeqeval,                          Check User Guide for details
		output wire                                        o_txpipe5_rxeqinprogress,                    //                                       .o_txpipe5_rxeqinprogress,                    Check User Guide for details
		output wire                                        o_txpipe5_rxeqtraining,                      //                                       .o_txpipe5_rxeqtraining,                      Check User Guide for details
		output wire                                        o_txpipe5_rxpolarity,                        //                                       .o_txpipe5_rxpolarity,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe5_rxpresethint,                      //                                       .o_txpipe5_rxpresethint,                      Check User Guide for details
		output wire                                        o_txpipe5_rxstandby,                         //                                       .o_txpipe5_rxstandby,                         Check User Guide for details
		output wire                                        o_txpipe5_rxtermination,                     //                                       .o_txpipe5_rxtermination,                     Check User Guide for details
		output wire                                        o_txpipe5_srisenable,                        //                                       .o_txpipe5_srisenable,                        Check User Guide for details
		output wire                                        o_txpipe5_txcmnmode_disable_a,               //                                       .o_txpipe5_txcmnmode_disable_a,               Check User Guide for details
		output wire                                        o_txpipe5_txcompliance,                      //                                       .o_txpipe5_txcompliance,                      Check User Guide for details
		output wire [39:0]                                 o_txpipe5_txdata,                            //                                       .o_txpipe5_txdata,                            Check User Guide for details
		output wire [3:0]                                  o_txpipe5_txdatak,                           //                                       .o_txpipe5_txdatak,                           Check User Guide for details
		output wire                                        o_txpipe5_txdatavalid,                       //                                       .o_txpipe5_txdatavalid,                       Check User Guide for details
		output wire [17:0]                                 o_txpipe5_txdeemph,                          //                                       .o_txpipe5_txdeemph,                          Check User Guide for details
		output wire                                        o_txpipe5_txdtctrx_lb,                       //                                       .o_txpipe5_txdtctrx_lb,                       Check User Guide for details
		output wire                                        o_txpipe5_txelecidle,                        //                                       .o_txpipe5_txelecidle,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe5_txmargin,                          //                                       .o_txpipe5_txmargin,                          Check User Guide for details
		output wire                                        o_txpipe5_txoneszeros,                       //                                       .o_txpipe5_txoneszeros,                       Check User Guide for details
		output wire                                        o_txpipe5_txstartblock,                      //                                       .o_txpipe5_txstartblock,                      Check User Guide for details
		output wire                                        o_txpipe5_txswing,                           //                                       .o_txpipe5_txswing,                           Check User Guide for details
		output wire [3:0]                                  o_txpipe5_txsyncheader,                      //                                       .o_txpipe5_txsyncheader,                      Check User Guide for details
		output wire [2:0]                                  o_txpipe5_width,                             //                                       .o_txpipe5_width,                             Check User Guide for details
		output wire                                        o_pcs6_pipe_rst_n,                           //                                       .o_pcs6_pipe_rst_n,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe6_dirfeedback,                       //                                       .i_rxpipe6_dirfeedback,                       Check User Guide for details
		input  wire [7:0]                                  i_rxpipe6_linkevaluationfeedbackfiguremerit, //                                       .i_rxpipe6_linkevaluationfeedbackfiguremerit, Check User Guide for details
		input  wire [5:0]                                  i_rxpipe6_localfs,                           //                                       .i_rxpipe6_localfs,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe6_locallf,                           //                                       .i_rxpipe6_locallf,                           Check User Guide for details
		input  wire                                        i_rxpipe6_localtxcoefficientsvalid,          //                                       .i_rxpipe6_localtxcoefficientsvalid,          Check User Guide for details
		input  wire [17:0]                                 i_rxpipe6_localtxpresetcoefficients,         //                                       .i_rxpipe6_localtxpresetcoefficients,         Check User Guide for details
		input  wire [7:0]                                  i_rxpipe6_p2m_bus,                           //                                       .i_rxpipe6_p2m_bus,                           Check User Guide for details
		input  wire                                        i_rxpipe6_pclkchangeok,                      //                                       .i_rxpipe6_pclkchangeok,                      Check User Guide for details
		input  wire                                        i_rxpipe6_phystatus,                         //                                       .i_rxpipe6_phystatus,                         Check User Guide for details
		input  wire [39:0]                                 i_rxpipe6_rxdata,                            //                                       .i_rxpipe6_rxdata,                            Check User Guide for details
		input  wire [3:0]                                  i_rxpipe6_rxdatak,                           //                                       .i_rxpipe6_rxdatak,                           Check User Guide for details
		input  wire                                        i_rxpipe6_rxdatavalid,                       //                                       .i_rxpipe6_rxdatavalid,                       Check User Guide for details
		input  wire                                        i_rxpipe6_rxelecidlea,                       //                                       .i_rxpipe6_rxelecidlea,                       Check User Guide for details
		input  wire                                        i_rxpipe6_rxstandbystatus,                   //                                       .i_rxpipe6_rxstandbystatus,                   Check User Guide for details
		input  wire                                        i_rxpipe6_rxstartblock,                      //                                       .i_rxpipe6_rxstartblock,                      Check User Guide for details
		input  wire [2:0]                                  i_rxpipe6_rxstatus,                          //                                       .i_rxpipe6_rxstatus,                          Check User Guide for details
		input  wire [3:0]                                  i_rxpipe6_rxsyncheader,                      //                                       .i_rxpipe6_rxsyncheader,                      Check User Guide for details
		input  wire                                        i_rxpipe6_rxvalid,                           //                                       .i_rxpipe6_rxvalid,                           Check User Guide for details
		output wire                                        o_txpipe6_asyncpowerchangeack,               //                                       .o_txpipe6_asyncpowerchangeack,               Check User Guide for details
		output wire                                        o_txpipe6_blockaligncontrol,                 //                                       .o_txpipe6_blockaligncontrol,                 Check User Guide for details
		output wire                                        o_txpipe6_cfg_hw_auto_sp_dis,                //                                       .o_txpipe6_cfg_hw_auto_sp_dis,                Check User Guide for details
		output wire                                        o_txpipe6_dirchange,                         //                                       .o_txpipe6_dirchange,                         Check User Guide for details
		output wire                                        o_txpipe6_ebuf_mode,                         //                                       .o_txpipe6_ebuf_mode,                         Check User Guide for details
		output wire                                        o_txpipe6_encodedecodebypass,                //                                       .o_txpipe6_encodedecodebypass,                Check User Guide for details
		output wire [5:0]                                  o_txpipe6_fs,                                //                                       .o_txpipe6_fs,                                Check User Guide for details
		output wire                                        o_txpipe6_getlocalpresetcoefficients,        //                                       .o_txpipe6_getlocalpresetcoefficients,        Check User Guide for details
		output wire                                        o_txpipe6_invalidrequest,                    //                                       .o_txpipe6_invalidrequest,                    Check User Guide for details
		output wire [5:0]                                  o_txpipe6_lf,                                //                                       .o_txpipe6_lf,                                Check User Guide for details
		output wire [4:0]                                  o_txpipe6_localpresetindex,                  //                                       .o_txpipe6_localpresetindex,                  Check User Guide for details
		output wire                                        o_txpipe6_lowpin_nt,                         //                                       .o_txpipe6_lowpin_nt,                         Check User Guide for details
		output wire [7:0]                                  o_txpipe6_m2p_bus,                           //                                       .o_txpipe6_m2p_bus,                           Check User Guide for details
		output wire [2:0]                                  o_txpipe6_pclk_rate,                         //                                       .o_txpipe6_pclk_rate,                         Check User Guide for details
		output wire                                        o_txpipe6_pclkchangeack,                     //                                       .o_txpipe6_pclkchangeack,                     Check User Guide for details
		output wire [3:0]                                  o_txpipe6_phy_mode_nt,                       //                                       .o_txpipe6_phy_mode_nt,                       Check User Guide for details
		output wire [3:0]                                  o_txpipe6_powerdown,                         //                                       .o_txpipe6_powerdown,                         Check User Guide for details
		output wire [2:0]                                  o_txpipe6_rate,                              //                                       .o_txpipe6_rate,                              Check User Guide for details
		output wire                                        o_txpipe6_rxelecidle_disable_a,              //                                       .o_txpipe6_rxelecidle_disable_a,              Check User Guide for details
		output wire                                        o_txpipe6_rxeqclr,                           //                                       .o_txpipe6_rxeqclr,                           Check User Guide for details
		output wire                                        o_txpipe6_rxeqeval,                          //                                       .o_txpipe6_rxeqeval,                          Check User Guide for details
		output wire                                        o_txpipe6_rxeqinprogress,                    //                                       .o_txpipe6_rxeqinprogress,                    Check User Guide for details
		output wire                                        o_txpipe6_rxeqtraining,                      //                                       .o_txpipe6_rxeqtraining,                      Check User Guide for details
		output wire                                        o_txpipe6_rxpolarity,                        //                                       .o_txpipe6_rxpolarity,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe6_rxpresethint,                      //                                       .o_txpipe6_rxpresethint,                      Check User Guide for details
		output wire                                        o_txpipe6_rxstandby,                         //                                       .o_txpipe6_rxstandby,                         Check User Guide for details
		output wire                                        o_txpipe6_rxtermination,                     //                                       .o_txpipe6_rxtermination,                     Check User Guide for details
		output wire                                        o_txpipe6_srisenable,                        //                                       .o_txpipe6_srisenable,                        Check User Guide for details
		output wire                                        o_txpipe6_txcmnmode_disable_a,               //                                       .o_txpipe6_txcmnmode_disable_a,               Check User Guide for details
		output wire                                        o_txpipe6_txcompliance,                      //                                       .o_txpipe6_txcompliance,                      Check User Guide for details
		output wire [39:0]                                 o_txpipe6_txdata,                            //                                       .o_txpipe6_txdata,                            Check User Guide for details
		output wire [3:0]                                  o_txpipe6_txdatak,                           //                                       .o_txpipe6_txdatak,                           Check User Guide for details
		output wire                                        o_txpipe6_txdatavalid,                       //                                       .o_txpipe6_txdatavalid,                       Check User Guide for details
		output wire [17:0]                                 o_txpipe6_txdeemph,                          //                                       .o_txpipe6_txdeemph,                          Check User Guide for details
		output wire                                        o_txpipe6_txdtctrx_lb,                       //                                       .o_txpipe6_txdtctrx_lb,                       Check User Guide for details
		output wire                                        o_txpipe6_txelecidle,                        //                                       .o_txpipe6_txelecidle,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe6_txmargin,                          //                                       .o_txpipe6_txmargin,                          Check User Guide for details
		output wire                                        o_txpipe6_txoneszeros,                       //                                       .o_txpipe6_txoneszeros,                       Check User Guide for details
		output wire                                        o_txpipe6_txstartblock,                      //                                       .o_txpipe6_txstartblock,                      Check User Guide for details
		output wire                                        o_txpipe6_txswing,                           //                                       .o_txpipe6_txswing,                           Check User Guide for details
		output wire [3:0]                                  o_txpipe6_txsyncheader,                      //                                       .o_txpipe6_txsyncheader,                      Check User Guide for details
		output wire [2:0]                                  o_txpipe6_width,                             //                                       .o_txpipe6_width,                             Check User Guide for details
		output wire                                        o_pcs7_pipe_rst_n,                           //                                       .o_pcs7_pipe_rst_n,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe7_dirfeedback,                       //                                       .i_rxpipe7_dirfeedback,                       Check User Guide for details
		input  wire [7:0]                                  i_rxpipe7_linkevaluationfeedbackfiguremerit, //                                       .i_rxpipe7_linkevaluationfeedbackfiguremerit, Check User Guide for details
		input  wire [5:0]                                  i_rxpipe7_localfs,                           //                                       .i_rxpipe7_localfs,                           Check User Guide for details
		input  wire [5:0]                                  i_rxpipe7_locallf,                           //                                       .i_rxpipe7_locallf,                           Check User Guide for details
		input  wire                                        i_rxpipe7_localtxcoefficientsvalid,          //                                       .i_rxpipe7_localtxcoefficientsvalid,          Check User Guide for details
		input  wire [17:0]                                 i_rxpipe7_localtxpresetcoefficients,         //                                       .i_rxpipe7_localtxpresetcoefficients,         Check User Guide for details
		input  wire [7:0]                                  i_rxpipe7_p2m_bus,                           //                                       .i_rxpipe7_p2m_bus,                           Check User Guide for details
		input  wire                                        i_rxpipe7_pclkchangeok,                      //                                       .i_rxpipe7_pclkchangeok,                      Check User Guide for details
		input  wire                                        i_rxpipe7_phystatus,                         //                                       .i_rxpipe7_phystatus,                         Check User Guide for details
		input  wire [39:0]                                 i_rxpipe7_rxdata,                            //                                       .i_rxpipe7_rxdata,                            Check User Guide for details
		input  wire [3:0]                                  i_rxpipe7_rxdatak,                           //                                       .i_rxpipe7_rxdatak,                           Check User Guide for details
		input  wire                                        i_rxpipe7_rxdatavalid,                       //                                       .i_rxpipe7_rxdatavalid,                       Check User Guide for details
		input  wire                                        i_rxpipe7_rxelecidlea,                       //                                       .i_rxpipe7_rxelecidlea,                       Check User Guide for details
		input  wire                                        i_rxpipe7_rxstandbystatus,                   //                                       .i_rxpipe7_rxstandbystatus,                   Check User Guide for details
		input  wire                                        i_rxpipe7_rxstartblock,                      //                                       .i_rxpipe7_rxstartblock,                      Check User Guide for details
		input  wire [2:0]                                  i_rxpipe7_rxstatus,                          //                                       .i_rxpipe7_rxstatus,                          Check User Guide for details
		input  wire [3:0]                                  i_rxpipe7_rxsyncheader,                      //                                       .i_rxpipe7_rxsyncheader,                      Check User Guide for details
		input  wire                                        i_rxpipe7_rxvalid,                           //                                       .i_rxpipe7_rxvalid,                           Check User Guide for details
		output wire                                        o_txpipe7_asyncpowerchangeack,               //                                       .o_txpipe7_asyncpowerchangeack,               Check User Guide for details
		output wire                                        o_txpipe7_blockaligncontrol,                 //                                       .o_txpipe7_blockaligncontrol,                 Check User Guide for details
		output wire                                        o_txpipe7_cfg_hw_auto_sp_dis,                //                                       .o_txpipe7_cfg_hw_auto_sp_dis,                Check User Guide for details
		output wire                                        o_txpipe7_dirchange,                         //                                       .o_txpipe7_dirchange,                         Check User Guide for details
		output wire                                        o_txpipe7_ebuf_mode,                         //                                       .o_txpipe7_ebuf_mode,                         Check User Guide for details
		output wire                                        o_txpipe7_encodedecodebypass,                //                                       .o_txpipe7_encodedecodebypass,                Check User Guide for details
		output wire [5:0]                                  o_txpipe7_fs,                                //                                       .o_txpipe7_fs,                                Check User Guide for details
		output wire                                        o_txpipe7_getlocalpresetcoefficients,        //                                       .o_txpipe7_getlocalpresetcoefficients,        Check User Guide for details
		output wire                                        o_txpipe7_invalidrequest,                    //                                       .o_txpipe7_invalidrequest,                    Check User Guide for details
		output wire [5:0]                                  o_txpipe7_lf,                                //                                       .o_txpipe7_lf,                                Check User Guide for details
		output wire [4:0]                                  o_txpipe7_localpresetindex,                  //                                       .o_txpipe7_localpresetindex,                  Check User Guide for details
		output wire                                        o_txpipe7_lowpin_nt,                         //                                       .o_txpipe7_lowpin_nt,                         Check User Guide for details
		output wire [7:0]                                  o_txpipe7_m2p_bus,                           //                                       .o_txpipe7_m2p_bus,                           Check User Guide for details
		output wire [2:0]                                  o_txpipe7_pclk_rate,                         //                                       .o_txpipe7_pclk_rate,                         Check User Guide for details
		output wire                                        o_txpipe7_pclkchangeack,                     //                                       .o_txpipe7_pclkchangeack,                     Check User Guide for details
		output wire [3:0]                                  o_txpipe7_phy_mode_nt,                       //                                       .o_txpipe7_phy_mode_nt,                       Check User Guide for details
		output wire [3:0]                                  o_txpipe7_powerdown,                         //                                       .o_txpipe7_powerdown,                         Check User Guide for details
		output wire [2:0]                                  o_txpipe7_rate,                              //                                       .o_txpipe7_rate,                              Check User Guide for details
		output wire                                        o_txpipe7_rxelecidle_disable_a,              //                                       .o_txpipe7_rxelecidle_disable_a,              Check User Guide for details
		output wire                                        o_txpipe7_rxeqclr,                           //                                       .o_txpipe7_rxeqclr,                           Check User Guide for details
		output wire                                        o_txpipe7_rxeqeval,                          //                                       .o_txpipe7_rxeqeval,                          Check User Guide for details
		output wire                                        o_txpipe7_rxeqinprogress,                    //                                       .o_txpipe7_rxeqinprogress,                    Check User Guide for details
		output wire                                        o_txpipe7_rxeqtraining,                      //                                       .o_txpipe7_rxeqtraining,                      Check User Guide for details
		output wire                                        o_txpipe7_rxpolarity,                        //                                       .o_txpipe7_rxpolarity,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe7_rxpresethint,                      //                                       .o_txpipe7_rxpresethint,                      Check User Guide for details
		output wire                                        o_txpipe7_rxstandby,                         //                                       .o_txpipe7_rxstandby,                         Check User Guide for details
		output wire                                        o_txpipe7_rxtermination,                     //                                       .o_txpipe7_rxtermination,                     Check User Guide for details
		output wire                                        o_txpipe7_srisenable,                        //                                       .o_txpipe7_srisenable,                        Check User Guide for details
		output wire                                        o_txpipe7_txcmnmode_disable_a,               //                                       .o_txpipe7_txcmnmode_disable_a,               Check User Guide for details
		output wire                                        o_txpipe7_txcompliance,                      //                                       .o_txpipe7_txcompliance,                      Check User Guide for details
		output wire [39:0]                                 o_txpipe7_txdata,                            //                                       .o_txpipe7_txdata,                            Check User Guide for details
		output wire [3:0]                                  o_txpipe7_txdatak,                           //                                       .o_txpipe7_txdatak,                           Check User Guide for details
		output wire                                        o_txpipe7_txdatavalid,                       //                                       .o_txpipe7_txdatavalid,                       Check User Guide for details
		output wire [17:0]                                 o_txpipe7_txdeemph,                          //                                       .o_txpipe7_txdeemph,                          Check User Guide for details
		output wire                                        o_txpipe7_txdtctrx_lb,                       //                                       .o_txpipe7_txdtctrx_lb,                       Check User Guide for details
		output wire                                        o_txpipe7_txelecidle,                        //                                       .o_txpipe7_txelecidle,                        Check User Guide for details
		output wire [2:0]                                  o_txpipe7_txmargin,                          //                                       .o_txpipe7_txmargin,                          Check User Guide for details
		output wire                                        o_txpipe7_txoneszeros,                       //                                       .o_txpipe7_txoneszeros,                       Check User Guide for details
		output wire                                        o_txpipe7_txstartblock,                      //                                       .o_txpipe7_txstartblock,                      Check User Guide for details
		output wire                                        o_txpipe7_txswing,                           //                                       .o_txpipe7_txswing,                           Check User Guide for details
		output wire [3:0]                                  o_txpipe7_txsyncheader,                      //                                       .o_txpipe7_txsyncheader,                      Check User Guide for details
		output wire [2:0]                                  o_txpipe7_width,                             //                                       .o_txpipe7_width,                             Check User Guide for details
		input  wire                                        i_pin_perst_n,                               //                                       .i_pin_perst_n,                               Check User Guide for details
		input  wire                                        i_hio_ch0_lavmm_clk,                         //                    i_hio_ch0_lavmm_clk.clk
		input  wire                                        i_hio_ch0_lavmm_rstn,                        //                   i_hio_ch0_lavmm_rstn.reset
		input  wire [20:0]                                 i_hio_ch0_lavmm_addr,                        //                          hio_ch0_lavmm.address
		input  wire [3:0]                                  i_hio_ch0_lavmm_be,                          //                                       .byteenable
		output wire                                        o_hio_ch0_lavmm_rdata_valid,                 //                                       .readdatavalid
		input  wire                                        i_hio_ch0_lavmm_read,                        //                                       .read
		input  wire                                        i_hio_ch0_lavmm_write,                       //                                       .write
		output wire [31:0]                                 o_hio_ch0_lavmm_rdata,                       //                                       .readdata
		input  wire [31:0]                                 i_hio_ch0_lavmm_wdata,                       //                                       .writedata
		output wire                                        o_hio_ch0_lavmm_waitreq,                     //                                       .waitrequest
		input  wire                                        i_hio_ch0_pld_rx_clk_in_row_clk,             //        i_hio_ch0_pld_rx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch0_pld_tx_clk_in_row_clk,             //        i_hio_ch0_pld_tx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch0_det_lat_rx_dl_clk,                 //            i_hio_ch0_det_lat_rx_dl_clk.clk
		input  wire                                        i_hio_ch0_det_lat_rx_mux_select,             //        i_hio_ch0_det_lat_rx_mux_select.clk
		input  wire                                        i_hio_ch0_det_lat_rx_sclk_flop,              //         i_hio_ch0_det_lat_rx_sclk_flop.clk
		input  wire                                        i_hio_ch0_det_lat_rx_sclk_gen_clk,           //      i_hio_ch0_det_lat_rx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch0_det_lat_rx_trig_flop,              //         i_hio_ch0_det_lat_rx_trig_flop.clk
		input  wire                                        i_hio_ch0_det_lat_sampling_clk,              //         i_hio_ch0_det_lat_sampling_clk.clk
		input  wire                                        i_hio_ch0_det_lat_tx_dl_clk,                 //            i_hio_ch0_det_lat_tx_dl_clk.clk
		input  wire                                        i_hio_ch0_det_lat_tx_mux_select,             //        i_hio_ch0_det_lat_tx_mux_select.clk
		input  wire                                        i_hio_ch0_det_lat_tx_sclk_flop,              //         i_hio_ch0_det_lat_tx_sclk_flop.clk
		input  wire                                        i_hio_ch0_det_lat_tx_sclk_gen_clk,           //      i_hio_ch0_det_lat_tx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch0_det_lat_tx_trig_flop,              //         i_hio_ch0_det_lat_tx_trig_flop.clk
		output wire                                        o_hio_ch0_user_rx_clk1_clk,                  //             o_hio_ch0_user_rx_clk1_clk.clk
		output wire                                        o_hio_ch0_user_rx_clk2_clk,                  //             o_hio_ch0_user_rx_clk2_clk.clk
		output wire                                        o_hio_ch0_user_tx_clk1_clk,                  //             o_hio_ch0_user_tx_clk1_clk.clk
		output wire                                        o_hio_ch0_user_tx_clk2_clk,                  //             o_hio_ch0_user_tx_clk2_clk.clk
		output wire                                        o_hio_ch0_ux_chnl_refclk_mux,                //           o_hio_ch0_ux_chnl_refclk_mux.clk
		output wire                                        o_hio_ch0_det_lat_rx_async_dl_sync,          //     o_hio_ch0_det_lat_rx_async_dl_sync.clk
		output wire                                        o_hio_ch0_det_lat_rx_async_pulse,            //       o_hio_ch0_det_lat_rx_async_pulse.clk
		output wire                                        o_hio_ch0_det_lat_rx_async_sample_sync,      // o_hio_ch0_det_lat_rx_async_sample_sync.clk
		output wire                                        o_hio_ch0_det_lat_rx_sclk_sample_sync,       //  o_hio_ch0_det_lat_rx_sclk_sample_sync.clk
		output wire                                        o_hio_ch0_det_lat_rx_trig_sample_sync,       //  o_hio_ch0_det_lat_rx_trig_sample_sync.clk
		output wire                                        o_hio_ch0_det_lat_tx_async_dl_sync,          //     o_hio_ch0_det_lat_tx_async_dl_sync.clk
		output wire                                        o_hio_ch0_det_lat_tx_async_pulse,            //       o_hio_ch0_det_lat_tx_async_pulse.clk
		output wire                                        o_hio_ch0_det_lat_tx_async_sample_sync,      // o_hio_ch0_det_lat_tx_async_sample_sync.clk
		output wire                                        o_hio_ch0_det_lat_tx_sclk_sample_sync,       //  o_hio_ch0_det_lat_tx_sclk_sample_sync.clk
		output wire                                        o_hio_ch0_det_lat_tx_trig_sample_sync,       //  o_hio_ch0_det_lat_tx_trig_sample_sync.clk
		output wire                                        o_hio_ch0_xcvrif_rx_latency_pulse,           //      o_hio_ch0_xcvrif_rx_latency_pulse.clk
		output wire                                        o_hio_ch0_xcvrif_tx_latency_pulse,           //      o_hio_ch0_xcvrif_tx_latency_pulse.clk
		input  wire                                        i_hio_ch1_lavmm_clk,                         //                    i_hio_ch1_lavmm_clk.clk
		input  wire                                        i_hio_ch1_lavmm_rstn,                        //                   i_hio_ch1_lavmm_rstn.reset
		input  wire [20:0]                                 i_hio_ch1_lavmm_addr,                        //                          hio_ch1_lavmm.address
		input  wire [3:0]                                  i_hio_ch1_lavmm_be,                          //                                       .byteenable
		output wire                                        o_hio_ch1_lavmm_rdata_valid,                 //                                       .readdatavalid
		input  wire                                        i_hio_ch1_lavmm_read,                        //                                       .read
		input  wire                                        i_hio_ch1_lavmm_write,                       //                                       .write
		output wire [31:0]                                 o_hio_ch1_lavmm_rdata,                       //                                       .readdata
		input  wire [31:0]                                 i_hio_ch1_lavmm_wdata,                       //                                       .writedata
		output wire                                        o_hio_ch1_lavmm_waitreq,                     //                                       .waitrequest
		input  wire                                        i_hio_ch1_pld_rx_clk_in_row_clk,             //        i_hio_ch1_pld_rx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch1_pld_tx_clk_in_row_clk,             //        i_hio_ch1_pld_tx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch1_det_lat_rx_dl_clk,                 //            i_hio_ch1_det_lat_rx_dl_clk.clk
		input  wire                                        i_hio_ch1_det_lat_rx_mux_select,             //        i_hio_ch1_det_lat_rx_mux_select.clk
		input  wire                                        i_hio_ch1_det_lat_rx_sclk_flop,              //         i_hio_ch1_det_lat_rx_sclk_flop.clk
		input  wire                                        i_hio_ch1_det_lat_rx_sclk_gen_clk,           //      i_hio_ch1_det_lat_rx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch1_det_lat_rx_trig_flop,              //         i_hio_ch1_det_lat_rx_trig_flop.clk
		input  wire                                        i_hio_ch1_det_lat_sampling_clk,              //         i_hio_ch1_det_lat_sampling_clk.clk
		input  wire                                        i_hio_ch1_det_lat_tx_dl_clk,                 //            i_hio_ch1_det_lat_tx_dl_clk.clk
		input  wire                                        i_hio_ch1_det_lat_tx_mux_select,             //        i_hio_ch1_det_lat_tx_mux_select.clk
		input  wire                                        i_hio_ch1_det_lat_tx_sclk_flop,              //         i_hio_ch1_det_lat_tx_sclk_flop.clk
		input  wire                                        i_hio_ch1_det_lat_tx_sclk_gen_clk,           //      i_hio_ch1_det_lat_tx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch1_det_lat_tx_trig_flop,              //         i_hio_ch1_det_lat_tx_trig_flop.clk
		output wire                                        o_hio_ch1_user_rx_clk1_clk,                  //             o_hio_ch1_user_rx_clk1_clk.clk
		output wire                                        o_hio_ch1_user_rx_clk2_clk,                  //             o_hio_ch1_user_rx_clk2_clk.clk
		output wire                                        o_hio_ch1_user_tx_clk1_clk,                  //             o_hio_ch1_user_tx_clk1_clk.clk
		output wire                                        o_hio_ch1_user_tx_clk2_clk,                  //             o_hio_ch1_user_tx_clk2_clk.clk
		output wire                                        o_hio_ch1_ux_chnl_refclk_mux,                //           o_hio_ch1_ux_chnl_refclk_mux.clk
		output wire                                        o_hio_ch1_det_lat_rx_async_dl_sync,          //     o_hio_ch1_det_lat_rx_async_dl_sync.clk
		output wire                                        o_hio_ch1_det_lat_rx_async_pulse,            //       o_hio_ch1_det_lat_rx_async_pulse.clk
		output wire                                        o_hio_ch1_det_lat_rx_async_sample_sync,      // o_hio_ch1_det_lat_rx_async_sample_sync.clk
		output wire                                        o_hio_ch1_det_lat_rx_sclk_sample_sync,       //  o_hio_ch1_det_lat_rx_sclk_sample_sync.clk
		output wire                                        o_hio_ch1_det_lat_rx_trig_sample_sync,       //  o_hio_ch1_det_lat_rx_trig_sample_sync.clk
		output wire                                        o_hio_ch1_det_lat_tx_async_dl_sync,          //     o_hio_ch1_det_lat_tx_async_dl_sync.clk
		output wire                                        o_hio_ch1_det_lat_tx_async_pulse,            //       o_hio_ch1_det_lat_tx_async_pulse.clk
		output wire                                        o_hio_ch1_det_lat_tx_async_sample_sync,      // o_hio_ch1_det_lat_tx_async_sample_sync.clk
		output wire                                        o_hio_ch1_det_lat_tx_sclk_sample_sync,       //  o_hio_ch1_det_lat_tx_sclk_sample_sync.clk
		output wire                                        o_hio_ch1_det_lat_tx_trig_sample_sync,       //  o_hio_ch1_det_lat_tx_trig_sample_sync.clk
		output wire                                        o_hio_ch1_xcvrif_rx_latency_pulse,           //      o_hio_ch1_xcvrif_rx_latency_pulse.clk
		output wire                                        o_hio_ch1_xcvrif_tx_latency_pulse,           //      o_hio_ch1_xcvrif_tx_latency_pulse.clk
		input  wire                                        i_hio_ch2_lavmm_clk,                         //                    i_hio_ch2_lavmm_clk.clk
		input  wire                                        i_hio_ch2_lavmm_rstn,                        //                   i_hio_ch2_lavmm_rstn.reset
		input  wire [20:0]                                 i_hio_ch2_lavmm_addr,                        //                          hio_ch2_lavmm.address
		input  wire [3:0]                                  i_hio_ch2_lavmm_be,                          //                                       .byteenable
		output wire                                        o_hio_ch2_lavmm_rdata_valid,                 //                                       .readdatavalid
		input  wire                                        i_hio_ch2_lavmm_read,                        //                                       .read
		input  wire                                        i_hio_ch2_lavmm_write,                       //                                       .write
		output wire [31:0]                                 o_hio_ch2_lavmm_rdata,                       //                                       .readdata
		input  wire [31:0]                                 i_hio_ch2_lavmm_wdata,                       //                                       .writedata
		output wire                                        o_hio_ch2_lavmm_waitreq,                     //                                       .waitrequest
		input  wire                                        i_hio_ch2_pld_rx_clk_in_row_clk,             //        i_hio_ch2_pld_rx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch2_pld_tx_clk_in_row_clk,             //        i_hio_ch2_pld_tx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch2_det_lat_rx_dl_clk,                 //            i_hio_ch2_det_lat_rx_dl_clk.clk
		input  wire                                        i_hio_ch2_det_lat_rx_mux_select,             //        i_hio_ch2_det_lat_rx_mux_select.clk
		input  wire                                        i_hio_ch2_det_lat_rx_sclk_flop,              //         i_hio_ch2_det_lat_rx_sclk_flop.clk
		input  wire                                        i_hio_ch2_det_lat_rx_sclk_gen_clk,           //      i_hio_ch2_det_lat_rx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch2_det_lat_rx_trig_flop,              //         i_hio_ch2_det_lat_rx_trig_flop.clk
		input  wire                                        i_hio_ch2_det_lat_sampling_clk,              //         i_hio_ch2_det_lat_sampling_clk.clk
		input  wire                                        i_hio_ch2_det_lat_tx_dl_clk,                 //            i_hio_ch2_det_lat_tx_dl_clk.clk
		input  wire                                        i_hio_ch2_det_lat_tx_mux_select,             //        i_hio_ch2_det_lat_tx_mux_select.clk
		input  wire                                        i_hio_ch2_det_lat_tx_sclk_flop,              //         i_hio_ch2_det_lat_tx_sclk_flop.clk
		input  wire                                        i_hio_ch2_det_lat_tx_sclk_gen_clk,           //      i_hio_ch2_det_lat_tx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch2_det_lat_tx_trig_flop,              //         i_hio_ch2_det_lat_tx_trig_flop.clk
		output wire                                        o_hio_ch2_user_rx_clk1_clk,                  //             o_hio_ch2_user_rx_clk1_clk.clk
		output wire                                        o_hio_ch2_user_rx_clk2_clk,                  //             o_hio_ch2_user_rx_clk2_clk.clk
		output wire                                        o_hio_ch2_user_tx_clk1_clk,                  //             o_hio_ch2_user_tx_clk1_clk.clk
		output wire                                        o_hio_ch2_user_tx_clk2_clk,                  //             o_hio_ch2_user_tx_clk2_clk.clk
		output wire                                        o_hio_ch2_ux_chnl_refclk_mux,                //           o_hio_ch2_ux_chnl_refclk_mux.clk
		output wire                                        o_hio_ch2_det_lat_rx_async_dl_sync,          //     o_hio_ch2_det_lat_rx_async_dl_sync.clk
		output wire                                        o_hio_ch2_det_lat_rx_async_pulse,            //       o_hio_ch2_det_lat_rx_async_pulse.clk
		output wire                                        o_hio_ch2_det_lat_rx_async_sample_sync,      // o_hio_ch2_det_lat_rx_async_sample_sync.clk
		output wire                                        o_hio_ch2_det_lat_rx_sclk_sample_sync,       //  o_hio_ch2_det_lat_rx_sclk_sample_sync.clk
		output wire                                        o_hio_ch2_det_lat_rx_trig_sample_sync,       //  o_hio_ch2_det_lat_rx_trig_sample_sync.clk
		output wire                                        o_hio_ch2_det_lat_tx_async_dl_sync,          //     o_hio_ch2_det_lat_tx_async_dl_sync.clk
		output wire                                        o_hio_ch2_det_lat_tx_async_pulse,            //       o_hio_ch2_det_lat_tx_async_pulse.clk
		output wire                                        o_hio_ch2_det_lat_tx_async_sample_sync,      // o_hio_ch2_det_lat_tx_async_sample_sync.clk
		output wire                                        o_hio_ch2_det_lat_tx_sclk_sample_sync,       //  o_hio_ch2_det_lat_tx_sclk_sample_sync.clk
		output wire                                        o_hio_ch2_det_lat_tx_trig_sample_sync,       //  o_hio_ch2_det_lat_tx_trig_sample_sync.clk
		output wire                                        o_hio_ch2_xcvrif_rx_latency_pulse,           //      o_hio_ch2_xcvrif_rx_latency_pulse.clk
		output wire                                        o_hio_ch2_xcvrif_tx_latency_pulse,           //      o_hio_ch2_xcvrif_tx_latency_pulse.clk
		input  wire                                        i_hio_ch3_lavmm_clk,                         //                    i_hio_ch3_lavmm_clk.clk
		input  wire                                        i_hio_ch3_lavmm_rstn,                        //                   i_hio_ch3_lavmm_rstn.reset
		input  wire [20:0]                                 i_hio_ch3_lavmm_addr,                        //                          hio_ch3_lavmm.address
		input  wire [3:0]                                  i_hio_ch3_lavmm_be,                          //                                       .byteenable
		output wire                                        o_hio_ch3_lavmm_rdata_valid,                 //                                       .readdatavalid
		input  wire                                        i_hio_ch3_lavmm_read,                        //                                       .read
		input  wire                                        i_hio_ch3_lavmm_write,                       //                                       .write
		output wire [31:0]                                 o_hio_ch3_lavmm_rdata,                       //                                       .readdata
		input  wire [31:0]                                 i_hio_ch3_lavmm_wdata,                       //                                       .writedata
		output wire                                        o_hio_ch3_lavmm_waitreq,                     //                                       .waitrequest
		input  wire                                        i_hio_ch3_pld_rx_clk_in_row_clk,             //        i_hio_ch3_pld_rx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch3_pld_tx_clk_in_row_clk,             //        i_hio_ch3_pld_tx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch3_det_lat_rx_dl_clk,                 //            i_hio_ch3_det_lat_rx_dl_clk.clk
		input  wire                                        i_hio_ch3_det_lat_rx_mux_select,             //        i_hio_ch3_det_lat_rx_mux_select.clk
		input  wire                                        i_hio_ch3_det_lat_rx_sclk_flop,              //         i_hio_ch3_det_lat_rx_sclk_flop.clk
		input  wire                                        i_hio_ch3_det_lat_rx_sclk_gen_clk,           //      i_hio_ch3_det_lat_rx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch3_det_lat_rx_trig_flop,              //         i_hio_ch3_det_lat_rx_trig_flop.clk
		input  wire                                        i_hio_ch3_det_lat_sampling_clk,              //         i_hio_ch3_det_lat_sampling_clk.clk
		input  wire                                        i_hio_ch3_det_lat_tx_dl_clk,                 //            i_hio_ch3_det_lat_tx_dl_clk.clk
		input  wire                                        i_hio_ch3_det_lat_tx_mux_select,             //        i_hio_ch3_det_lat_tx_mux_select.clk
		input  wire                                        i_hio_ch3_det_lat_tx_sclk_flop,              //         i_hio_ch3_det_lat_tx_sclk_flop.clk
		input  wire                                        i_hio_ch3_det_lat_tx_sclk_gen_clk,           //      i_hio_ch3_det_lat_tx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch3_det_lat_tx_trig_flop,              //         i_hio_ch3_det_lat_tx_trig_flop.clk
		output wire                                        o_hio_ch3_user_rx_clk1_clk,                  //             o_hio_ch3_user_rx_clk1_clk.clk
		output wire                                        o_hio_ch3_user_rx_clk2_clk,                  //             o_hio_ch3_user_rx_clk2_clk.clk
		output wire                                        o_hio_ch3_user_tx_clk1_clk,                  //             o_hio_ch3_user_tx_clk1_clk.clk
		output wire                                        o_hio_ch3_user_tx_clk2_clk,                  //             o_hio_ch3_user_tx_clk2_clk.clk
		output wire                                        o_hio_ch3_ux_chnl_refclk_mux,                //           o_hio_ch3_ux_chnl_refclk_mux.clk
		output wire                                        o_hio_ch3_det_lat_rx_async_dl_sync,          //     o_hio_ch3_det_lat_rx_async_dl_sync.clk
		output wire                                        o_hio_ch3_det_lat_rx_async_pulse,            //       o_hio_ch3_det_lat_rx_async_pulse.clk
		output wire                                        o_hio_ch3_det_lat_rx_async_sample_sync,      // o_hio_ch3_det_lat_rx_async_sample_sync.clk
		output wire                                        o_hio_ch3_det_lat_rx_sclk_sample_sync,       //  o_hio_ch3_det_lat_rx_sclk_sample_sync.clk
		output wire                                        o_hio_ch3_det_lat_rx_trig_sample_sync,       //  o_hio_ch3_det_lat_rx_trig_sample_sync.clk
		output wire                                        o_hio_ch3_det_lat_tx_async_dl_sync,          //     o_hio_ch3_det_lat_tx_async_dl_sync.clk
		output wire                                        o_hio_ch3_det_lat_tx_async_pulse,            //       o_hio_ch3_det_lat_tx_async_pulse.clk
		output wire                                        o_hio_ch3_det_lat_tx_async_sample_sync,      // o_hio_ch3_det_lat_tx_async_sample_sync.clk
		output wire                                        o_hio_ch3_det_lat_tx_sclk_sample_sync,       //  o_hio_ch3_det_lat_tx_sclk_sample_sync.clk
		output wire                                        o_hio_ch3_det_lat_tx_trig_sample_sync,       //  o_hio_ch3_det_lat_tx_trig_sample_sync.clk
		output wire                                        o_hio_ch3_xcvrif_rx_latency_pulse,           //      o_hio_ch3_xcvrif_rx_latency_pulse.clk
		output wire                                        o_hio_ch3_xcvrif_tx_latency_pulse,           //      o_hio_ch3_xcvrif_tx_latency_pulse.clk
		input  wire                                        i_hio_ch4_lavmm_clk,                         //                    i_hio_ch4_lavmm_clk.clk
		input  wire                                        i_hio_ch4_lavmm_rstn,                        //                   i_hio_ch4_lavmm_rstn.reset
		input  wire [20:0]                                 i_hio_ch4_lavmm_addr,                        //                          hio_ch4_lavmm.address
		input  wire [3:0]                                  i_hio_ch4_lavmm_be,                          //                                       .byteenable
		output wire                                        o_hio_ch4_lavmm_rdata_valid,                 //                                       .readdatavalid
		input  wire                                        i_hio_ch4_lavmm_read,                        //                                       .read
		input  wire                                        i_hio_ch4_lavmm_write,                       //                                       .write
		output wire [31:0]                                 o_hio_ch4_lavmm_rdata,                       //                                       .readdata
		input  wire [31:0]                                 i_hio_ch4_lavmm_wdata,                       //                                       .writedata
		output wire                                        o_hio_ch4_lavmm_waitreq,                     //                                       .waitrequest
		input  wire                                        i_hio_ch4_pld_rx_clk_in_row_clk,             //        i_hio_ch4_pld_rx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch4_pld_tx_clk_in_row_clk,             //        i_hio_ch4_pld_tx_clk_in_row_clk.clk
		input  wire                                        i_hio_ch4_det_lat_rx_dl_clk,                 //            i_hio_ch4_det_lat_rx_dl_clk.clk
		input  wire                                        i_hio_ch4_det_lat_rx_mux_select,             //        i_hio_ch4_det_lat_rx_mux_select.clk
		input  wire                                        i_hio_ch4_det_lat_rx_sclk_flop,              //         i_hio_ch4_det_lat_rx_sclk_flop.clk
		input  wire                                        i_hio_ch4_det_lat_rx_sclk_gen_clk,           //      i_hio_ch4_det_lat_rx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch4_det_lat_rx_trig_flop,              //         i_hio_ch4_det_lat_rx_trig_flop.clk
		input  wire                                        i_hio_ch4_det_lat_sampling_clk,              //         i_hio_ch4_det_lat_sampling_clk.clk
		input  wire                                        i_hio_ch4_det_lat_tx_dl_clk,                 //            i_hio_ch4_det_lat_tx_dl_clk.clk
		input  wire                                        i_hio_ch4_det_lat_tx_mux_select,             //        i_hio_ch4_det_lat_tx_mux_select.clk
		input  wire                                        i_hio_ch4_det_lat_tx_sclk_flop,              //         i_hio_ch4_det_lat_tx_sclk_flop.clk
		input  wire                                        i_hio_ch4_det_lat_tx_sclk_gen_clk,           //      i_hio_ch4_det_lat_tx_sclk_gen_clk.clk
		input  wire                                        i_hio_ch4_det_lat_tx_trig_flop,              //         i_hio_ch4_det_lat_tx_trig_flop.clk
		output wire                                        o_hio_ch4_user_rx_clk1_clk,                  //             o_hio_ch4_user_rx_clk1_clk.clk
		output wire                                        o_hio_ch4_user_rx_clk2_clk,                  //             o_hio_ch4_user_rx_clk2_clk.clk
		output wire                                        o_hio_ch4_user_tx_clk1_clk,                  //             o_hio_ch4_user_tx_clk1_clk.clk
		output wire                                        o_hio_ch4_user_tx_clk2_clk,                  //             o_hio_ch4_user_tx_clk2_clk.clk
		output wire                                        o_hio_ch4_ux_chnl_refclk_mux,                //           o_hio_ch4_ux_chnl_refclk_mux.clk
		output wire                                        o_hio_ch4_det_lat_rx_async_dl_sync,          //     o_hio_ch4_det_lat_rx_async_dl_sync.clk
		output wire                                        o_hio_ch4_det_lat_rx_async_pulse,            //       o_hio_ch4_det_lat_rx_async_pulse.clk
		output wire                                        o_hio_ch4_det_lat_rx_async_sample_sync,      // o_hio_ch4_det_lat_rx_async_sample_sync.clk
		output wire                                        o_hio_ch4_det_lat_rx_sclk_sample_sync,       //  o_hio_ch4_det_lat_rx_sclk_sample_sync.clk
		output wire                                        o_hio_ch4_det_lat_rx_trig_sample_sync,       //  o_hio_ch4_det_lat_rx_trig_sample_sync.clk
		output wire                                        o_hio_ch4_det_lat_tx_async_dl_sync,          //     o_hio_ch4_det_lat_tx_async_dl_sync.clk
		output wire                                        o_hio_ch4_det_lat_tx_async_pulse,            //       o_hio_ch4_det_lat_tx_async_pulse.clk
		output wire                                        o_hio_ch4_det_lat_tx_async_sample_sync,      // o_hio_ch4_det_lat_tx_async_sample_sync.clk
		output wire                                        o_hio_ch4_det_lat_tx_sclk_sample_sync,       //  o_hio_ch4_det_lat_tx_sclk_sample_sync.clk
		output wire                                        o_hio_ch4_det_lat_tx_trig_sample_sync,       //  o_hio_ch4_det_lat_tx_trig_sample_sync.clk
		output wire                                        o_hio_ch4_xcvrif_rx_latency_pulse,           //      o_hio_ch4_xcvrif_rx_latency_pulse.clk
		output wire                                        o_hio_ch4_xcvrif_tx_latency_pulse            //      o_hio_ch4_xcvrif_tx_latency_pulse.clk
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (ch0_pcs_l_tx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_pcs_l_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch0_pcs_l_rx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_pcs_l_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_loopback_mode_atom != "CH0_LOOPBACK_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_dyn_tx_mux_atom != "CH0_DYN_TX_MUX_ETHPCS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_dyn_tx_mux_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_error_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_error_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_rx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_tx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_mode_atom != "CH0_FEC_MODE_RSFEC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_pcs_l_tx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_pcs_l_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch1_pcs_l_rx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_pcs_l_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_loopback_mode_atom != "CH1_LOOPBACK_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_dyn_tx_mux_atom != "CH1_DYN_TX_MUX_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_dyn_tx_mux_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_error_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_error_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_rx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_tx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_mode_atom != "CH1_FEC_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_pcs_l_tx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_pcs_l_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch2_pcs_l_rx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_pcs_l_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_loopback_mode_atom != "CH2_LOOPBACK_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_dyn_tx_mux_atom != "CH2_DYN_TX_MUX_ETHPCS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_dyn_tx_mux_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_error_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_error_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_rx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_tx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_mode_atom != "CH2_FEC_MODE_RSFEC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_pcs_l_tx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_pcs_l_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch3_pcs_l_rx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_pcs_l_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_loopback_mode_atom != "CH3_LOOPBACK_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_dyn_tx_mux_atom != "CH3_DYN_TX_MUX_DESKEW")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_dyn_tx_mux_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_error_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_error_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_rx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_tx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_mode_atom != "CH3_FEC_MODE_RSFEC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_rx_prbs_monitor_en_atom != "CH0_RX_PRBS_MONITOR_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_rx_prbs_monitor_en_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_rx_prbs_monitor_en_atom != "CH1_RX_PRBS_MONITOR_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_rx_prbs_monitor_en_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_rx_prbs_monitor_en_atom != "CH2_RX_PRBS_MONITOR_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_rx_prbs_monitor_en_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_rx_prbs_monitor_en_atom != "CH3_RX_PRBS_MONITOR_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_rx_prbs_monitor_en_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_prbs_gen_en_atom != "CH0_TX_PRBS_GEN_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_prbs_gen_en_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_prbs_gen_en_atom != "CH1_TX_PRBS_GEN_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_prbs_gen_en_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_prbs_gen_en_atom != "CH2_TX_PRBS_GEN_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_prbs_gen_en_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_prbs_gen_en_atom != "CH3_TX_PRBS_GEN_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_prbs_gen_en_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_user1_clk_mux_dynamic_sel_atom != "CH0_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_user2_clk_mux_dynamic_sel_atom != "CH0_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_user1_clk_mux_dynamic_sel_atom != "CH0_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_user2_clk_mux_dynamic_sel_atom != "CH0_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_user1_clk_mux_dynamic_sel_atom != "CH1_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_user2_clk_mux_dynamic_sel_atom != "CH1_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_user1_clk_mux_dynamic_sel_atom != "CH1_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_user2_clk_mux_dynamic_sel_atom != "CH1_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_user1_clk_mux_dynamic_sel_atom != "CH2_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_user2_clk_mux_dynamic_sel_atom != "CH2_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_user1_clk_mux_dynamic_sel_atom != "CH2_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_user2_clk_mux_dynamic_sel_atom != "CH2_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_user1_clk_mux_dynamic_sel_atom != "CH3_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_user2_clk_mux_dynamic_sel_atom != "CH3_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_user1_clk_mux_dynamic_sel_atom != "CH3_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_user2_clk_mux_dynamic_sel_atom != "CH3_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch0_pcie_mode_atom != "CH0_PCIE_MODE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_pcie_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_pcie_mode_atom != "CH1_PCIE_MODE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_pcie_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_pcie_mode_atom != "CH2_PCIE_MODE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_pcie_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_pcie_mode_atom != "CH3_PCIE_MODE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_pcie_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_rx_protocol_hint_atom != "CH0_RX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_rx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_rx_protocol_hint_atom != "CH1_RX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_rx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_rx_protocol_hint_atom != "CH2_RX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_rx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_rx_protocol_hint_atom != "CH3_RX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_rx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch0_clkrx_refclk_cssm_fw_control_atom != "CH0_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_clkrx_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch1_clkrx_refclk_cssm_fw_control_atom != "CH1_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_clkrx_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch2_clkrx_refclk_cssm_fw_control_atom != "CH2_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_clkrx_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch3_clkrx_refclk_cssm_fw_control_atom != "CH3_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_clkrx_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch0_clkrx_refclk_sector_specifies_refclk_ready_atom != "CH0_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_clkrx_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch1_clkrx_refclk_sector_specifies_refclk_ready_atom != "CH1_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_clkrx_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch2_clkrx_refclk_sector_specifies_refclk_ready_atom != "CH2_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_clkrx_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch3_clkrx_refclk_sector_specifies_refclk_ready_atom != "CH3_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_clkrx_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch0_local_refclk_cssm_fw_control_atom != "CH0_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_local_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch1_local_refclk_cssm_fw_control_atom != "CH1_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_local_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch2_local_refclk_cssm_fw_control_atom != "CH2_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_local_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch3_local_refclk_cssm_fw_control_atom != "CH3_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_local_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch0_local_refclk_sector_specifies_refclk_ready_atom != "CH0_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_local_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch1_local_refclk_sector_specifies_refclk_ready_atom != "CH1_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_local_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch2_local_refclk_sector_specifies_refclk_ready_atom != "CH2_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_local_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch3_local_refclk_sector_specifies_refclk_ready_atom != "CH3_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_local_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_bonding_category_atom != "CH0_TX_BONDING_CATEGORY_BONDING_LEADER")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_bonding_category_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_bonding_category_atom != "CH1_TX_BONDING_CATEGORY_BONDING_FOLLOWER")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_bonding_category_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_bonding_category_atom != "CH2_TX_BONDING_CATEGORY_BONDING_FOLLOWER")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_bonding_category_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_bonding_category_atom != "CH3_TX_BONDING_CATEGORY_BONDING_FOLLOWER")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_bonding_category_atom_check ( .error(1'b1) );
		end
		if (hal_num_of_lanes_hwtcl != 4)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					hal_num_of_lanes_hwtcl_check ( .error(1'b1) );
		end
		if (ch0_duplex_mode_atom != "CH0_DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_fec_spec_atom != "CH0_FEC_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fec_spec_atom_check ( .error(1'b1) );
		end
		if (ch0_fracture_atom != "CH0_FRACTURE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_fracture_atom_check ( .error(1'b1) );
		end
		if (ch0_dr_enabled_atom != "CH0_DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch0_sup_mode_atom != "CH0_SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_sup_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_sim_mode_atom != "CH0_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_duplex_mode_atom != "CH1_DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_fec_spec_atom != "CH1_FEC_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fec_spec_atom_check ( .error(1'b1) );
		end
		if (ch1_fracture_atom != "CH1_FRACTURE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_fracture_atom_check ( .error(1'b1) );
		end
		if (ch1_dr_enabled_atom != "CH1_DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch1_sup_mode_atom != "CH1_SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_sup_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_sim_mode_atom != "CH1_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_duplex_mode_atom != "CH2_DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_fec_spec_atom != "CH2_FEC_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fec_spec_atom_check ( .error(1'b1) );
		end
		if (ch2_fracture_atom != "CH2_FRACTURE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_fracture_atom_check ( .error(1'b1) );
		end
		if (ch2_dr_enabled_atom != "CH2_DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch2_sup_mode_atom != "CH2_SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_sup_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_sim_mode_atom != "CH2_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_duplex_mode_atom != "CH3_DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_fec_spec_atom != "CH3_FEC_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fec_spec_atom_check ( .error(1'b1) );
		end
		if (ch3_fracture_atom != "CH3_FRACTURE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_fracture_atom_check ( .error(1'b1) );
		end
		if (ch3_dr_enabled_atom != "CH3_DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch3_sup_mode_atom != "CH3_SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_sup_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_sim_mode_atom != "CH3_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_tx_preloaded_hardware_configs_atom != "CH0_TX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_tx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_rx_preloaded_hardware_configs_atom != "CH0_RX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_rx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch0_lc_postdiv_sel_atom != "CH0_LC_POSTDIV_SEL_SYNTH2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_lc_postdiv_sel_atom_check ( .error(1'b1) );
		end
		if (ch0_sequencer_reg_en_atom != "CH0_SEQUENCER_REG_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_sequencer_reg_en_atom_check ( .error(1'b1) );
		end
		if (ch0_rst_mux_static_sel_atom != "CH0_RST_MUX_STATIC_SEL_HRC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rst_mux_static_sel_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_tx_prbs_pattern_atom != 4'b0000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_tx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_rx_prbs_pattern_atom != 4'b0000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_rx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_tx_user_clk_only_mode_atom != "CH0_TX_USER_CLK_ONLY_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_tx_user_clk_only_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_tx_width_atom != "CH0_TX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_tx_width_atom_check ( .error(1'b1) );
		end
		if (ch0_xcvr_rx_width_atom != "CH0_RX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_xcvr_rx_width_atom_check ( .error(1'b1) );
		end
		if (ch0_phy_loopback_mode_atom != "CH0_LOOPBACK_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_phy_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_flux_mode_atom != "CH0_FLUX_MODE_FLUX_MODE_BYPASS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_flux_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_sim_mode_atom != "CH0_TX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_sim_mode_atom != "CH0_RX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_dl_enable_atom != "CH0_TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_dl_enable_atom != "CH0_RX_DL_ENABLE_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_fec_type_used_atom != "CH0_RX_FEC_TYPE_USED_RS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_fec_type_used_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_tx_preloaded_hardware_configs_atom != "CH1_TX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_tx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_rx_preloaded_hardware_configs_atom != "CH1_RX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_rx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch1_lc_postdiv_sel_atom != "CH1_LC_POSTDIV_SEL_SYNTH2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_lc_postdiv_sel_atom_check ( .error(1'b1) );
		end
		if (ch1_sequencer_reg_en_atom != "CH1_SEQUENCER_REG_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_sequencer_reg_en_atom_check ( .error(1'b1) );
		end
		if (ch1_rst_mux_static_sel_atom != "CH1_RST_MUX_STATIC_SEL_HRC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rst_mux_static_sel_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_tx_prbs_pattern_atom != 4'b0000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_tx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_rx_prbs_pattern_atom != 4'b0001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_rx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_tx_user_clk_only_mode_atom != "CH1_TX_USER_CLK_ONLY_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_tx_user_clk_only_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_tx_width_atom != "CH1_TX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_tx_width_atom_check ( .error(1'b1) );
		end
		if (ch1_xcvr_rx_width_atom != "CH1_RX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_xcvr_rx_width_atom_check ( .error(1'b1) );
		end
		if (ch1_phy_loopback_mode_atom != "CH1_LOOPBACK_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_phy_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_flux_mode_atom != "CH1_FLUX_MODE_FLUX_MODE_BYPASS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_flux_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_sim_mode_atom != "CH1_TX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_sim_mode_atom != "CH1_RX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_dl_enable_atom != "CH1_TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_dl_enable_atom != "CH1_RX_DL_ENABLE_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_fec_type_used_atom != "CH1_RX_FEC_TYPE_USED_NONE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_fec_type_used_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_tx_preloaded_hardware_configs_atom != "CH2_TX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_tx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_rx_preloaded_hardware_configs_atom != "CH2_RX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_rx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch2_lc_postdiv_sel_atom != "CH2_LC_POSTDIV_SEL_SYNTH2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_lc_postdiv_sel_atom_check ( .error(1'b1) );
		end
		if (ch2_sequencer_reg_en_atom != "CH2_SEQUENCER_REG_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_sequencer_reg_en_atom_check ( .error(1'b1) );
		end
		if (ch2_rst_mux_static_sel_atom != "CH2_RST_MUX_STATIC_SEL_HRC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rst_mux_static_sel_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_tx_prbs_pattern_atom != 4'b0000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_tx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_rx_prbs_pattern_atom != 4'b0011)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_rx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_tx_user_clk_only_mode_atom != "CH2_TX_USER_CLK_ONLY_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_tx_user_clk_only_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_tx_width_atom != "CH2_TX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_tx_width_atom_check ( .error(1'b1) );
		end
		if (ch2_xcvr_rx_width_atom != "CH2_RX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_xcvr_rx_width_atom_check ( .error(1'b1) );
		end
		if (ch2_phy_loopback_mode_atom != "CH2_LOOPBACK_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_phy_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_flux_mode_atom != "CH2_FLUX_MODE_FLUX_MODE_BYPASS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_flux_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_sim_mode_atom != "CH2_TX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_sim_mode_atom != "CH2_RX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_dl_enable_atom != "CH2_TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_dl_enable_atom != "CH2_RX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_fec_type_used_atom != "CH2_RX_FEC_TYPE_USED_RS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_fec_type_used_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_tx_preloaded_hardware_configs_atom != "CH3_TX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_tx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_rx_preloaded_hardware_configs_atom != "CH3_RX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_rx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch3_lc_postdiv_sel_atom != "CH3_LC_POSTDIV_SEL_SYNTH2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_lc_postdiv_sel_atom_check ( .error(1'b1) );
		end
		if (ch3_sequencer_reg_en_atom != "CH3_SEQUENCER_REG_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_sequencer_reg_en_atom_check ( .error(1'b1) );
		end
		if (ch3_rst_mux_static_sel_atom != "CH3_RST_MUX_STATIC_SEL_HRC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rst_mux_static_sel_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_tx_prbs_pattern_atom != 4'b0000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_tx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_rx_prbs_pattern_atom != 4'b0111)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_rx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_tx_user_clk_only_mode_atom != "CH3_TX_USER_CLK_ONLY_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_tx_user_clk_only_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_tx_width_atom != "CH3_TX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_tx_width_atom_check ( .error(1'b1) );
		end
		if (ch3_xcvr_rx_width_atom != "CH3_RX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_xcvr_rx_width_atom_check ( .error(1'b1) );
		end
		if (ch3_phy_loopback_mode_atom != "CH3_LOOPBACK_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_phy_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_flux_mode_atom != "CH3_FLUX_MODE_FLUX_MODE_BYPASS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_flux_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_sim_mode_atom != "CH3_TX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_sim_mode_atom != "CH3_RX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_dl_enable_atom != "CH3_TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_dl_enable_atom != "CH3_RX_DL_ENABLE_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_fec_type_used_atom != "CH3_RX_FEC_TYPE_USED_RS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_fec_type_used_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_pll_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_pll_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch0_cdr_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_cdr_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_pll_refclk_select_atom != "CH0_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_pll_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch0_cdr_refclk_select_atom != "CH0_CDR_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_cdr_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_pll_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_pll_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch1_cdr_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_cdr_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_pll_refclk_select_atom != "CH1_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_pll_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch1_cdr_refclk_select_atom != "CH1_CDR_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_cdr_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_pll_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_pll_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch2_cdr_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_cdr_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_pll_refclk_select_atom != "CH2_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_pll_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch2_cdr_refclk_select_atom != "CH2_CDR_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_cdr_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_pll_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_pll_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch3_cdr_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_cdr_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_pll_refclk_select_atom != "CH3_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_pll_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch3_cdr_refclk_select_atom != "CH3_CDR_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_cdr_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_dl_rx_lat_bit_for_async_atom != 18'b010100000100010011)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_dl_rx_lat_bit_for_async_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_dl_rxbit_cntr_pma_atom != "CH0_RX_DL_RXBIT_CNTR_PMA_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_dl_rxbit_cntr_pma_atom_check ( .error(1'b1) );
		end
		if (ch0_rx_dl_rxbit_rollover_atom != 18'b111110100100001111)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_rx_dl_rxbit_rollover_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_dl_rx_lat_bit_for_async_atom != 18'b111110100110100101)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_dl_rx_lat_bit_for_async_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_dl_rxbit_cntr_pma_atom != "CH1_RX_DL_RXBIT_CNTR_PMA_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_dl_rxbit_cntr_pma_atom_check ( .error(1'b1) );
		end
		if (ch1_rx_dl_rxbit_rollover_atom != 18'b001001111001000101)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_rx_dl_rxbit_rollover_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_dl_rx_lat_bit_for_async_atom != 18'b111010100000111101)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_dl_rx_lat_bit_for_async_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_dl_rxbit_cntr_pma_atom != "CH2_RX_DL_RXBIT_CNTR_PMA_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_dl_rxbit_cntr_pma_atom_check ( .error(1'b1) );
		end
		if (ch2_rx_dl_rxbit_rollover_atom != 18'b111000111110011110)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_rx_dl_rxbit_rollover_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_dl_rx_lat_bit_for_async_atom != 18'b100000100111100001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_dl_rx_lat_bit_for_async_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_dl_rxbit_cntr_pma_atom != "CH3_RX_DL_RXBIT_CNTR_PMA_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_dl_rxbit_cntr_pma_atom_check ( .error(1'b1) );
		end
		if (ch3_rx_dl_rxbit_rollover_atom != 18'b001101111001101011)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_rx_dl_rxbit_rollover_atom_check ( .error(1'b1) );
		end
		if (ch0_tx_bond_size_atom != "CH0_TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch0_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch1_tx_bond_size_atom != "CH1_TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch1_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch2_tx_bond_size_atom != "CH2_TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch2_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch3_tx_bond_size_atom != "CH3_TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch3_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (pcie_parity_bypass != "true")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pcie_parity_bypass_check ( .error(1'b1) );
		end
		if (rxbuf_limit_bypass != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					rxbuf_limit_bypass_check ( .error(1'b1) );
		end
		if (maxpayload_size != "MAXPAYLOAD_SIZE_MAX_PAYLOAD_512")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					maxpayload_size_check ( .error(1'b1) );
		end
		if (pldclk_rate != "PLDCLK_RATE_FAST")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pldclk_rate_check ( .error(1'b1) );
		end
		if (port_type != "PORT_TYPE_NATIVE_EP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					port_type_check ( .error(1'b1) );
		end
		if (sris_enable != "SRIS_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sris_enable_check ( .error(1'b1) );
		end
		if (sris_mode != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sris_mode_check ( .error(1'b1) );
		end
		if (sim_mode != "SIM_MODE_DISABLE_VSIM_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sim_mode_check ( .error(1'b1) );
		end
		if (sup_mode != "SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sup_mode_check ( .error(1'b1) );
		end
		if (cvp_enable != "CVP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					cvp_enable_check ( .error(1'b1) );
		end
		if (cii_monitor_en != "CII_MONITOR_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					cii_monitor_en_check ( .error(1'b1) );
		end
		if (pclk_clk_hz != 32'b00111011100110101100101000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pclk_clk_hz_check ( .error(1'b1) );
		end
		if (pf0_cap_link_surprise_down_err_cap != "PF0_CAP_LINK_SURPRISE_DOWN_ERR_CAP_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_cap_link_surprise_down_err_cap_check ( .error(1'b1) );
		end
		if (sys_clk_hz != 32'b00010100110111001001001110000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sys_clk_hz_check ( .error(1'b1) );
		end
		if (link_rate != "LINK_RATE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					link_rate_check ( .error(1'b1) );
		end
		if (link_width != "LINK_WIDTH_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					link_width_check ( .error(1'b1) );
		end
		if (num_of_lanes != "NUM_OF_LANES_NUM_4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					num_of_lanes_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset0 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset0_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset1 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset1_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset2 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset2_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset3 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset3_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset4 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset4_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset5 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset5_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset6 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset6_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset7 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset7_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset8 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset8_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset9 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset9_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset10 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset10_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset11 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset11_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset12 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset12_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset13 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset13_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset14 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset14_check ( .error(1'b1) );
		end
		if (pf0_dsp_16g_tx_preset15 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_16g_tx_preset15_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset0 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset0_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset1 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset1_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset2 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset2_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset3 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset3_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset4 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset4_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset5 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset5_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset6 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset6_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset7 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset7_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset8 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset8_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset9 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset9_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset10 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset10_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset11 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset11_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset12 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset12_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset13 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset13_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset14 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset14_check ( .error(1'b1) );
		end
		if (pf0_dsp_tx_preset15 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_dsp_tx_preset15_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset0 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset0_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset1 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset1_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset2 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset2_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset3 != 7)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset3_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset4 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset4_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset5 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset5_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset6 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset6_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset7 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset7_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset8 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset8_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset9 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset9_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset10 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset10_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset11 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset11_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset12 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset12_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset13 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset13_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset14 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset14_check ( .error(1'b1) );
		end
		if (pf0_usp_16g_tx_preset15 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_16g_tx_preset15_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset0 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset0_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset1 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset1_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset2 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset2_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset3 != 9)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset3_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset4 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset4_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset5 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset5_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset6 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset6_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset7 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset7_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset8 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset8_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset9 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset9_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset10 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset10_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset11 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset11_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset12 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset12_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset13 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset13_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset14 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset14_check ( .error(1'b1) );
		end
		if (pf0_usp_tx_preset15 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_usp_tx_preset15_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar0_enabled != "PF0_PCI_TYPE0_BAR0_ENABLED_ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar0_mask_31_1 != 32'b00000000000000000111111111111111)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar0_mask_31_1_check ( .error(1'b1) );
		end
		if (pf0_bar0_prefetch != "true")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf0_bar0_type != "PF0_BAR0_TYPE_BAR_MEM64")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar0_type_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar1_enabled != "PF0_PCI_TYPE0_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar1_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar1_mask_31_0_check ( .error(1'b1) );
		end
		if (pf0_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar2_enabled != "PF0_PCI_TYPE0_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar2_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar2_mask_31_1_check ( .error(1'b1) );
		end
		if (pf0_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf0_bar2_type != "PF0_BAR2_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar2_type_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar3_enabled != "PF0_PCI_TYPE0_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar3_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar3_mask_31_0_check ( .error(1'b1) );
		end
		if (pf0_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar4_enabled != "PF0_PCI_TYPE0_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar4_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar4_mask_31_1_check ( .error(1'b1) );
		end
		if (pf0_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf0_bar4_type != "PF0_BAR4_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar4_type_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar5_enabled != "PF0_PCI_TYPE0_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_bar5_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_bar5_mask_31_0_check ( .error(1'b1) );
		end
		if (pf0_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf0_rom_bar_enable != "PF0_ROM_BAR_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_rom_bar_enable_check ( .error(1'b1) );
		end
		if (pf0_rom_mask != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_rom_mask_check ( .error(1'b1) );
		end
		if (pf0_rom_bar_enabled != "PF0_ROM_BAR_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_rom_bar_enabled_check ( .error(1'b1) );
		end
		if (pf0_rp_rom_bar_enabled != "PF0_RP_ROM_BAR_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_rp_rom_bar_enabled_check ( .error(1'b1) );
		end
		if (pf0_rp_rom_mask != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_rp_rom_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar0_enabled != "PF0_SRIOV_VF_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar0_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar0_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar0_type != "PF0_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar0_type_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar1_enabled != "PF0_SRIOV_VF_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar1_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar1_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar2_enabled != "PF0_SRIOV_VF_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar2_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar2_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar2_type != "PF0_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar2_type_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar3_enabled != "PF0_SRIOV_VF_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar3_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar3_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar4_enabled != "PF0_SRIOV_VF_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar4_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar4_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar4_type != "PF0_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar4_type_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar5_enabled != "PF0_SRIOV_VF_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar5_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar5_mask_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar0_enabled != "PF1_PCI_TYPE0_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar0_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar0_mask_31_1_check ( .error(1'b1) );
		end
		if (pf1_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf1_bar0_type != "PF1_BAR0_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar0_type_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar1_enabled != "PF1_PCI_TYPE0_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar1_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar1_mask_31_0_check ( .error(1'b1) );
		end
		if (pf1_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar2_enabled != "PF1_PCI_TYPE0_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar2_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar2_mask_31_1_check ( .error(1'b1) );
		end
		if (pf1_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf1_bar2_type != "PF1_BAR2_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar2_type_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar3_enabled != "PF1_PCI_TYPE0_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar3_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar3_mask_31_0_check ( .error(1'b1) );
		end
		if (pf1_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar4_enabled != "PF1_PCI_TYPE0_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar4_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar4_mask_31_1_check ( .error(1'b1) );
		end
		if (pf1_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf1_bar4_type != "PF1_BAR4_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar4_type_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar5_enabled != "PF1_PCI_TYPE0_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_bar5_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_bar5_mask_31_0_check ( .error(1'b1) );
		end
		if (pf1_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf1_rom_bar_enable != "PF1_ROM_BAR_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_rom_bar_enable_check ( .error(1'b1) );
		end
		if (pf1_rom_mask != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_rom_mask_check ( .error(1'b1) );
		end
		if (pf1_rom_bar_enabled != "PF1_ROM_BAR_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_rom_bar_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar0_enabled != "PF1_SRIOV_VF_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar0_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar0_mask_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar0_type != "PF1_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar0_type_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar1_enabled != "PF1_SRIOV_VF_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar1_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar1_mask_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar2_enabled != "PF1_SRIOV_VF_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar2_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar2_mask_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar2_type != "PF1_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar2_type_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar3_enabled != "PF1_SRIOV_VF_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar3_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar3_mask_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar4_enabled != "PF1_SRIOV_VF_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar4_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar4_mask_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar4_type != "PF1_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar4_type_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar5_enabled != "PF1_SRIOV_VF_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar5_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar5_mask_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar0_enabled != "PF2_PCI_TYPE0_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar0_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar0_mask_31_1_check ( .error(1'b1) );
		end
		if (pf2_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf2_bar0_type != "PF2_BAR0_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar0_type_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar1_enabled != "PF2_PCI_TYPE0_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar1_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar1_mask_31_0_check ( .error(1'b1) );
		end
		if (pf2_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar2_enabled != "PF2_PCI_TYPE0_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar2_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar2_mask_31_1_check ( .error(1'b1) );
		end
		if (pf2_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf2_bar2_type != "PF2_BAR2_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar2_type_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar3_enabled != "PF2_PCI_TYPE0_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar3_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar3_mask_31_0_check ( .error(1'b1) );
		end
		if (pf2_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar4_enabled != "PF2_PCI_TYPE0_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar4_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar4_mask_31_1_check ( .error(1'b1) );
		end
		if (pf2_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf2_bar4_type != "PF2_BAR4_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar4_type_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar5_enabled != "PF2_PCI_TYPE0_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_bar5_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_bar5_mask_31_0_check ( .error(1'b1) );
		end
		if (pf2_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf2_rom_bar_enable != "PF2_ROM_BAR_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_rom_bar_enable_check ( .error(1'b1) );
		end
		if (pf2_rom_mask != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_rom_mask_check ( .error(1'b1) );
		end
		if (pf2_rom_bar_enabled != "PF2_ROM_BAR_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_rom_bar_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar0_enabled != "PF2_SRIOV_VF_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar0_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar0_mask_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar0_type != "PF2_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar0_type_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar1_enabled != "PF2_SRIOV_VF_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar1_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar1_mask_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar2_enabled != "PF2_SRIOV_VF_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar2_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar2_mask_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar2_type != "PF2_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar2_type_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar3_enabled != "PF2_SRIOV_VF_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar3_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar3_mask_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar4_enabled != "PF2_SRIOV_VF_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar4_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar4_mask_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar4_type != "PF2_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar4_type_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar5_enabled != "PF2_SRIOV_VF_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar5_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar5_mask_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar0_enabled != "PF3_PCI_TYPE0_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar0_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar0_mask_31_1_check ( .error(1'b1) );
		end
		if (pf3_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf3_bar0_type != "PF3_BAR0_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar0_type_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar1_enabled != "PF3_PCI_TYPE0_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar1_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar1_mask_31_0_check ( .error(1'b1) );
		end
		if (pf3_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar2_enabled != "PF3_PCI_TYPE0_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar2_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar2_mask_31_1_check ( .error(1'b1) );
		end
		if (pf3_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf3_bar2_type != "PF3_BAR2_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar2_type_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar3_enabled != "PF3_PCI_TYPE0_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar3_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar3_mask_31_0_check ( .error(1'b1) );
		end
		if (pf3_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar4_enabled != "PF3_PCI_TYPE0_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar4_mask_31_1 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar4_mask_31_1_check ( .error(1'b1) );
		end
		if (pf3_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf3_bar4_type != "PF3_BAR4_TYPE_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar4_type_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar5_enabled != "PF3_PCI_TYPE0_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_bar5_mask_31_0 != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_bar5_mask_31_0_check ( .error(1'b1) );
		end
		if (pf3_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf3_rom_bar_enable != "PF3_ROM_BAR_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_rom_bar_enable_check ( .error(1'b1) );
		end
		if (pf3_rom_mask != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_rom_mask_check ( .error(1'b1) );
		end
		if (pf3_rom_bar_enabled != "PF3_ROM_BAR_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_rom_bar_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar0_enabled != "PF3_SRIOV_VF_BAR0_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar0_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar0_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar0_mask_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar0_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar0_prefetch_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar0_type != "PF3_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar0_type_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar1_enabled != "PF3_SRIOV_VF_BAR1_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar1_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar1_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar1_mask_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar1_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar1_prefetch_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar2_enabled != "PF3_SRIOV_VF_BAR2_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar2_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar2_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar2_mask_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar2_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar2_prefetch_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar2_type != "PF3_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar2_type_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar3_enabled != "PF3_SRIOV_VF_BAR3_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar3_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar3_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar3_mask_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar3_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar3_prefetch_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar4_enabled != "PF3_SRIOV_VF_BAR4_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar4_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar4_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar4_mask_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar4_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar4_prefetch_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar4_type != "PF3_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar4_type_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar5_enabled != "PF3_SRIOV_VF_BAR5_ENABLED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar5_enabled_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar5_mask != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar5_mask_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_bar5_prefetch != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_bar5_prefetch_check ( .error(1'b1) );
		end
		if (pf1_enable != "PF1_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_enable_check ( .error(1'b1) );
		end
		if (pf2_enable != "PF2_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_enable_check ( .error(1'b1) );
		end
		if (pf3_enable != "PF3_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_enable_check ( .error(1'b1) );
		end
		if (pf0_sriov_enable != "PF0_SRIOV_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_enable_check ( .error(1'b1) );
		end
		if (pf1_sriov_enable != "PF1_SRIOV_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_enable_check ( .error(1'b1) );
		end
		if (pf2_sriov_enable != "PF2_SRIOV_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_enable_check ( .error(1'b1) );
		end
		if (pf3_sriov_enable != "PF3_SRIOV_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_enable_check ( .error(1'b1) );
		end
		if (pf0_sriov_cap_sup_page_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_cap_sup_page_size_check ( .error(1'b1) );
		end
		if (pf1_sriov_cap_sup_page_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_cap_sup_page_size_check ( .error(1'b1) );
		end
		if (pf2_sriov_cap_sup_page_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_cap_sup_page_size_check ( .error(1'b1) );
		end
		if (pf3_sriov_cap_sup_page_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_cap_sup_page_size_check ( .error(1'b1) );
		end
		if (pf0_sriov_num_vf != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_num_vf_check ( .error(1'b1) );
		end
		if (pf1_sriov_num_vf != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_num_vf_check ( .error(1'b1) );
		end
		if (pf2_sriov_num_vf != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_num_vf_check ( .error(1'b1) );
		end
		if (pf3_sriov_num_vf != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_num_vf_check ( .error(1'b1) );
		end
		if (pf0_msi_enable != "PF0_MSI_ENABLE_ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_msi_enable_check ( .error(1'b1) );
		end
		if (pf0_pci_msi_ext_data_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msi_ext_data_cap_check ( .error(1'b1) );
		end
		if (pf0_pci_msi_ext_data_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msi_ext_data_en_check ( .error(1'b1) );
		end
		if (pf0_pci_msi_64_bit_addr_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msi_64_bit_addr_cap_check ( .error(1'b1) );
		end
		if (pf0_pci_msi_multiple_msg_cap != "PF0_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msi_multiple_msg_cap_check ( .error(1'b1) );
		end
		if (pf0_msix_enable != "PF0_MSIX_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_msix_enable_check ( .error(1'b1) );
		end
		if (pf0_pci_msix_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msix_table_size_check ( .error(1'b1) );
		end
		if (pf0_pci_msix_table_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msix_table_offset_check ( .error(1'b1) );
		end
		if (pf0_pci_msix_bir != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msix_bir_check ( .error(1'b1) );
		end
		if (pf0_pci_msix_pba != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msix_pba_check ( .error(1'b1) );
		end
		if (pf0_pci_msix_pba_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msix_pba_offset_check ( .error(1'b1) );
		end
		if (pf0_pci_msix_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_msix_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf0_exvf_msix_cap_enable != "PF0_EXVF_MSIX_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_exvf_msix_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_msix_tablesize_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msix_tablesize_pf0_check ( .error(1'b1) );
		end
		if (exvf_msixtable_offset_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_offset_pf0_check ( .error(1'b1) );
		end
		if (exvf_msixtable_bir_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_bir_pf0_check ( .error(1'b1) );
		end
		if (exvf_msixpba_offset_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_offset_pf0_check ( .error(1'b1) );
		end
		if (exvf_msixpba_bir_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_bir_pf0_check ( .error(1'b1) );
		end
		if (pf1_msi_enable != "PF1_MSI_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_msi_enable_check ( .error(1'b1) );
		end
		if (pf1_pci_msi_ext_data_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msi_ext_data_cap_check ( .error(1'b1) );
		end
		if (pf1_pci_msi_ext_data_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msi_ext_data_en_check ( .error(1'b1) );
		end
		if (pf1_pci_msi_64_bit_addr_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msi_64_bit_addr_cap_check ( .error(1'b1) );
		end
		if (pf1_pci_msi_multiple_msg_cap != "PF1_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msi_multiple_msg_cap_check ( .error(1'b1) );
		end
		if (pf1_msix_enable != "PF1_MSIX_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_msix_enable_check ( .error(1'b1) );
		end
		if (pf1_pci_msix_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msix_table_size_check ( .error(1'b1) );
		end
		if (pf1_pci_msix_table_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msix_table_offset_check ( .error(1'b1) );
		end
		if (pf1_pci_msix_bir != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msix_bir_check ( .error(1'b1) );
		end
		if (pf1_pci_msix_pba != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msix_pba_check ( .error(1'b1) );
		end
		if (pf1_pci_msix_pba_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msix_pba_offset_check ( .error(1'b1) );
		end
		if (pf1_pci_msix_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_msix_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf1_exvf_msix_cap_enable != "PF1_EXVF_MSIX_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_exvf_msix_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_msix_tablesize_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msix_tablesize_pf1_check ( .error(1'b1) );
		end
		if (exvf_msixtable_offset_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_offset_pf1_check ( .error(1'b1) );
		end
		if (exvf_msixtable_bir_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_bir_pf1_check ( .error(1'b1) );
		end
		if (exvf_msixpba_offset_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_offset_pf1_check ( .error(1'b1) );
		end
		if (exvf_msixpba_bir_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_bir_pf1_check ( .error(1'b1) );
		end
		if (pf2_msi_enable != "PF2_MSI_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_msi_enable_check ( .error(1'b1) );
		end
		if (pf2_pci_msi_ext_data_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msi_ext_data_cap_check ( .error(1'b1) );
		end
		if (pf2_pci_msi_ext_data_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msi_ext_data_en_check ( .error(1'b1) );
		end
		if (pf2_pci_msi_64_bit_addr_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msi_64_bit_addr_cap_check ( .error(1'b1) );
		end
		if (pf2_pci_msi_multiple_msg_cap != "PF2_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msi_multiple_msg_cap_check ( .error(1'b1) );
		end
		if (pf2_msix_enable != "PF2_MSIX_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_msix_enable_check ( .error(1'b1) );
		end
		if (pf2_pci_msix_bir != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msix_bir_check ( .error(1'b1) );
		end
		if (pf2_pci_msix_pba != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msix_pba_check ( .error(1'b1) );
		end
		if (pf2_pci_msix_pba_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msix_pba_offset_check ( .error(1'b1) );
		end
		if (pf2_pci_msix_table_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msix_table_offset_check ( .error(1'b1) );
		end
		if (pf2_pci_msix_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msix_table_size_check ( .error(1'b1) );
		end
		if (pf2_pci_msix_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_msix_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf2_exvf_msix_cap_enable != "PF2_EXVF_MSIX_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_exvf_msix_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_msix_tablesize_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msix_tablesize_pf2_check ( .error(1'b1) );
		end
		if (exvf_msixtable_offset_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_offset_pf2_check ( .error(1'b1) );
		end
		if (exvf_msixtable_bir_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_bir_pf2_check ( .error(1'b1) );
		end
		if (exvf_msixpba_offset_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_offset_pf2_check ( .error(1'b1) );
		end
		if (exvf_msixpba_bir_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_bir_pf2_check ( .error(1'b1) );
		end
		if (pf3_msi_enable != "PF3_MSI_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_msi_enable_check ( .error(1'b1) );
		end
		if (pf3_pci_msi_ext_data_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msi_ext_data_cap_check ( .error(1'b1) );
		end
		if (pf3_pci_msi_ext_data_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msi_ext_data_en_check ( .error(1'b1) );
		end
		if (pf3_pci_msi_64_bit_addr_cap != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msi_64_bit_addr_cap_check ( .error(1'b1) );
		end
		if (pf3_pci_msi_multiple_msg_cap != "PF3_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msi_multiple_msg_cap_check ( .error(1'b1) );
		end
		if (pf3_msix_enable != "PF3_MSIX_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_msix_enable_check ( .error(1'b1) );
		end
		if (pf3_pci_msix_bir != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msix_bir_check ( .error(1'b1) );
		end
		if (pf3_pci_msix_pba != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msix_pba_check ( .error(1'b1) );
		end
		if (pf3_pci_msix_pba_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msix_pba_offset_check ( .error(1'b1) );
		end
		if (pf3_pci_msix_table_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msix_table_offset_check ( .error(1'b1) );
		end
		if (pf3_pci_msix_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msix_table_size_check ( .error(1'b1) );
		end
		if (pf3_pci_msix_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_msix_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf3_exvf_msix_cap_enable != "PF3_EXVF_MSIX_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_exvf_msix_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_msix_tablesize_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msix_tablesize_pf3_check ( .error(1'b1) );
		end
		if (exvf_msixtable_offset_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_offset_pf3_check ( .error(1'b1) );
		end
		if (exvf_msixtable_bir_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixtable_bir_pf3_check ( .error(1'b1) );
		end
		if (exvf_msixpba_offset_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_offset_pf3_check ( .error(1'b1) );
		end
		if (exvf_msixpba_bir_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_msixpba_bir_pf3_check ( .error(1'b1) );
		end
		if (pf0_prs_ext_cap_enable != "PF0_PRS_EXT_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_prs_ext_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_prs_ext_cap_outstanding_capacity != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_prs_ext_cap_outstanding_capacity_check ( .error(1'b1) );
		end
		if (pf1_prs_ext_cap_enable != "PF1_PRS_EXT_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_prs_ext_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_prs_ext_cap_outstanding_capacity != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_prs_ext_cap_outstanding_capacity_check ( .error(1'b1) );
		end
		if (pf2_prs_ext_cap_enable != "PF2_PRS_EXT_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_prs_ext_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_prs_ext_cap_outstanding_capacity != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_prs_ext_cap_outstanding_capacity_check ( .error(1'b1) );
		end
		if (pf3_prs_ext_cap_enable != "PF3_PRS_EXT_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_prs_ext_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_prs_ext_cap_outstanding_capacity != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_prs_ext_cap_outstanding_capacity_check ( .error(1'b1) );
		end
		if (pf0_pasid_cap_enable != "PF0_PASID_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pasid_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_pasid_cap_execute_permission_supported != "PF0_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pasid_cap_execute_permission_supported_check ( .error(1'b1) );
		end
		if (pf0_pasid_cap_max_pasid_width != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pasid_cap_max_pasid_width_check ( .error(1'b1) );
		end
		if (pf0_pasid_cap_privileged_mode_supported != "PF0_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pasid_cap_privileged_mode_supported_check ( .error(1'b1) );
		end
		if (pf1_pasid_cap_enable != "PF1_PASID_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pasid_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_pasid_cap_execute_permission_supported != "PF1_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pasid_cap_execute_permission_supported_check ( .error(1'b1) );
		end
		if (pf1_pasid_cap_max_pasid_width != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pasid_cap_max_pasid_width_check ( .error(1'b1) );
		end
		if (pf1_pasid_cap_privileged_mode_supported != "PF1_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pasid_cap_privileged_mode_supported_check ( .error(1'b1) );
		end
		if (pf2_pasid_cap_enable != "PF2_PASID_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pasid_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_pasid_cap_execute_permission_supported != "PF2_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pasid_cap_execute_permission_supported_check ( .error(1'b1) );
		end
		if (pf2_pasid_cap_max_pasid_width != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pasid_cap_max_pasid_width_check ( .error(1'b1) );
		end
		if (pf2_pasid_cap_privileged_mode_supported != "PF2_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pasid_cap_privileged_mode_supported_check ( .error(1'b1) );
		end
		if (pf3_pasid_cap_enable != "PF3_PASID_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pasid_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_pasid_cap_execute_permission_supported != "PF3_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pasid_cap_execute_permission_supported_check ( .error(1'b1) );
		end
		if (pf3_pasid_cap_max_pasid_width != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pasid_cap_max_pasid_width_check ( .error(1'b1) );
		end
		if (pf3_pasid_cap_privileged_mode_supported != "PF3_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pasid_cap_privileged_mode_supported_check ( .error(1'b1) );
		end
		if (pf0_sn_cap_enable != "PF0_SN_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sn_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_sn_ser_num_reg_1_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sn_ser_num_reg_1_dw_check ( .error(1'b1) );
		end
		if (pf0_sn_ser_num_reg_2_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sn_ser_num_reg_2_dw_check ( .error(1'b1) );
		end
		if (pf1_sn_cap_enable != "PF1_SN_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sn_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_sn_ser_num_reg_1_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sn_ser_num_reg_1_dw_check ( .error(1'b1) );
		end
		if (pf1_sn_ser_num_reg_2_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sn_ser_num_reg_2_dw_check ( .error(1'b1) );
		end
		if (pf2_sn_cap_enable != "PF2_SN_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sn_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_sn_ser_num_reg_1_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sn_ser_num_reg_1_dw_check ( .error(1'b1) );
		end
		if (pf2_sn_ser_num_reg_2_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sn_ser_num_reg_2_dw_check ( .error(1'b1) );
		end
		if (pf3_sn_cap_enable != "PF3_SN_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sn_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_sn_ser_num_reg_1_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sn_ser_num_reg_1_dw_check ( .error(1'b1) );
		end
		if (pf3_sn_ser_num_reg_2_dw != 32'b00000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sn_ser_num_reg_2_dw_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_ep_l0s_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_ep_l0s_accpt_latency_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_ep_l1_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_ep_l1_accpt_latency_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_l0s_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_l0s_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_l1_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_l1_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_ep_l0s_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_ep_l0s_accpt_latency_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_ep_l1_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_ep_l1_accpt_latency_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_l0s_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_l0s_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_l1_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_l1_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_ep_l0s_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_ep_l0s_accpt_latency_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_ep_l1_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_ep_l1_accpt_latency_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_l0s_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_l0s_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_l1_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_l1_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_ep_l0s_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_ep_l0s_accpt_latency_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_ep_l1_accpt_latency != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_ep_l1_accpt_latency_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_l0s_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_l0s_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_l1_exit_latency_commclk_dis != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_l1_exit_latency_commclk_dis_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_flr_cap != "PF0_PCIE_CAP_FLR_CAP_NOT_CAPABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_flr_cap_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_flr_cap != "PF1_PCIE_CAP_FLR_CAP_NOT_CAPABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_flr_cap_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_flr_cap != "PF2_PCIE_CAP_FLR_CAP_NOT_CAPABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_flr_cap_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_flr_cap != "PF3_PCIE_CAP_FLR_CAP_NOT_CAPABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_flr_cap_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_port_num != 1)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_port_num_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_port_num != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_port_num_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_port_num != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_port_num_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_port_num != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_port_num_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_slot_clk_config != "true")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_slot_clk_config_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_slot_clk_config != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_slot_clk_config_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_slot_clk_config != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_slot_clk_config_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_slot_clk_config != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_slot_clk_config_check ( .error(1'b1) );
		end
		if (pf0_ltr_cap_enable != "PF0_LTR_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_ltr_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_pcie_slot_imp != "PF0_PCIE_SLOT_IMP_NOT_IMPLEMENTED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_slot_imp_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_slot_power_limit_scale != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_slot_power_limit_scale_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_slot_power_limit_value != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_slot_power_limit_value_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_phy_slot_num != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_phy_slot_num_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_hot_plug_capable != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_hot_plug_capable_check ( .error(1'b1) );
		end
		if (pf0_pcie_cap_ext_tag_en != "true")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pcie_cap_ext_tag_en_check ( .error(1'b1) );
		end
		if (pf1_pcie_cap_ext_tag_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pcie_cap_ext_tag_en_check ( .error(1'b1) );
		end
		if (pf2_pcie_cap_ext_tag_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pcie_cap_ext_tag_en_check ( .error(1'b1) );
		end
		if (pf3_pcie_cap_ext_tag_en != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pcie_cap_ext_tag_en_check ( .error(1'b1) );
		end
		if (cfg_ptm_auto_update_signal != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					cfg_ptm_auto_update_signal_check ( .error(1'b1) );
		end
		if (ptm_autoupdate != "PTM_AUTOUPDATE_AUTOUPDATE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ptm_autoupdate_check ( .error(1'b1) );
		end
		if (ptm_enable != "PTM_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ptm_enable_check ( .error(1'b1) );
		end
		if (pf0_ats_cap_enable != "PF0_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_exvf_ats_cap_enable != "PF0_EXVF_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_exvf_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_ats_cap_invalidate_q_depth != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_ats_cap_invalidate_q_depth_check ( .error(1'b1) );
		end
		if (pf0_ats_exvf_align_request != "PF0_ATS_EXVF_ALIGN_REQUEST_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_ats_exvf_align_request_check ( .error(1'b1) );
		end
		if (pf1_ats_cap_enable != "PF1_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_exvf_ats_cap_enable != "PF1_EXVF_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_exvf_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_ats_cap_invalidate_q_depth != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_ats_cap_invalidate_q_depth_check ( .error(1'b1) );
		end
		if (pf1_ats_exvf_align_request != "PF1_ATS_EXVF_ALIGN_REQUEST_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_ats_exvf_align_request_check ( .error(1'b1) );
		end
		if (pf2_ats_cap_enable != "PF2_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_exvf_ats_cap_enable != "PF2_EXVF_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_exvf_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_ats_cap_invalidate_q_depth != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_ats_cap_invalidate_q_depth_check ( .error(1'b1) );
		end
		if (pf2_ats_exvf_align_request != "PF2_ATS_EXVF_ALIGN_REQUEST_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_ats_exvf_align_request_check ( .error(1'b1) );
		end
		if (pf3_ats_cap_enable != "PF3_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_exvf_ats_cap_enable != "PF3_EXVF_ATS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_exvf_ats_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_ats_cap_invalidate_q_depth != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_ats_cap_invalidate_q_depth_check ( .error(1'b1) );
		end
		if (pf3_ats_exvf_align_request != "PF3_ATS_EXVF_ALIGN_REQUEST_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_ats_exvf_align_request_check ( .error(1'b1) );
		end
		if (pf0_tph_cap_enable != "PF0_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_int_vec != "PF0_TPH_REQ_CAP_INT_VEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_int_vec_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_int_vec_vfcomm_cs2 != "PF0_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_int_vec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_st_table_loc_0_vfcomm_cs2 != "PF0_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_st_table_loc_0_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_st_table_loc_1 != "PF0_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_st_table_loc_1_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_st_table_loc_1_vfcomm_cs2 != "PF0_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_st_table_loc_1_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_st_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_st_table_size_check ( .error(1'b1) );
		end
		if (pf0_tph_req_cap_st_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_cap_st_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf0_tph_req_device_spec != "PF0_TPH_REQ_DEVICE_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_device_spec_check ( .error(1'b1) );
		end
		if (pf0_tph_req_device_spec_vfcomm_cs2 != "PF0_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_tph_req_device_spec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf0_exvf_tph_cap_enable != "PF0_EXVF_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_exvf_tph_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablelocation_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablelocation_pf0_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablesize_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablesize_pf0_check ( .error(1'b1) );
		end
		if (pf1_tph_cap_enable != "PF1_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_int_vec != "PF1_TPH_REQ_CAP_INT_VEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_int_vec_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_int_vec_vfcomm_cs2 != "PF1_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_int_vec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_st_table_loc_0_vfcomm_cs2 != "PF1_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_st_table_loc_0_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_st_table_loc_1 != "PF1_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_st_table_loc_1_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_st_table_loc_1_vfcomm_cs2 != "PF1_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_st_table_loc_1_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_st_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_st_table_size_check ( .error(1'b1) );
		end
		if (pf1_tph_req_cap_st_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_cap_st_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf1_tph_req_device_spec != "PF1_TPH_REQ_DEVICE_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_device_spec_check ( .error(1'b1) );
		end
		if (pf1_tph_req_device_spec_vfcomm_cs2 != "PF1_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_tph_req_device_spec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf1_exvf_tph_cap_enable != "PF1_EXVF_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_exvf_tph_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablelocation_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablelocation_pf1_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablesize_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablesize_pf1_check ( .error(1'b1) );
		end
		if (pf2_tph_cap_enable != "PF2_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_int_vec != "PF2_TPH_REQ_CAP_INT_VEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_int_vec_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_int_vec_vfcomm_cs2 != "PF2_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_int_vec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_st_table_loc_0_vfcomm_cs2 != "PF2_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_st_table_loc_0_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_st_table_loc_1 != "PF2_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_st_table_loc_1_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_st_table_loc_1_vfcomm_cs2 != "PF2_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_st_table_loc_1_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_st_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_st_table_size_check ( .error(1'b1) );
		end
		if (pf2_tph_req_cap_st_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_cap_st_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf2_tph_req_device_spec != "PF2_TPH_REQ_DEVICE_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_device_spec_check ( .error(1'b1) );
		end
		if (pf2_tph_req_device_spec_vfcomm_cs2 != "PF2_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_tph_req_device_spec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf2_exvf_tph_cap_enable != "PF2_EXVF_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_exvf_tph_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablelocation_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablelocation_pf2_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablesize_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablesize_pf2_check ( .error(1'b1) );
		end
		if (pf3_tph_cap_enable != "PF3_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_int_vec != "PF3_TPH_REQ_CAP_INT_VEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_int_vec_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_int_vec_vfcomm_cs2 != "PF3_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_int_vec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_st_table_loc_0_vfcomm_cs2 != "PF3_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_st_table_loc_0_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_st_table_loc_1 != "PF3_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_st_table_loc_1_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_st_table_loc_1_vfcomm_cs2 != "PF3_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_st_table_loc_1_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_st_table_size != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_st_table_size_check ( .error(1'b1) );
		end
		if (pf3_tph_req_cap_st_table_size_vfcomm_cs2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_cap_st_table_size_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf3_tph_req_device_spec != "PF3_TPH_REQ_DEVICE_SPEC_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_device_spec_check ( .error(1'b1) );
		end
		if (pf3_tph_req_device_spec_vfcomm_cs2 != "PF3_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_tph_req_device_spec_vfcomm_cs2_check ( .error(1'b1) );
		end
		if (pf3_exvf_tph_cap_enable != "PF3_EXVF_TPH_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_exvf_tph_cap_enable_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablelocation_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablelocation_pf3_check ( .error(1'b1) );
		end
		if (exvf_tph_sttablesize_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_tph_sttablesize_pf3_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_enable != "PF0_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_exvf_acs_cap_enable != "PF0_EXVF_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_exvf_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_src_valid != "PF0_ACS_CAP_ACS_SRC_VALID_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_src_valid_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_at_block != "PF0_ACS_CAP_ACS_AT_BLOCK_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_at_block_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_p2p_req_redirect != "PF0_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_p2p_req_redirect_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_p2p_cpl_redirect != "PF0_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_p2p_cpl_redirect_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_usp_forwarding != "PF0_ACS_CAP_ACS_USP_FORWARDING_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_usp_forwarding_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_p2p_egress_control != "PF0_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_p2p_egress_control_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_egress_ctrl_size != 8)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_egress_ctrl_size_check ( .error(1'b1) );
		end
		if (pf0_acs_cap_acs_direct_translated_p2p != "PF0_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_acs_cap_acs_direct_translated_p2p_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_enable != "PF1_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_exvf_acs_cap_enable != "PF1_EXVF_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_exvf_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_src_valid != "PF1_ACS_CAP_ACS_SRC_VALID_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_src_valid_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_at_block != "PF1_ACS_CAP_ACS_AT_BLOCK_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_at_block_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_p2p_req_redirect != "PF1_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_p2p_req_redirect_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_p2p_cpl_redirect != "PF1_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_p2p_cpl_redirect_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_usp_forwarding != "PF1_ACS_CAP_ACS_USP_FORWARDING_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_usp_forwarding_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_p2p_egress_control != "PF1_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_p2p_egress_control_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_egress_ctrl_size != 8)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_egress_ctrl_size_check ( .error(1'b1) );
		end
		if (pf1_acs_cap_acs_direct_translated_p2p != "PF1_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_acs_cap_acs_direct_translated_p2p_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_enable != "PF2_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_exvf_acs_cap_enable != "PF2_EXVF_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_exvf_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_src_valid != "PF2_ACS_CAP_ACS_SRC_VALID_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_src_valid_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_at_block != "PF2_ACS_CAP_ACS_AT_BLOCK_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_at_block_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_p2p_req_redirect != "PF2_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_p2p_req_redirect_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_p2p_cpl_redirect != "PF2_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_p2p_cpl_redirect_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_usp_forwarding != "PF2_ACS_CAP_ACS_USP_FORWARDING_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_usp_forwarding_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_p2p_egress_control != "PF2_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_p2p_egress_control_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_egress_ctrl_size != 8)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_egress_ctrl_size_check ( .error(1'b1) );
		end
		if (pf2_acs_cap_acs_direct_translated_p2p != "PF2_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_acs_cap_acs_direct_translated_p2p_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_enable != "PF3_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_exvf_acs_cap_enable != "PF3_EXVF_ACS_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_exvf_acs_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_src_valid != "PF3_ACS_CAP_ACS_SRC_VALID_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_src_valid_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_at_block != "PF3_ACS_CAP_ACS_AT_BLOCK_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_at_block_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_p2p_req_redirect != "PF3_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_p2p_req_redirect_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_p2p_cpl_redirect != "PF3_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_p2p_cpl_redirect_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_usp_forwarding != "PF3_ACS_CAP_ACS_USP_FORWARDING_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_usp_forwarding_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_p2p_egress_control != "PF3_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_p2p_egress_control_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_egress_ctrl_size != 8)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_egress_ctrl_size_check ( .error(1'b1) );
		end
		if (pf3_acs_cap_acs_direct_translated_p2p != "PF3_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_acs_cap_acs_direct_translated_p2p_check ( .error(1'b1) );
		end
		if (pf0_virtio_en != "PF0_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_virtio_en_check ( .error(1'b1) );
		end
		if (pf1_virtio_en != "PF1_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_virtio_en_check ( .error(1'b1) );
		end
		if (pf2_virtio_en != "PF2_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_virtio_en_check ( .error(1'b1) );
		end
		if (pf3_virtio_en != "PF3_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_virtio_en_check ( .error(1'b1) );
		end
		if (pf0_exvf_virtio_en != "PF0_EXVF_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_exvf_virtio_en_check ( .error(1'b1) );
		end
		if (pf1_exvf_virtio_en != "PF1_EXVF_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_exvf_virtio_en_check ( .error(1'b1) );
		end
		if (pf2_exvf_virtio_en != "PF2_EXVF_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_exvf_virtio_en_check ( .error(1'b1) );
		end
		if (pf3_exvf_virtio_en != "PF3_EXVF_VIRTIO_EN_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_exvf_virtio_en_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_device_id_check ( .error(1'b1) );
		end
		if (pf0_pci_type0_vendor_id != 4466)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_pci_type0_vendor_id_check ( .error(1'b1) );
		end
		if (pf0_revision_id != 1)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_revision_id_check ( .error(1'b1) );
		end
		if (pf0_base_class_code != 255)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_base_class_code_check ( .error(1'b1) );
		end
		if (pf0_subclass_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_subclass_code_check ( .error(1'b1) );
		end
		if (pf0_program_interface != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_program_interface_check ( .error(1'b1) );
		end
		if (pf0_subsys_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_subsys_vendor_id_check ( .error(1'b1) );
		end
		if (pf0_subsys_dev_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_subsys_dev_id_check ( .error(1'b1) );
		end
		if (pf0_sriov_vf_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_sriov_vf_device_id_check ( .error(1'b1) );
		end
		if (exvf_subsysid_pf0 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_subsysid_pf0_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_vendor_id_check ( .error(1'b1) );
		end
		if (pf1_pci_type0_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_pci_type0_device_id_check ( .error(1'b1) );
		end
		if (pf1_revision_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_revision_id_check ( .error(1'b1) );
		end
		if (pf1_base_class_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_base_class_code_check ( .error(1'b1) );
		end
		if (pf1_subclass_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_subclass_code_check ( .error(1'b1) );
		end
		if (pf1_program_interface != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_program_interface_check ( .error(1'b1) );
		end
		if (pf1_subsys_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_subsys_vendor_id_check ( .error(1'b1) );
		end
		if (pf1_subsys_dev_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_subsys_dev_id_check ( .error(1'b1) );
		end
		if (pf1_sriov_vf_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_sriov_vf_device_id_check ( .error(1'b1) );
		end
		if (exvf_subsysid_pf1 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_subsysid_pf1_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_vendor_id_check ( .error(1'b1) );
		end
		if (pf2_pci_type0_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_pci_type0_device_id_check ( .error(1'b1) );
		end
		if (pf2_revision_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_revision_id_check ( .error(1'b1) );
		end
		if (pf2_base_class_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_base_class_code_check ( .error(1'b1) );
		end
		if (pf2_subclass_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_subclass_code_check ( .error(1'b1) );
		end
		if (pf2_program_interface != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_program_interface_check ( .error(1'b1) );
		end
		if (pf2_subsys_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_subsys_vendor_id_check ( .error(1'b1) );
		end
		if (pf2_subsys_dev_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_subsys_dev_id_check ( .error(1'b1) );
		end
		if (pf2_sriov_vf_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_sriov_vf_device_id_check ( .error(1'b1) );
		end
		if (exvf_subsysid_pf2 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_subsysid_pf2_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_vendor_id_check ( .error(1'b1) );
		end
		if (pf3_pci_type0_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_pci_type0_device_id_check ( .error(1'b1) );
		end
		if (pf3_revision_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_revision_id_check ( .error(1'b1) );
		end
		if (pf3_base_class_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_base_class_code_check ( .error(1'b1) );
		end
		if (pf3_subclass_code != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_subclass_code_check ( .error(1'b1) );
		end
		if (pf3_program_interface != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_program_interface_check ( .error(1'b1) );
		end
		if (pf3_subsys_vendor_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_subsys_vendor_id_check ( .error(1'b1) );
		end
		if (pf3_subsys_dev_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_subsys_dev_id_check ( .error(1'b1) );
		end
		if (pf3_sriov_vf_device_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_sriov_vf_device_id_check ( .error(1'b1) );
		end
		if (exvf_subsysid_pf3 != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					exvf_subsysid_pf3_check ( .error(1'b1) );
		end
		if (vsec_select != "false")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					vsec_select_check ( .error(1'b1) );
		end
		if (pf0_user_vsec_cap_enable != "PF0_USER_VSEC_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_user_vsec_cap_enable_check ( .error(1'b1) );
		end
		if (pf1_user_vsec_cap_enable != "PF1_USER_VSEC_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_user_vsec_cap_enable_check ( .error(1'b1) );
		end
		if (pf2_user_vsec_cap_enable != "PF2_USER_VSEC_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_user_vsec_cap_enable_check ( .error(1'b1) );
		end
		if (pf3_user_vsec_cap_enable != "PF3_USER_VSEC_CAP_ENABLE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_user_vsec_cap_enable_check ( .error(1'b1) );
		end
		if (vsec_next_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					vsec_next_offset_check ( .error(1'b1) );
		end
		if (pf1_user_vsec_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_user_vsec_offset_check ( .error(1'b1) );
		end
		if (pf2_user_vsec_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_user_vsec_offset_check ( .error(1'b1) );
		end
		if (pf3_user_vsec_offset != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_user_vsec_offset_check ( .error(1'b1) );
		end
		if (cvp_vendor_specific_header_id != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					cvp_vendor_specific_header_id_check ( .error(1'b1) );
		end
		if (drop_vendor0_msg != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					drop_vendor0_msg_check ( .error(1'b1) );
		end
		if (drop_vendor1_msg != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					drop_vendor1_msg_check ( .error(1'b1) );
		end
		if (pf0_int_pin != "PF0_INT_PIN_NO_INT")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_int_pin_check ( .error(1'b1) );
		end
		if (pf1_int_pin != "PF1_INT_PIN_NO_INT")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf1_int_pin_check ( .error(1'b1) );
		end
		if (pf2_int_pin != "PF2_INT_PIN_NO_INT")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf2_int_pin_check ( .error(1'b1) );
		end
		if (pf3_int_pin != "PF3_INT_PIN_NO_INT")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf3_int_pin_check ( .error(1'b1) );
		end
		if (dtk_mode_en != "DTK_MODE_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					dtk_mode_en_check ( .error(1'b1) );
		end
		if (hrc_arb_sel != "HRC_ARB_SEL_LOCAL_QUAD_ARB")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					hrc_arb_sel_check ( .error(1'b1) );
		end
		if (num_arb_ip != 1)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					num_arb_ip_check ( .error(1'b1) );
		end
		if (pcie_hrc_pulse_sel != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pcie_hrc_pulse_sel_check ( .error(1'b1) );
		end
		if (pf0_port_logic_fast_link_mode != "PF0_PORT_LOGIC_FAST_LINK_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_port_logic_fast_link_mode_check ( .error(1'b1) );
		end
		if (pf0_prefetch_decode != "PF0_PREFETCH_DECODE_PREF64")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pf0_prefetch_decode_check ( .error(1'b1) );
		end
		if (usb_hrc_pulse_sel != 0)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					usb_hrc_pulse_sel_check ( .error(1'b1) );
		end
		if (pcie_pcs_mode != "PCIE_PCS_MODE_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					pcie_pcs_mode_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_clk_mux_0_sel != "SEL_SAME_QUAD_PCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_clk_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_clk_mux_1_sel != "SEL_SAME_QUAD_PCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_clk_mux_1_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_clk_mux_2_sel != "SEL_SAME_QUAD_PCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_clk_mux_2_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_clk_mux_3_sel != "SEL_SAME_QUAD_PCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_clk_mux_3_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_hps_clkmux_0_sel != "SEL_HPS_PCS1_ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_hps_clkmux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rst_mux_0_sel != "SEL_SAME_QUAD_PCS_RST")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rst_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rst_mux_1_sel != "SEL_SAME_QUAD_PCS_RST")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rst_mux_1_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rst_mux_2_sel != "SEL_SAME_QUAD_PCS_RST")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rst_mux_2_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rst_mux_3_sel != "SEL_SAME_QUAD_PCS_RST")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rst_mux_3_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_tx_mux_0_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_tx_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_tx_mux_1_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_tx_mux_1_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_tx_mux_2_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_tx_mux_2_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_tx_mux_3_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_tx_mux_3_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_hps_demux_0_sel != "SEL_HPS_PCS1_ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_hps_demux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_hps_mux_0_sel != "SEL_HPS_PCS1_ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_hps_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rx_demux_0_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rx_demux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rx_demux_1_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rx_demux_1_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rx_demux_2_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rx_demux_2_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_pcs_rx_demux_3_sel != "SEL_SAME_QUAD_PCIE_CTRL")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_pcs_rx_demux_3_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_clk_mux_0_sel != "SEL_MIDDLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_clk_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pcie_data_mux_0_sel != "SEL_MIDDLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pcie_data_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_dr_enabled != "DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_dr_enabled_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_duplex_mode != "DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_duplex_mode_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_pld_channel_identifier != "PLD_CHANNEL_IDENTIFIER_PHIP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_pld_channel_identifier_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_clkout1_divider != "RX_CLKOUT1_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_clkout1_divider_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_clkout2_divider != "RX_CLKOUT2_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_clkout2_divider_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_en != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_en_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_fifo_mode != "RX_FIFO_MODE_PHASE_COMP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_fifo_mode_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_fifo_width != "RX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_fifo_width_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_fifo_wr_clk_hz != 36'b000000010001111000011010001100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_fifo_wr_clk_hz_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_user1_clk_dynamic_mux != "RX_USER1_CLK_DYNAMIC_MUX_C2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_user1_clk_dynamic_mux_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_rx_user2_clk_dynamic_mux != "RX_USER2_CLK_DYNAMIC_MUX_UX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_rx_user2_clk_dynamic_mux_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_sup_mode != "SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_sup_mode_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_clkout1_divider != "TX_CLKOUT1_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_clkout1_divider_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_clkout2_divider != "TX_CLKOUT2_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_clkout2_divider_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_en != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_en_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_fifo_mode != "TX_FIFO_MODE_PHASE_COMP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_fifo_mode_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_fifo_rd_clk_hz != 36'b000000010001111000011010001100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_fifo_rd_clk_hz_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_fifo_width != "TX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_fifo_width_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_user1_clk_dynamic_mux != "TX_USER1_CLK_DYNAMIC_MUX_C1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_user1_clk_dynamic_mux_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_tx_user2_clk_dynamic_mux != "TX_USER2_CLK_DYNAMIC_MUX_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_tx_user2_clk_dynamic_mux_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_dp_0_vc_rx_pldif_wm_en != "VC_RX_PLDIF_WM_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_dp_0_vc_rx_pldif_wm_en_check ( .error(1'b1) );
		end
		if (sm_pld_rx_mux_0_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_pld_rx_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_pld_tx_demux_0_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_pld_tx_demux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_sel_check ( .error(1'b1) );
		end
		if (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_sel_check ( .error(1'b1) );
		end
	endgenerate

	system_intel_pcie_gts_0_pcie_hal_top_2100_okrywsy #(
		.ch0_pcs_l_tx_en_atom                                ("FALSE"),
		.ch0_pcs_l_rx_en_atom                                ("FALSE"),
		.ch0_fec_loopback_mode_atom                          ("CH0_LOOPBACK_MODE_DISABLE"),
		.ch0_fec_dyn_tx_mux_atom                             ("CH0_DYN_TX_MUX_ETHPCS"),
		.ch0_fec_error_atom                                  ("FALSE"),
		.ch0_fec_rx_en_atom                                  ("TRUE"),
		.ch0_fec_tx_en_atom                                  ("TRUE"),
		.ch0_fec_mode_atom                                   ("CH0_FEC_MODE_RSFEC"),
		.ch1_pcs_l_tx_en_atom                                ("FALSE"),
		.ch1_pcs_l_rx_en_atom                                ("FALSE"),
		.ch1_fec_loopback_mode_atom                          ("CH1_LOOPBACK_MODE_DISABLE"),
		.ch1_fec_dyn_tx_mux_atom                             ("CH1_DYN_TX_MUX_UNUSED"),
		.ch1_fec_error_atom                                  ("FALSE"),
		.ch1_fec_rx_en_atom                                  ("FALSE"),
		.ch1_fec_tx_en_atom                                  ("FALSE"),
		.ch1_fec_mode_atom                                   ("CH1_FEC_MODE_DISABLED"),
		.ch2_pcs_l_tx_en_atom                                ("FALSE"),
		.ch2_pcs_l_rx_en_atom                                ("FALSE"),
		.ch2_fec_loopback_mode_atom                          ("CH2_LOOPBACK_MODE_DISABLE"),
		.ch2_fec_dyn_tx_mux_atom                             ("CH2_DYN_TX_MUX_ETHPCS"),
		.ch2_fec_error_atom                                  ("FALSE"),
		.ch2_fec_rx_en_atom                                  ("TRUE"),
		.ch2_fec_tx_en_atom                                  ("TRUE"),
		.ch2_fec_mode_atom                                   ("CH2_FEC_MODE_RSFEC"),
		.ch3_pcs_l_tx_en_atom                                ("FALSE"),
		.ch3_pcs_l_rx_en_atom                                ("FALSE"),
		.ch3_fec_loopback_mode_atom                          ("CH3_LOOPBACK_MODE_DISABLE"),
		.ch3_fec_dyn_tx_mux_atom                             ("CH3_DYN_TX_MUX_DESKEW"),
		.ch3_fec_error_atom                                  ("FALSE"),
		.ch3_fec_rx_en_atom                                  ("TRUE"),
		.ch3_fec_tx_en_atom                                  ("TRUE"),
		.ch3_fec_mode_atom                                   ("CH3_FEC_MODE_RSFEC"),
		.ch0_xcvr_rx_prbs_monitor_en_atom                    ("CH0_RX_PRBS_MONITOR_EN_DISABLE"),
		.ch1_xcvr_rx_prbs_monitor_en_atom                    ("CH1_RX_PRBS_MONITOR_EN_ENABLE"),
		.ch2_xcvr_rx_prbs_monitor_en_atom                    ("CH2_RX_PRBS_MONITOR_EN_ENABLE"),
		.ch3_xcvr_rx_prbs_monitor_en_atom                    ("CH3_RX_PRBS_MONITOR_EN_ENABLE"),
		.ch0_tx_prbs_gen_en_atom                             ("CH0_TX_PRBS_GEN_EN_DISABLE"),
		.ch1_tx_prbs_gen_en_atom                             ("CH1_TX_PRBS_GEN_EN_DISABLE"),
		.ch2_tx_prbs_gen_en_atom                             ("CH2_TX_PRBS_GEN_EN_DISABLE"),
		.ch3_tx_prbs_gen_en_atom                             ("CH3_TX_PRBS_GEN_EN_DISABLE"),
		.ch0_rx_user1_clk_mux_dynamic_sel_atom               ("CH0_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch0_rx_user2_clk_mux_dynamic_sel_atom               ("CH0_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch0_tx_user1_clk_mux_dynamic_sel_atom               ("CH0_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch0_tx_user2_clk_mux_dynamic_sel_atom               ("CH0_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch1_rx_user1_clk_mux_dynamic_sel_atom               ("CH1_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch1_rx_user2_clk_mux_dynamic_sel_atom               ("CH1_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch1_tx_user1_clk_mux_dynamic_sel_atom               ("CH1_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch1_tx_user2_clk_mux_dynamic_sel_atom               ("CH1_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch2_rx_user1_clk_mux_dynamic_sel_atom               ("CH2_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch2_rx_user2_clk_mux_dynamic_sel_atom               ("CH2_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch2_tx_user1_clk_mux_dynamic_sel_atom               ("CH2_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch2_tx_user2_clk_mux_dynamic_sel_atom               ("CH2_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch3_rx_user1_clk_mux_dynamic_sel_atom               ("CH3_RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch3_rx_user2_clk_mux_dynamic_sel_atom               ("CH3_RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch3_tx_user1_clk_mux_dynamic_sel_atom               ("CH3_TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch3_tx_user2_clk_mux_dynamic_sel_atom               ("CH3_TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch0_pcie_mode_atom                                  ("CH0_PCIE_MODE_GEN4"),
		.ch1_pcie_mode_atom                                  ("CH1_PCIE_MODE_GEN4"),
		.ch2_pcie_mode_atom                                  ("CH2_PCIE_MODE_GEN4"),
		.ch3_pcie_mode_atom                                  ("CH3_PCIE_MODE_GEN4"),
		.ch0_xcvr_rx_protocol_hint_atom                      ("CH0_RX_PROTOCOL_HINT_DISABLED"),
		.ch1_xcvr_rx_protocol_hint_atom                      ("CH1_RX_PROTOCOL_HINT_DISABLED"),
		.ch2_xcvr_rx_protocol_hint_atom                      ("CH2_RX_PROTOCOL_HINT_DISABLED"),
		.ch3_xcvr_rx_protocol_hint_atom                      ("CH3_RX_PROTOCOL_HINT_DISABLED"),
		.ch0_clkrx_refclk_cssm_fw_control_atom               ("CH0_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch1_clkrx_refclk_cssm_fw_control_atom               ("CH1_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch2_clkrx_refclk_cssm_fw_control_atom               ("CH2_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch3_clkrx_refclk_cssm_fw_control_atom               ("CH3_CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch0_clkrx_refclk_sector_specifies_refclk_ready_atom ("CH0_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch1_clkrx_refclk_sector_specifies_refclk_ready_atom ("CH1_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch2_clkrx_refclk_sector_specifies_refclk_ready_atom ("CH2_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch3_clkrx_refclk_sector_specifies_refclk_ready_atom ("CH3_CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch0_local_refclk_cssm_fw_control_atom               ("CH0_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch1_local_refclk_cssm_fw_control_atom               ("CH1_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch2_local_refclk_cssm_fw_control_atom               ("CH2_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch3_local_refclk_cssm_fw_control_atom               ("CH3_LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch0_local_refclk_sector_specifies_refclk_ready_atom ("CH0_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch1_local_refclk_sector_specifies_refclk_ready_atom ("CH1_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch2_local_refclk_sector_specifies_refclk_ready_atom ("CH2_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch3_local_refclk_sector_specifies_refclk_ready_atom ("CH3_LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch0_tx_bonding_category_atom                        ("CH0_TX_BONDING_CATEGORY_BONDING_LEADER"),
		.ch1_tx_bonding_category_atom                        ("CH1_TX_BONDING_CATEGORY_BONDING_FOLLOWER"),
		.ch2_tx_bonding_category_atom                        ("CH2_TX_BONDING_CATEGORY_BONDING_FOLLOWER"),
		.ch3_tx_bonding_category_atom                        ("CH3_TX_BONDING_CATEGORY_BONDING_FOLLOWER"),
		.hal_num_of_lanes_hwtcl                              (4),
		.ch0_duplex_mode_atom                                ("CH0_DUPLEX_MODE_DUPLEX"),
		.ch0_fec_spec_atom                                   ("CH0_FEC_SPEC_DISABLED"),
		.ch0_fracture_atom                                   ("CH0_FRACTURE_UNUSED"),
		.ch0_dr_enabled_atom                                 ("CH0_DR_ENABLED_DR_DISABLED"),
		.ch0_sup_mode_atom                                   ("CH0_SUP_MODE_USER_MODE"),
		.ch0_sim_mode_atom                                   ("CH0_SIM_MODE_DISABLE"),
		.ch1_duplex_mode_atom                                ("CH1_DUPLEX_MODE_DUPLEX"),
		.ch1_fec_spec_atom                                   ("CH1_FEC_SPEC_DISABLED"),
		.ch1_fracture_atom                                   ("CH1_FRACTURE_UNUSED"),
		.ch1_dr_enabled_atom                                 ("CH1_DR_ENABLED_DR_DISABLED"),
		.ch1_sup_mode_atom                                   ("CH1_SUP_MODE_USER_MODE"),
		.ch1_sim_mode_atom                                   ("CH1_SIM_MODE_DISABLE"),
		.ch2_duplex_mode_atom                                ("CH2_DUPLEX_MODE_DUPLEX"),
		.ch2_fec_spec_atom                                   ("CH2_FEC_SPEC_DISABLED"),
		.ch2_fracture_atom                                   ("CH2_FRACTURE_UNUSED"),
		.ch2_dr_enabled_atom                                 ("CH2_DR_ENABLED_DR_DISABLED"),
		.ch2_sup_mode_atom                                   ("CH2_SUP_MODE_USER_MODE"),
		.ch2_sim_mode_atom                                   ("CH2_SIM_MODE_DISABLE"),
		.ch3_duplex_mode_atom                                ("CH3_DUPLEX_MODE_DUPLEX"),
		.ch3_fec_spec_atom                                   ("CH3_FEC_SPEC_DISABLED"),
		.ch3_fracture_atom                                   ("CH3_FRACTURE_UNUSED"),
		.ch3_dr_enabled_atom                                 ("CH3_DR_ENABLED_DR_DISABLED"),
		.ch3_sup_mode_atom                                   ("CH3_SUP_MODE_USER_MODE"),
		.ch3_sim_mode_atom                                   ("CH3_SIM_MODE_DISABLE"),
		.ch0_xcvr_tx_preloaded_hardware_configs_atom         ("CH0_TX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch0_xcvr_rx_preloaded_hardware_configs_atom         ("CH0_RX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch0_lc_postdiv_sel_atom                             ("CH0_LC_POSTDIV_SEL_SYNTH2"),
		.ch0_sequencer_reg_en_atom                           ("CH0_SEQUENCER_REG_EN_ENABLE"),
		.ch0_rst_mux_static_sel_atom                         ("CH0_RST_MUX_STATIC_SEL_HRC"),
		.ch0_xcvr_tx_prbs_pattern_atom                       (4'b0000),
		.ch0_xcvr_rx_prbs_pattern_atom                       (4'b0000),
		.ch0_xcvr_tx_user_clk_only_mode_atom                 ("CH0_TX_USER_CLK_ONLY_MODE_DISABLE"),
		.ch0_xcvr_tx_width_atom                              ("CH0_TX_WIDTH_X16"),
		.ch0_xcvr_rx_width_atom                              ("CH0_RX_WIDTH_X16"),
		.ch0_phy_loopback_mode_atom                          ("CH0_LOOPBACK_MODE_DISABLED"),
		.ch0_flux_mode_atom                                  ("CH0_FLUX_MODE_FLUX_MODE_BYPASS"),
		.ch0_tx_sim_mode_atom                                ("CH0_TX_SIM_MODE_DISABLE"),
		.ch0_rx_sim_mode_atom                                ("CH0_RX_SIM_MODE_DISABLE"),
		.ch0_tx_dl_enable_atom                               ("CH0_TX_DL_ENABLE_DISABLE"),
		.ch0_rx_dl_enable_atom                               ("CH0_RX_DL_ENABLE_ENABLE"),
		.ch0_rx_fec_type_used_atom                           ("CH0_RX_FEC_TYPE_USED_RS"),
		.ch1_xcvr_tx_preloaded_hardware_configs_atom         ("CH1_TX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch1_xcvr_rx_preloaded_hardware_configs_atom         ("CH1_RX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch1_lc_postdiv_sel_atom                             ("CH1_LC_POSTDIV_SEL_SYNTH2"),
		.ch1_sequencer_reg_en_atom                           ("CH1_SEQUENCER_REG_EN_DISABLE"),
		.ch1_rst_mux_static_sel_atom                         ("CH1_RST_MUX_STATIC_SEL_HRC"),
		.ch1_xcvr_tx_prbs_pattern_atom                       (4'b0000),
		.ch1_xcvr_rx_prbs_pattern_atom                       (4'b0001),
		.ch1_xcvr_tx_user_clk_only_mode_atom                 ("CH1_TX_USER_CLK_ONLY_MODE_DISABLE"),
		.ch1_xcvr_tx_width_atom                              ("CH1_TX_WIDTH_X16"),
		.ch1_xcvr_rx_width_atom                              ("CH1_RX_WIDTH_X16"),
		.ch1_phy_loopback_mode_atom                          ("CH1_LOOPBACK_MODE_DISABLED"),
		.ch1_flux_mode_atom                                  ("CH1_FLUX_MODE_FLUX_MODE_BYPASS"),
		.ch1_tx_sim_mode_atom                                ("CH1_TX_SIM_MODE_DISABLE"),
		.ch1_rx_sim_mode_atom                                ("CH1_RX_SIM_MODE_DISABLE"),
		.ch1_tx_dl_enable_atom                               ("CH1_TX_DL_ENABLE_DISABLE"),
		.ch1_rx_dl_enable_atom                               ("CH1_RX_DL_ENABLE_ENABLE"),
		.ch1_rx_fec_type_used_atom                           ("CH1_RX_FEC_TYPE_USED_NONE"),
		.ch2_xcvr_tx_preloaded_hardware_configs_atom         ("CH2_TX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch2_xcvr_rx_preloaded_hardware_configs_atom         ("CH2_RX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch2_lc_postdiv_sel_atom                             ("CH2_LC_POSTDIV_SEL_SYNTH2"),
		.ch2_sequencer_reg_en_atom                           ("CH2_SEQUENCER_REG_EN_DISABLE"),
		.ch2_rst_mux_static_sel_atom                         ("CH2_RST_MUX_STATIC_SEL_HRC"),
		.ch2_xcvr_tx_prbs_pattern_atom                       (4'b0000),
		.ch2_xcvr_rx_prbs_pattern_atom                       (4'b0011),
		.ch2_xcvr_tx_user_clk_only_mode_atom                 ("CH2_TX_USER_CLK_ONLY_MODE_DISABLE"),
		.ch2_xcvr_tx_width_atom                              ("CH2_TX_WIDTH_X16"),
		.ch2_xcvr_rx_width_atom                              ("CH2_RX_WIDTH_X16"),
		.ch2_phy_loopback_mode_atom                          ("CH2_LOOPBACK_MODE_DISABLED"),
		.ch2_flux_mode_atom                                  ("CH2_FLUX_MODE_FLUX_MODE_BYPASS"),
		.ch2_tx_sim_mode_atom                                ("CH2_TX_SIM_MODE_DISABLE"),
		.ch2_rx_sim_mode_atom                                ("CH2_RX_SIM_MODE_DISABLE"),
		.ch2_tx_dl_enable_atom                               ("CH2_TX_DL_ENABLE_DISABLE"),
		.ch2_rx_dl_enable_atom                               ("CH2_RX_DL_ENABLE_DISABLE"),
		.ch2_rx_fec_type_used_atom                           ("CH2_RX_FEC_TYPE_USED_RS"),
		.ch3_xcvr_tx_preloaded_hardware_configs_atom         ("CH3_TX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch3_xcvr_rx_preloaded_hardware_configs_atom         ("CH3_RX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch3_lc_postdiv_sel_atom                             ("CH3_LC_POSTDIV_SEL_SYNTH2"),
		.ch3_sequencer_reg_en_atom                           ("CH3_SEQUENCER_REG_EN_ENABLE"),
		.ch3_rst_mux_static_sel_atom                         ("CH3_RST_MUX_STATIC_SEL_HRC"),
		.ch3_xcvr_tx_prbs_pattern_atom                       (4'b0000),
		.ch3_xcvr_rx_prbs_pattern_atom                       (4'b0111),
		.ch3_xcvr_tx_user_clk_only_mode_atom                 ("CH3_TX_USER_CLK_ONLY_MODE_DISABLE"),
		.ch3_xcvr_tx_width_atom                              ("CH3_TX_WIDTH_X16"),
		.ch3_xcvr_rx_width_atom                              ("CH3_RX_WIDTH_X16"),
		.ch3_phy_loopback_mode_atom                          ("CH3_LOOPBACK_MODE_DISABLED"),
		.ch3_flux_mode_atom                                  ("CH3_FLUX_MODE_FLUX_MODE_BYPASS"),
		.ch3_tx_sim_mode_atom                                ("CH3_TX_SIM_MODE_DISABLE"),
		.ch3_rx_sim_mode_atom                                ("CH3_RX_SIM_MODE_DISABLE"),
		.ch3_tx_dl_enable_atom                               ("CH3_TX_DL_ENABLE_DISABLE"),
		.ch3_rx_dl_enable_atom                               ("CH3_RX_DL_ENABLE_ENABLE"),
		.ch3_rx_fec_type_used_atom                           ("CH3_RX_FEC_TYPE_USED_RS"),
		.ch0_tx_pll_l_counter_atom                           (6'b000001),
		.ch0_cdr_l_counter_atom                              (6'b000001),
		.ch0_tx_pll_refclk_select_atom                       ("CH0_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch0_cdr_refclk_select_atom                          ("CH0_CDR_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch1_tx_pll_l_counter_atom                           (6'b000001),
		.ch1_cdr_l_counter_atom                              (6'b000001),
		.ch1_tx_pll_refclk_select_atom                       ("CH1_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch1_cdr_refclk_select_atom                          ("CH1_CDR_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch2_tx_pll_l_counter_atom                           (6'b000001),
		.ch2_cdr_l_counter_atom                              (6'b000001),
		.ch2_tx_pll_refclk_select_atom                       ("CH2_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch2_cdr_refclk_select_atom                          ("CH2_CDR_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch3_tx_pll_l_counter_atom                           (6'b000001),
		.ch3_cdr_l_counter_atom                              (6'b000001),
		.ch3_tx_pll_refclk_select_atom                       ("CH3_TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch3_cdr_refclk_select_atom                          ("CH3_CDR_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch0_rx_dl_rx_lat_bit_for_async_atom                 (18'b010100000100010011),
		.ch0_rx_dl_rxbit_cntr_pma_atom                       ("CH0_RX_DL_RXBIT_CNTR_PMA_DISABLE"),
		.ch0_rx_dl_rxbit_rollover_atom                       (18'b111110100100001111),
		.ch1_rx_dl_rx_lat_bit_for_async_atom                 (18'b111110100110100101),
		.ch1_rx_dl_rxbit_cntr_pma_atom                       ("CH1_RX_DL_RXBIT_CNTR_PMA_ENABLE"),
		.ch1_rx_dl_rxbit_rollover_atom                       (18'b001001111001000101),
		.ch2_rx_dl_rx_lat_bit_for_async_atom                 (18'b111010100000111101),
		.ch2_rx_dl_rxbit_cntr_pma_atom                       ("CH2_RX_DL_RXBIT_CNTR_PMA_DISABLE"),
		.ch2_rx_dl_rxbit_rollover_atom                       (18'b111000111110011110),
		.ch3_rx_dl_rx_lat_bit_for_async_atom                 (18'b100000100111100001),
		.ch3_rx_dl_rxbit_cntr_pma_atom                       ("CH3_RX_DL_RXBIT_CNTR_PMA_DISABLE"),
		.ch3_rx_dl_rxbit_rollover_atom                       (18'b001101111001101011),
		.ch0_tx_bond_size_atom                               ("CH0_TX_BOND_SIZE_X4"),
		.ch1_tx_bond_size_atom                               ("CH1_TX_BOND_SIZE_X4"),
		.ch2_tx_bond_size_atom                               ("CH2_TX_BOND_SIZE_X4"),
		.ch3_tx_bond_size_atom                               ("CH3_TX_BOND_SIZE_X4"),
		.pcie_parity_bypass                                  ("true"),
		.rxbuf_limit_bypass                                  (7),
		.maxpayload_size                                     ("MAXPAYLOAD_SIZE_MAX_PAYLOAD_512"),
		.pldclk_rate                                         ("PLDCLK_RATE_FAST"),
		.port_type                                           ("PORT_TYPE_NATIVE_EP"),
		.sris_enable                                         ("SRIS_ENABLE_DISABLED"),
		.sris_mode                                           ("false"),
		.sim_mode                                            ("SIM_MODE_DISABLE_VSIM_MODE"),
		.sup_mode                                            ("SUP_MODE_USER_MODE"),
		.cvp_enable                                          ("CVP_ENABLE_DISABLED"),
		.cii_monitor_en                                      ("CII_MONITOR_EN_DISABLE"),
		.pclk_clk_hz                                         (32'b00111011100110101100101000000000),
		.pf0_cap_link_surprise_down_err_cap                  ("PF0_CAP_LINK_SURPRISE_DOWN_ERR_CAP_DISABLE"),
		.sys_clk_hz                                          (32'b00010100110111001001001110000000),
		.link_rate                                           ("LINK_RATE_GEN4"),
		.link_width                                          ("LINK_WIDTH_X4"),
		.num_of_lanes                                        ("NUM_OF_LANES_NUM_4"),
		.pf0_dsp_16g_tx_preset0                              (7),
		.pf0_dsp_16g_tx_preset1                              (7),
		.pf0_dsp_16g_tx_preset2                              (7),
		.pf0_dsp_16g_tx_preset3                              (7),
		.pf0_dsp_16g_tx_preset4                              (0),
		.pf0_dsp_16g_tx_preset5                              (0),
		.pf0_dsp_16g_tx_preset6                              (0),
		.pf0_dsp_16g_tx_preset7                              (0),
		.pf0_dsp_16g_tx_preset8                              (0),
		.pf0_dsp_16g_tx_preset9                              (0),
		.pf0_dsp_16g_tx_preset10                             (0),
		.pf0_dsp_16g_tx_preset11                             (0),
		.pf0_dsp_16g_tx_preset12                             (0),
		.pf0_dsp_16g_tx_preset13                             (0),
		.pf0_dsp_16g_tx_preset14                             (0),
		.pf0_dsp_16g_tx_preset15                             (0),
		.pf0_dsp_tx_preset0                                  (9),
		.pf0_dsp_tx_preset1                                  (9),
		.pf0_dsp_tx_preset2                                  (9),
		.pf0_dsp_tx_preset3                                  (9),
		.pf0_dsp_tx_preset4                                  (0),
		.pf0_dsp_tx_preset5                                  (0),
		.pf0_dsp_tx_preset6                                  (0),
		.pf0_dsp_tx_preset7                                  (0),
		.pf0_dsp_tx_preset8                                  (0),
		.pf0_dsp_tx_preset9                                  (0),
		.pf0_dsp_tx_preset10                                 (0),
		.pf0_dsp_tx_preset11                                 (0),
		.pf0_dsp_tx_preset12                                 (0),
		.pf0_dsp_tx_preset13                                 (0),
		.pf0_dsp_tx_preset14                                 (0),
		.pf0_dsp_tx_preset15                                 (0),
		.pf0_usp_16g_tx_preset0                              (7),
		.pf0_usp_16g_tx_preset1                              (7),
		.pf0_usp_16g_tx_preset2                              (7),
		.pf0_usp_16g_tx_preset3                              (7),
		.pf0_usp_16g_tx_preset4                              (0),
		.pf0_usp_16g_tx_preset5                              (0),
		.pf0_usp_16g_tx_preset6                              (0),
		.pf0_usp_16g_tx_preset7                              (0),
		.pf0_usp_16g_tx_preset8                              (0),
		.pf0_usp_16g_tx_preset9                              (0),
		.pf0_usp_16g_tx_preset10                             (0),
		.pf0_usp_16g_tx_preset11                             (0),
		.pf0_usp_16g_tx_preset12                             (0),
		.pf0_usp_16g_tx_preset13                             (0),
		.pf0_usp_16g_tx_preset14                             (0),
		.pf0_usp_16g_tx_preset15                             (0),
		.pf0_usp_tx_preset0                                  (9),
		.pf0_usp_tx_preset1                                  (9),
		.pf0_usp_tx_preset2                                  (9),
		.pf0_usp_tx_preset3                                  (9),
		.pf0_usp_tx_preset4                                  (0),
		.pf0_usp_tx_preset5                                  (0),
		.pf0_usp_tx_preset6                                  (0),
		.pf0_usp_tx_preset7                                  (0),
		.pf0_usp_tx_preset8                                  (0),
		.pf0_usp_tx_preset9                                  (0),
		.pf0_usp_tx_preset10                                 (0),
		.pf0_usp_tx_preset11                                 (0),
		.pf0_usp_tx_preset12                                 (0),
		.pf0_usp_tx_preset13                                 (0),
		.pf0_usp_tx_preset14                                 (0),
		.pf0_usp_tx_preset15                                 (0),
		.pf0_pci_type0_bar0_enabled                          ("PF0_PCI_TYPE0_BAR0_ENABLED_ENABLED"),
		.pf0_pci_type0_bar0_mask_31_1                        (32'b00000000000000000111111111111111),
		.pf0_bar0_prefetch                                   ("true"),
		.pf0_bar0_type                                       ("PF0_BAR0_TYPE_BAR_MEM64"),
		.pf0_pci_type0_bar1_enabled                          ("PF0_PCI_TYPE0_BAR1_ENABLED_DISABLED"),
		.pf0_pci_type0_bar1_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf0_bar1_prefetch                                   ("false"),
		.pf0_pci_type0_bar2_enabled                          ("PF0_PCI_TYPE0_BAR2_ENABLED_DISABLED"),
		.pf0_pci_type0_bar2_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf0_bar2_prefetch                                   ("false"),
		.pf0_bar2_type                                       ("PF0_BAR2_TYPE_BAR_MEM32"),
		.pf0_pci_type0_bar3_enabled                          ("PF0_PCI_TYPE0_BAR3_ENABLED_DISABLED"),
		.pf0_pci_type0_bar3_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf0_bar3_prefetch                                   ("false"),
		.pf0_pci_type0_bar4_enabled                          ("PF0_PCI_TYPE0_BAR4_ENABLED_DISABLED"),
		.pf0_pci_type0_bar4_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf0_bar4_prefetch                                   ("false"),
		.pf0_bar4_type                                       ("PF0_BAR4_TYPE_BAR_MEM32"),
		.pf0_pci_type0_bar5_enabled                          ("PF0_PCI_TYPE0_BAR5_ENABLED_DISABLED"),
		.pf0_pci_type0_bar5_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf0_bar5_prefetch                                   ("false"),
		.pf0_rom_bar_enable                                  ("PF0_ROM_BAR_ENABLE_DISABLED"),
		.pf0_rom_mask                                        (0),
		.pf0_rom_bar_enabled                                 ("PF0_ROM_BAR_ENABLED_DISABLED"),
		.pf0_rp_rom_bar_enabled                              ("PF0_RP_ROM_BAR_ENABLED_DISABLED"),
		.pf0_rp_rom_mask                                     (0),
		.pf0_sriov_vf_bar0_enabled                           ("PF0_SRIOV_VF_BAR0_ENABLED_DISABLED"),
		.pf0_sriov_vf_bar0_mask                              (32'b00000000000000000000000000000000),
		.pf0_sriov_vf_bar0_prefetch                          ("false"),
		.pf0_sriov_vf_bar0_type                              ("PF0_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf0_sriov_vf_bar1_enabled                           ("PF0_SRIOV_VF_BAR1_ENABLED_DISABLED"),
		.pf0_sriov_vf_bar1_mask                              (32'b00000000000000000000000000000000),
		.pf0_sriov_vf_bar1_prefetch                          ("false"),
		.pf0_sriov_vf_bar2_enabled                           ("PF0_SRIOV_VF_BAR2_ENABLED_DISABLED"),
		.pf0_sriov_vf_bar2_mask                              (32'b00000000000000000000000000000000),
		.pf0_sriov_vf_bar2_prefetch                          ("false"),
		.pf0_sriov_vf_bar2_type                              ("PF0_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf0_sriov_vf_bar3_enabled                           ("PF0_SRIOV_VF_BAR3_ENABLED_DISABLED"),
		.pf0_sriov_vf_bar3_mask                              (32'b00000000000000000000000000000000),
		.pf0_sriov_vf_bar3_prefetch                          ("false"),
		.pf0_sriov_vf_bar4_enabled                           ("PF0_SRIOV_VF_BAR4_ENABLED_DISABLED"),
		.pf0_sriov_vf_bar4_mask                              (32'b00000000000000000000000000000000),
		.pf0_sriov_vf_bar4_prefetch                          ("false"),
		.pf0_sriov_vf_bar4_type                              ("PF0_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf0_sriov_vf_bar5_enabled                           ("PF0_SRIOV_VF_BAR5_ENABLED_DISABLED"),
		.pf0_sriov_vf_bar5_mask                              (32'b00000000000000000000000000000000),
		.pf0_sriov_vf_bar5_prefetch                          ("false"),
		.pf1_pci_type0_bar0_enabled                          ("PF1_PCI_TYPE0_BAR0_ENABLED_DISABLED"),
		.pf1_pci_type0_bar0_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf1_bar0_prefetch                                   ("false"),
		.pf1_bar0_type                                       ("PF1_BAR0_TYPE_BAR_MEM32"),
		.pf1_pci_type0_bar1_enabled                          ("PF1_PCI_TYPE0_BAR1_ENABLED_DISABLED"),
		.pf1_pci_type0_bar1_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf1_bar1_prefetch                                   ("false"),
		.pf1_pci_type0_bar2_enabled                          ("PF1_PCI_TYPE0_BAR2_ENABLED_DISABLED"),
		.pf1_pci_type0_bar2_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf1_bar2_prefetch                                   ("false"),
		.pf1_bar2_type                                       ("PF1_BAR2_TYPE_BAR_MEM32"),
		.pf1_pci_type0_bar3_enabled                          ("PF1_PCI_TYPE0_BAR3_ENABLED_DISABLED"),
		.pf1_pci_type0_bar3_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf1_bar3_prefetch                                   ("false"),
		.pf1_pci_type0_bar4_enabled                          ("PF1_PCI_TYPE0_BAR4_ENABLED_DISABLED"),
		.pf1_pci_type0_bar4_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf1_bar4_prefetch                                   ("false"),
		.pf1_bar4_type                                       ("PF1_BAR4_TYPE_BAR_MEM32"),
		.pf1_pci_type0_bar5_enabled                          ("PF1_PCI_TYPE0_BAR5_ENABLED_DISABLED"),
		.pf1_pci_type0_bar5_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf1_bar5_prefetch                                   ("false"),
		.pf1_rom_bar_enable                                  ("PF1_ROM_BAR_ENABLE_DISABLED"),
		.pf1_rom_mask                                        (0),
		.pf1_rom_bar_enabled                                 ("PF1_ROM_BAR_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar0_enabled                           ("PF1_SRIOV_VF_BAR0_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar0_mask                              (32'b00000000000000000000000000000000),
		.pf1_sriov_vf_bar0_prefetch                          ("false"),
		.pf1_sriov_vf_bar0_type                              ("PF1_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf1_sriov_vf_bar1_enabled                           ("PF1_SRIOV_VF_BAR1_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar1_mask                              (32'b00000000000000000000000000000000),
		.pf1_sriov_vf_bar1_prefetch                          ("false"),
		.pf1_sriov_vf_bar2_enabled                           ("PF1_SRIOV_VF_BAR2_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar2_mask                              (32'b00000000000000000000000000000000),
		.pf1_sriov_vf_bar2_prefetch                          ("false"),
		.pf1_sriov_vf_bar2_type                              ("PF1_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf1_sriov_vf_bar3_enabled                           ("PF1_SRIOV_VF_BAR3_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar3_mask                              (32'b00000000000000000000000000000000),
		.pf1_sriov_vf_bar3_prefetch                          ("false"),
		.pf1_sriov_vf_bar4_enabled                           ("PF1_SRIOV_VF_BAR4_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar4_mask                              (32'b00000000000000000000000000000000),
		.pf1_sriov_vf_bar4_prefetch                          ("false"),
		.pf1_sriov_vf_bar4_type                              ("PF1_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf1_sriov_vf_bar5_enabled                           ("PF1_SRIOV_VF_BAR5_ENABLED_DISABLED"),
		.pf1_sriov_vf_bar5_mask                              (32'b00000000000000000000000000000000),
		.pf1_sriov_vf_bar5_prefetch                          ("false"),
		.pf2_pci_type0_bar0_enabled                          ("PF2_PCI_TYPE0_BAR0_ENABLED_DISABLED"),
		.pf2_pci_type0_bar0_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf2_bar0_prefetch                                   ("false"),
		.pf2_bar0_type                                       ("PF2_BAR0_TYPE_BAR_MEM32"),
		.pf2_pci_type0_bar1_enabled                          ("PF2_PCI_TYPE0_BAR1_ENABLED_DISABLED"),
		.pf2_pci_type0_bar1_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf2_bar1_prefetch                                   ("false"),
		.pf2_pci_type0_bar2_enabled                          ("PF2_PCI_TYPE0_BAR2_ENABLED_DISABLED"),
		.pf2_pci_type0_bar2_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf2_bar2_prefetch                                   ("false"),
		.pf2_bar2_type                                       ("PF2_BAR2_TYPE_BAR_MEM32"),
		.pf2_pci_type0_bar3_enabled                          ("PF2_PCI_TYPE0_BAR3_ENABLED_DISABLED"),
		.pf2_pci_type0_bar3_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf2_bar3_prefetch                                   ("false"),
		.pf2_pci_type0_bar4_enabled                          ("PF2_PCI_TYPE0_BAR4_ENABLED_DISABLED"),
		.pf2_pci_type0_bar4_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf2_bar4_prefetch                                   ("false"),
		.pf2_bar4_type                                       ("PF2_BAR4_TYPE_BAR_MEM32"),
		.pf2_pci_type0_bar5_enabled                          ("PF2_PCI_TYPE0_BAR5_ENABLED_DISABLED"),
		.pf2_pci_type0_bar5_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf2_bar5_prefetch                                   ("false"),
		.pf2_rom_bar_enable                                  ("PF2_ROM_BAR_ENABLE_DISABLED"),
		.pf2_rom_mask                                        (0),
		.pf2_rom_bar_enabled                                 ("PF2_ROM_BAR_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar0_enabled                           ("PF2_SRIOV_VF_BAR0_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar0_mask                              (32'b00000000000000000000000000000000),
		.pf2_sriov_vf_bar0_prefetch                          ("false"),
		.pf2_sriov_vf_bar0_type                              ("PF2_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf2_sriov_vf_bar1_enabled                           ("PF2_SRIOV_VF_BAR1_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar1_mask                              (32'b00000000000000000000000000000000),
		.pf2_sriov_vf_bar1_prefetch                          ("false"),
		.pf2_sriov_vf_bar2_enabled                           ("PF2_SRIOV_VF_BAR2_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar2_mask                              (32'b00000000000000000000000000000000),
		.pf2_sriov_vf_bar2_prefetch                          ("false"),
		.pf2_sriov_vf_bar2_type                              ("PF2_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf2_sriov_vf_bar3_enabled                           ("PF2_SRIOV_VF_BAR3_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar3_mask                              (32'b00000000000000000000000000000000),
		.pf2_sriov_vf_bar3_prefetch                          ("false"),
		.pf2_sriov_vf_bar4_enabled                           ("PF2_SRIOV_VF_BAR4_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar4_mask                              (32'b00000000000000000000000000000000),
		.pf2_sriov_vf_bar4_prefetch                          ("false"),
		.pf2_sriov_vf_bar4_type                              ("PF2_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf2_sriov_vf_bar5_enabled                           ("PF2_SRIOV_VF_BAR5_ENABLED_DISABLED"),
		.pf2_sriov_vf_bar5_mask                              (32'b00000000000000000000000000000000),
		.pf2_sriov_vf_bar5_prefetch                          ("false"),
		.pf3_pci_type0_bar0_enabled                          ("PF3_PCI_TYPE0_BAR0_ENABLED_DISABLED"),
		.pf3_pci_type0_bar0_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf3_bar0_prefetch                                   ("false"),
		.pf3_bar0_type                                       ("PF3_BAR0_TYPE_BAR_MEM32"),
		.pf3_pci_type0_bar1_enabled                          ("PF3_PCI_TYPE0_BAR1_ENABLED_DISABLED"),
		.pf3_pci_type0_bar1_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf3_bar1_prefetch                                   ("false"),
		.pf3_pci_type0_bar2_enabled                          ("PF3_PCI_TYPE0_BAR2_ENABLED_DISABLED"),
		.pf3_pci_type0_bar2_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf3_bar2_prefetch                                   ("false"),
		.pf3_bar2_type                                       ("PF3_BAR2_TYPE_BAR_MEM32"),
		.pf3_pci_type0_bar3_enabled                          ("PF3_PCI_TYPE0_BAR3_ENABLED_DISABLED"),
		.pf3_pci_type0_bar3_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf3_bar3_prefetch                                   ("false"),
		.pf3_pci_type0_bar4_enabled                          ("PF3_PCI_TYPE0_BAR4_ENABLED_DISABLED"),
		.pf3_pci_type0_bar4_mask_31_1                        (32'b00000000000000000000000000000000),
		.pf3_bar4_prefetch                                   ("false"),
		.pf3_bar4_type                                       ("PF3_BAR4_TYPE_BAR_MEM32"),
		.pf3_pci_type0_bar5_enabled                          ("PF3_PCI_TYPE0_BAR5_ENABLED_DISABLED"),
		.pf3_pci_type0_bar5_mask_31_0                        (32'b00000000000000000000000000000000),
		.pf3_bar5_prefetch                                   ("false"),
		.pf3_rom_bar_enable                                  ("PF3_ROM_BAR_ENABLE_DISABLED"),
		.pf3_rom_mask                                        (0),
		.pf3_rom_bar_enabled                                 ("PF3_ROM_BAR_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar0_enabled                           ("PF3_SRIOV_VF_BAR0_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar0_mask                              (32'b00000000000000000000000000000000),
		.pf3_sriov_vf_bar0_prefetch                          ("false"),
		.pf3_sriov_vf_bar0_type                              ("PF3_SRIOV_VF_BAR0_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf3_sriov_vf_bar1_enabled                           ("PF3_SRIOV_VF_BAR1_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar1_mask                              (32'b00000000000000000000000000000000),
		.pf3_sriov_vf_bar1_prefetch                          ("false"),
		.pf3_sriov_vf_bar2_enabled                           ("PF3_SRIOV_VF_BAR2_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar2_mask                              (32'b00000000000000000000000000000000),
		.pf3_sriov_vf_bar2_prefetch                          ("false"),
		.pf3_sriov_vf_bar2_type                              ("PF3_SRIOV_VF_BAR2_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf3_sriov_vf_bar3_enabled                           ("PF3_SRIOV_VF_BAR3_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar3_mask                              (32'b00000000000000000000000000000000),
		.pf3_sriov_vf_bar3_prefetch                          ("false"),
		.pf3_sriov_vf_bar4_enabled                           ("PF3_SRIOV_VF_BAR4_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar4_mask                              (32'b00000000000000000000000000000000),
		.pf3_sriov_vf_bar4_prefetch                          ("false"),
		.pf3_sriov_vf_bar4_type                              ("PF3_SRIOV_VF_BAR4_TYPE_SRIOV_VF_BAR_MEM32"),
		.pf3_sriov_vf_bar5_enabled                           ("PF3_SRIOV_VF_BAR5_ENABLED_DISABLED"),
		.pf3_sriov_vf_bar5_mask                              (32'b00000000000000000000000000000000),
		.pf3_sriov_vf_bar5_prefetch                          ("false"),
		.pf1_enable                                          ("PF1_ENABLE_DISABLED"),
		.pf2_enable                                          ("PF2_ENABLE_DISABLED"),
		.pf3_enable                                          ("PF3_ENABLE_DISABLED"),
		.pf0_sriov_enable                                    ("PF0_SRIOV_ENABLE_DISABLED"),
		.pf1_sriov_enable                                    ("PF1_SRIOV_ENABLE_DISABLED"),
		.pf2_sriov_enable                                    ("PF2_SRIOV_ENABLE_DISABLED"),
		.pf3_sriov_enable                                    ("PF3_SRIOV_ENABLE_DISABLED"),
		.pf0_sriov_cap_sup_page_size                         (0),
		.pf1_sriov_cap_sup_page_size                         (0),
		.pf2_sriov_cap_sup_page_size                         (0),
		.pf3_sriov_cap_sup_page_size                         (0),
		.pf0_sriov_num_vf                                    (0),
		.pf1_sriov_num_vf                                    (0),
		.pf2_sriov_num_vf                                    (0),
		.pf3_sriov_num_vf                                    (0),
		.pf0_msi_enable                                      ("PF0_MSI_ENABLE_ENABLED"),
		.pf0_pci_msi_ext_data_cap                            ("false"),
		.pf0_pci_msi_ext_data_en                             ("false"),
		.pf0_pci_msi_64_bit_addr_cap                         ("false"),
		.pf0_pci_msi_multiple_msg_cap                        ("PF0_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1"),
		.pf0_msix_enable                                     ("PF0_MSIX_ENABLE_DISABLED"),
		.pf0_pci_msix_table_size                             (0),
		.pf0_pci_msix_table_offset                           (0),
		.pf0_pci_msix_bir                                    (0),
		.pf0_pci_msix_pba                                    (0),
		.pf0_pci_msix_pba_offset                             (0),
		.pf0_pci_msix_table_size_vfcomm_cs2                  (0),
		.pf0_exvf_msix_cap_enable                            ("PF0_EXVF_MSIX_CAP_ENABLE_DISABLED"),
		.exvf_msix_tablesize_pf0                             (0),
		.exvf_msixtable_offset_pf0                           (0),
		.exvf_msixtable_bir_pf0                              (0),
		.exvf_msixpba_offset_pf0                             (0),
		.exvf_msixpba_bir_pf0                                (0),
		.pf1_msi_enable                                      ("PF1_MSI_ENABLE_DISABLED"),
		.pf1_pci_msi_ext_data_cap                            ("false"),
		.pf1_pci_msi_ext_data_en                             ("false"),
		.pf1_pci_msi_64_bit_addr_cap                         ("false"),
		.pf1_pci_msi_multiple_msg_cap                        ("PF1_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1"),
		.pf1_msix_enable                                     ("PF1_MSIX_ENABLE_DISABLED"),
		.pf1_pci_msix_table_size                             (0),
		.pf1_pci_msix_table_offset                           (0),
		.pf1_pci_msix_bir                                    (0),
		.pf1_pci_msix_pba                                    (0),
		.pf1_pci_msix_pba_offset                             (0),
		.pf1_pci_msix_table_size_vfcomm_cs2                  (0),
		.pf1_exvf_msix_cap_enable                            ("PF1_EXVF_MSIX_CAP_ENABLE_DISABLED"),
		.exvf_msix_tablesize_pf1                             (0),
		.exvf_msixtable_offset_pf1                           (0),
		.exvf_msixtable_bir_pf1                              (0),
		.exvf_msixpba_offset_pf1                             (0),
		.exvf_msixpba_bir_pf1                                (0),
		.pf2_msi_enable                                      ("PF2_MSI_ENABLE_DISABLED"),
		.pf2_pci_msi_ext_data_cap                            ("false"),
		.pf2_pci_msi_ext_data_en                             ("false"),
		.pf2_pci_msi_64_bit_addr_cap                         ("false"),
		.pf2_pci_msi_multiple_msg_cap                        ("PF2_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1"),
		.pf2_msix_enable                                     ("PF2_MSIX_ENABLE_DISABLED"),
		.pf2_pci_msix_bir                                    (0),
		.pf2_pci_msix_pba                                    (0),
		.pf2_pci_msix_pba_offset                             (0),
		.pf2_pci_msix_table_offset                           (0),
		.pf2_pci_msix_table_size                             (0),
		.pf2_pci_msix_table_size_vfcomm_cs2                  (0),
		.pf2_exvf_msix_cap_enable                            ("PF2_EXVF_MSIX_CAP_ENABLE_DISABLED"),
		.exvf_msix_tablesize_pf2                             (0),
		.exvf_msixtable_offset_pf2                           (0),
		.exvf_msixtable_bir_pf2                              (0),
		.exvf_msixpba_offset_pf2                             (0),
		.exvf_msixpba_bir_pf2                                (0),
		.pf3_msi_enable                                      ("PF3_MSI_ENABLE_DISABLED"),
		.pf3_pci_msi_ext_data_cap                            ("false"),
		.pf3_pci_msi_ext_data_en                             ("false"),
		.pf3_pci_msi_64_bit_addr_cap                         ("false"),
		.pf3_pci_msi_multiple_msg_cap                        ("PF3_PCI_MSI_MULTIPLE_MSG_CAP_MSI_VEC_1"),
		.pf3_msix_enable                                     ("PF3_MSIX_ENABLE_DISABLED"),
		.pf3_pci_msix_bir                                    (0),
		.pf3_pci_msix_pba                                    (0),
		.pf3_pci_msix_pba_offset                             (0),
		.pf3_pci_msix_table_offset                           (0),
		.pf3_pci_msix_table_size                             (0),
		.pf3_pci_msix_table_size_vfcomm_cs2                  (0),
		.pf3_exvf_msix_cap_enable                            ("PF3_EXVF_MSIX_CAP_ENABLE_DISABLED"),
		.exvf_msix_tablesize_pf3                             (0),
		.exvf_msixtable_offset_pf3                           (0),
		.exvf_msixtable_bir_pf3                              (0),
		.exvf_msixpba_offset_pf3                             (0),
		.exvf_msixpba_bir_pf3                                (0),
		.pf0_prs_ext_cap_enable                              ("PF0_PRS_EXT_CAP_ENABLE_DISABLED"),
		.pf0_prs_ext_cap_outstanding_capacity                (0),
		.pf1_prs_ext_cap_enable                              ("PF1_PRS_EXT_CAP_ENABLE_DISABLED"),
		.pf1_prs_ext_cap_outstanding_capacity                (0),
		.pf2_prs_ext_cap_enable                              ("PF2_PRS_EXT_CAP_ENABLE_DISABLED"),
		.pf2_prs_ext_cap_outstanding_capacity                (0),
		.pf3_prs_ext_cap_enable                              ("PF3_PRS_EXT_CAP_ENABLE_DISABLED"),
		.pf3_prs_ext_cap_outstanding_capacity                (0),
		.pf0_pasid_cap_enable                                ("PF0_PASID_CAP_ENABLE_DISABLED"),
		.pf0_pasid_cap_execute_permission_supported          ("PF0_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED"),
		.pf0_pasid_cap_max_pasid_width                       (0),
		.pf0_pasid_cap_privileged_mode_supported             ("PF0_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED"),
		.pf1_pasid_cap_enable                                ("PF1_PASID_CAP_ENABLE_DISABLED"),
		.pf1_pasid_cap_execute_permission_supported          ("PF1_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED"),
		.pf1_pasid_cap_max_pasid_width                       (0),
		.pf1_pasid_cap_privileged_mode_supported             ("PF1_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED"),
		.pf2_pasid_cap_enable                                ("PF2_PASID_CAP_ENABLE_DISABLED"),
		.pf2_pasid_cap_execute_permission_supported          ("PF2_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED"),
		.pf2_pasid_cap_max_pasid_width                       (0),
		.pf2_pasid_cap_privileged_mode_supported             ("PF2_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED"),
		.pf3_pasid_cap_enable                                ("PF3_PASID_CAP_ENABLE_DISABLED"),
		.pf3_pasid_cap_execute_permission_supported          ("PF3_PASID_CAP_EXECUTE_PERMISSION_SUPPORTED_DISABLED"),
		.pf3_pasid_cap_max_pasid_width                       (0),
		.pf3_pasid_cap_privileged_mode_supported             ("PF3_PASID_CAP_PRIVILEGED_MODE_SUPPORTED_DISABLED"),
		.pf0_sn_cap_enable                                   ("PF0_SN_CAP_ENABLE_DISABLED"),
		.pf0_sn_ser_num_reg_1_dw                             (32'b00000000000000000000000000000000),
		.pf0_sn_ser_num_reg_2_dw                             (32'b00000000000000000000000000000000),
		.pf1_sn_cap_enable                                   ("PF1_SN_CAP_ENABLE_DISABLED"),
		.pf1_sn_ser_num_reg_1_dw                             (32'b00000000000000000000000000000000),
		.pf1_sn_ser_num_reg_2_dw                             (32'b00000000000000000000000000000000),
		.pf2_sn_cap_enable                                   ("PF2_SN_CAP_ENABLE_DISABLED"),
		.pf2_sn_ser_num_reg_1_dw                             (32'b00000000000000000000000000000000),
		.pf2_sn_ser_num_reg_2_dw                             (32'b00000000000000000000000000000000),
		.pf3_sn_cap_enable                                   ("PF3_SN_CAP_ENABLE_DISABLED"),
		.pf3_sn_ser_num_reg_1_dw                             (32'b00000000000000000000000000000000),
		.pf3_sn_ser_num_reg_2_dw                             (32'b00000000000000000000000000000000),
		.pf0_pcie_cap_ep_l0s_accpt_latency                   (0),
		.pf0_pcie_cap_ep_l1_accpt_latency                    (0),
		.pf0_pcie_cap_l0s_exit_latency_commclk_dis           (0),
		.pf0_pcie_cap_l1_exit_latency_commclk_dis            (0),
		.pf1_pcie_cap_ep_l0s_accpt_latency                   (0),
		.pf1_pcie_cap_ep_l1_accpt_latency                    (0),
		.pf1_pcie_cap_l0s_exit_latency_commclk_dis           (0),
		.pf1_pcie_cap_l1_exit_latency_commclk_dis            (0),
		.pf2_pcie_cap_ep_l0s_accpt_latency                   (0),
		.pf2_pcie_cap_ep_l1_accpt_latency                    (0),
		.pf2_pcie_cap_l0s_exit_latency_commclk_dis           (0),
		.pf2_pcie_cap_l1_exit_latency_commclk_dis            (0),
		.pf3_pcie_cap_ep_l0s_accpt_latency                   (0),
		.pf3_pcie_cap_ep_l1_accpt_latency                    (0),
		.pf3_pcie_cap_l0s_exit_latency_commclk_dis           (0),
		.pf3_pcie_cap_l1_exit_latency_commclk_dis            (0),
		.pf0_pcie_cap_flr_cap                                ("PF0_PCIE_CAP_FLR_CAP_NOT_CAPABLE"),
		.pf1_pcie_cap_flr_cap                                ("PF1_PCIE_CAP_FLR_CAP_NOT_CAPABLE"),
		.pf2_pcie_cap_flr_cap                                ("PF2_PCIE_CAP_FLR_CAP_NOT_CAPABLE"),
		.pf3_pcie_cap_flr_cap                                ("PF3_PCIE_CAP_FLR_CAP_NOT_CAPABLE"),
		.pf0_pcie_cap_port_num                               (1),
		.pf1_pcie_cap_port_num                               (0),
		.pf2_pcie_cap_port_num                               (0),
		.pf3_pcie_cap_port_num                               (0),
		.pf0_pcie_cap_slot_clk_config                        ("true"),
		.pf1_pcie_cap_slot_clk_config                        ("false"),
		.pf2_pcie_cap_slot_clk_config                        ("false"),
		.pf3_pcie_cap_slot_clk_config                        ("false"),
		.pf0_ltr_cap_enable                                  ("PF0_LTR_CAP_ENABLE_DISABLED"),
		.pf0_pcie_slot_imp                                   ("PF0_PCIE_SLOT_IMP_NOT_IMPLEMENTED"),
		.pf0_pcie_cap_slot_power_limit_scale                 (0),
		.pf0_pcie_cap_slot_power_limit_value                 (0),
		.pf0_pcie_cap_phy_slot_num                           (0),
		.pf0_pcie_cap_hot_plug_capable                       ("false"),
		.pf0_pcie_cap_ext_tag_en                             ("true"),
		.pf1_pcie_cap_ext_tag_en                             ("false"),
		.pf2_pcie_cap_ext_tag_en                             ("false"),
		.pf3_pcie_cap_ext_tag_en                             ("false"),
		.cfg_ptm_auto_update_signal                          ("false"),
		.ptm_autoupdate                                      ("PTM_AUTOUPDATE_AUTOUPDATE_DISABLE"),
		.ptm_enable                                          ("PTM_ENABLE_DISABLE"),
		.pf0_ats_cap_enable                                  ("PF0_ATS_CAP_ENABLE_DISABLED"),
		.pf0_exvf_ats_cap_enable                             ("PF0_EXVF_ATS_CAP_ENABLE_DISABLED"),
		.pf0_ats_cap_invalidate_q_depth                      (0),
		.pf0_ats_exvf_align_request                          ("PF0_ATS_EXVF_ALIGN_REQUEST_DISABLE"),
		.pf1_ats_cap_enable                                  ("PF1_ATS_CAP_ENABLE_DISABLED"),
		.pf1_exvf_ats_cap_enable                             ("PF1_EXVF_ATS_CAP_ENABLE_DISABLED"),
		.pf1_ats_cap_invalidate_q_depth                      (0),
		.pf1_ats_exvf_align_request                          ("PF1_ATS_EXVF_ALIGN_REQUEST_DISABLE"),
		.pf2_ats_cap_enable                                  ("PF2_ATS_CAP_ENABLE_DISABLED"),
		.pf2_exvf_ats_cap_enable                             ("PF2_EXVF_ATS_CAP_ENABLE_DISABLED"),
		.pf2_ats_cap_invalidate_q_depth                      (0),
		.pf2_ats_exvf_align_request                          ("PF2_ATS_EXVF_ALIGN_REQUEST_DISABLE"),
		.pf3_ats_cap_enable                                  ("PF3_ATS_CAP_ENABLE_DISABLED"),
		.pf3_exvf_ats_cap_enable                             ("PF3_EXVF_ATS_CAP_ENABLE_DISABLED"),
		.pf3_ats_cap_invalidate_q_depth                      (0),
		.pf3_ats_exvf_align_request                          ("PF3_ATS_EXVF_ALIGN_REQUEST_DISABLE"),
		.pf0_tph_cap_enable                                  ("PF0_TPH_CAP_ENABLE_DISABLED"),
		.pf0_tph_req_cap_int_vec                             ("PF0_TPH_REQ_CAP_INT_VEC_DISABLED"),
		.pf0_tph_req_cap_int_vec_vfcomm_cs2                  ("PF0_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED"),
		.pf0_tph_req_cap_st_table_loc_0_vfcomm_cs2           ("PF0_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF"),
		.pf0_tph_req_cap_st_table_loc_1                      ("PF0_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE"),
		.pf0_tph_req_cap_st_table_loc_1_vfcomm_cs2           ("PF0_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF"),
		.pf0_tph_req_cap_st_table_size                       (0),
		.pf0_tph_req_cap_st_table_size_vfcomm_cs2            (0),
		.pf0_tph_req_device_spec                             ("PF0_TPH_REQ_DEVICE_SPEC_DISABLED"),
		.pf0_tph_req_device_spec_vfcomm_cs2                  ("PF0_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED"),
		.pf0_exvf_tph_cap_enable                             ("PF0_EXVF_TPH_CAP_ENABLE_DISABLED"),
		.exvf_tph_sttablelocation_pf0                        (0),
		.exvf_tph_sttablesize_pf0                            (0),
		.pf1_tph_cap_enable                                  ("PF1_TPH_CAP_ENABLE_DISABLED"),
		.pf1_tph_req_cap_int_vec                             ("PF1_TPH_REQ_CAP_INT_VEC_DISABLED"),
		.pf1_tph_req_cap_int_vec_vfcomm_cs2                  ("PF1_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED"),
		.pf1_tph_req_cap_st_table_loc_0_vfcomm_cs2           ("PF1_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF"),
		.pf1_tph_req_cap_st_table_loc_1                      ("PF1_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE"),
		.pf1_tph_req_cap_st_table_loc_1_vfcomm_cs2           ("PF1_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF"),
		.pf1_tph_req_cap_st_table_size                       (0),
		.pf1_tph_req_cap_st_table_size_vfcomm_cs2            (0),
		.pf1_tph_req_device_spec                             ("PF1_TPH_REQ_DEVICE_SPEC_DISABLED"),
		.pf1_tph_req_device_spec_vfcomm_cs2                  ("PF1_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED"),
		.pf1_exvf_tph_cap_enable                             ("PF1_EXVF_TPH_CAP_ENABLE_DISABLED"),
		.exvf_tph_sttablelocation_pf1                        (0),
		.exvf_tph_sttablesize_pf1                            (0),
		.pf2_tph_cap_enable                                  ("PF2_TPH_CAP_ENABLE_DISABLED"),
		.pf2_tph_req_cap_int_vec                             ("PF2_TPH_REQ_CAP_INT_VEC_DISABLED"),
		.pf2_tph_req_cap_int_vec_vfcomm_cs2                  ("PF2_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED"),
		.pf2_tph_req_cap_st_table_loc_0_vfcomm_cs2           ("PF2_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF"),
		.pf2_tph_req_cap_st_table_loc_1                      ("PF2_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE"),
		.pf2_tph_req_cap_st_table_loc_1_vfcomm_cs2           ("PF2_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF"),
		.pf2_tph_req_cap_st_table_size                       (0),
		.pf2_tph_req_cap_st_table_size_vfcomm_cs2            (0),
		.pf2_tph_req_device_spec                             ("PF2_TPH_REQ_DEVICE_SPEC_DISABLED"),
		.pf2_tph_req_device_spec_vfcomm_cs2                  ("PF2_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED"),
		.pf2_exvf_tph_cap_enable                             ("PF2_EXVF_TPH_CAP_ENABLE_DISABLED"),
		.exvf_tph_sttablelocation_pf2                        (0),
		.exvf_tph_sttablesize_pf2                            (0),
		.pf3_tph_cap_enable                                  ("PF3_TPH_CAP_ENABLE_DISABLED"),
		.pf3_tph_req_cap_int_vec                             ("PF3_TPH_REQ_CAP_INT_VEC_DISABLED"),
		.pf3_tph_req_cap_int_vec_vfcomm_cs2                  ("PF3_TPH_REQ_CAP_INT_VEC_VFCOMM_CS2_DISABLED"),
		.pf3_tph_req_cap_st_table_loc_0_vfcomm_cs2           ("PF3_TPH_REQ_CAP_ST_TABLE_LOC_0_VFCOMM_CS2_NOT_IN_TPH_STRUCT_VF"),
		.pf3_tph_req_cap_st_table_loc_1                      ("PF3_TPH_REQ_CAP_ST_TABLE_LOC_1_NOT_IN_MSIX_TABLE"),
		.pf3_tph_req_cap_st_table_loc_1_vfcomm_cs2           ("PF3_TPH_REQ_CAP_ST_TABLE_LOC_1_VFCOMM_CS2_NOT_IN_MSIX_TABLE_VF"),
		.pf3_tph_req_cap_st_table_size                       (0),
		.pf3_tph_req_cap_st_table_size_vfcomm_cs2            (0),
		.pf3_tph_req_device_spec                             ("PF3_TPH_REQ_DEVICE_SPEC_DISABLED"),
		.pf3_tph_req_device_spec_vfcomm_cs2                  ("PF3_TPH_REQ_DEVICE_SPEC_VFCOMM_CS2_DISABLED"),
		.pf3_exvf_tph_cap_enable                             ("PF3_EXVF_TPH_CAP_ENABLE_DISABLED"),
		.exvf_tph_sttablelocation_pf3                        (0),
		.exvf_tph_sttablesize_pf3                            (0),
		.pf0_acs_cap_enable                                  ("PF0_ACS_CAP_ENABLE_DISABLED"),
		.pf0_exvf_acs_cap_enable                             ("PF0_EXVF_ACS_CAP_ENABLE_DISABLED"),
		.pf0_acs_cap_acs_src_valid                           ("PF0_ACS_CAP_ACS_SRC_VALID_DISABLED"),
		.pf0_acs_cap_acs_at_block                            ("PF0_ACS_CAP_ACS_AT_BLOCK_DISABLED"),
		.pf0_acs_cap_acs_p2p_req_redirect                    ("PF0_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED"),
		.pf0_acs_cap_acs_p2p_cpl_redirect                    ("PF0_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED"),
		.pf0_acs_cap_acs_usp_forwarding                      ("PF0_ACS_CAP_ACS_USP_FORWARDING_DISABLED"),
		.pf0_acs_cap_acs_p2p_egress_control                  ("PF0_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED"),
		.pf0_acs_cap_acs_egress_ctrl_size                    (8),
		.pf0_acs_cap_acs_direct_translated_p2p               ("PF0_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED"),
		.pf1_acs_cap_enable                                  ("PF1_ACS_CAP_ENABLE_DISABLED"),
		.pf1_exvf_acs_cap_enable                             ("PF1_EXVF_ACS_CAP_ENABLE_DISABLED"),
		.pf1_acs_cap_acs_src_valid                           ("PF1_ACS_CAP_ACS_SRC_VALID_DISABLED"),
		.pf1_acs_cap_acs_at_block                            ("PF1_ACS_CAP_ACS_AT_BLOCK_DISABLED"),
		.pf1_acs_cap_acs_p2p_req_redirect                    ("PF1_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED"),
		.pf1_acs_cap_acs_p2p_cpl_redirect                    ("PF1_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED"),
		.pf1_acs_cap_acs_usp_forwarding                      ("PF1_ACS_CAP_ACS_USP_FORWARDING_DISABLED"),
		.pf1_acs_cap_acs_p2p_egress_control                  ("PF1_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED"),
		.pf1_acs_cap_acs_egress_ctrl_size                    (8),
		.pf1_acs_cap_acs_direct_translated_p2p               ("PF1_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED"),
		.pf2_acs_cap_enable                                  ("PF2_ACS_CAP_ENABLE_DISABLED"),
		.pf2_exvf_acs_cap_enable                             ("PF2_EXVF_ACS_CAP_ENABLE_DISABLED"),
		.pf2_acs_cap_acs_src_valid                           ("PF2_ACS_CAP_ACS_SRC_VALID_DISABLED"),
		.pf2_acs_cap_acs_at_block                            ("PF2_ACS_CAP_ACS_AT_BLOCK_DISABLED"),
		.pf2_acs_cap_acs_p2p_req_redirect                    ("PF2_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED"),
		.pf2_acs_cap_acs_p2p_cpl_redirect                    ("PF2_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED"),
		.pf2_acs_cap_acs_usp_forwarding                      ("PF2_ACS_CAP_ACS_USP_FORWARDING_DISABLED"),
		.pf2_acs_cap_acs_p2p_egress_control                  ("PF2_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED"),
		.pf2_acs_cap_acs_egress_ctrl_size                    (8),
		.pf2_acs_cap_acs_direct_translated_p2p               ("PF2_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED"),
		.pf3_acs_cap_enable                                  ("PF3_ACS_CAP_ENABLE_DISABLED"),
		.pf3_exvf_acs_cap_enable                             ("PF3_EXVF_ACS_CAP_ENABLE_DISABLED"),
		.pf3_acs_cap_acs_src_valid                           ("PF3_ACS_CAP_ACS_SRC_VALID_DISABLED"),
		.pf3_acs_cap_acs_at_block                            ("PF3_ACS_CAP_ACS_AT_BLOCK_DISABLED"),
		.pf3_acs_cap_acs_p2p_req_redirect                    ("PF3_ACS_CAP_ACS_P2P_REQ_REDIRECT_DISABLED"),
		.pf3_acs_cap_acs_p2p_cpl_redirect                    ("PF3_ACS_CAP_ACS_P2P_CPL_REDIRECT_DISABLED"),
		.pf3_acs_cap_acs_usp_forwarding                      ("PF3_ACS_CAP_ACS_USP_FORWARDING_DISABLED"),
		.pf3_acs_cap_acs_p2p_egress_control                  ("PF3_ACS_CAP_ACS_P2P_EGRESS_CONTROL_DISABLED"),
		.pf3_acs_cap_acs_egress_ctrl_size                    (8),
		.pf3_acs_cap_acs_direct_translated_p2p               ("PF3_ACS_CAP_ACS_DIRECT_TRANSLATED_P2P_DISABLED"),
		.pf0_virtio_en                                       ("PF0_VIRTIO_EN_DISABLED"),
		.pf1_virtio_en                                       ("PF1_VIRTIO_EN_DISABLED"),
		.pf2_virtio_en                                       ("PF2_VIRTIO_EN_DISABLED"),
		.pf3_virtio_en                                       ("PF3_VIRTIO_EN_DISABLED"),
		.pf0_exvf_virtio_en                                  ("PF0_EXVF_VIRTIO_EN_DISABLED"),
		.pf1_exvf_virtio_en                                  ("PF1_EXVF_VIRTIO_EN_DISABLED"),
		.pf2_exvf_virtio_en                                  ("PF2_EXVF_VIRTIO_EN_DISABLED"),
		.pf3_exvf_virtio_en                                  ("PF3_EXVF_VIRTIO_EN_DISABLED"),
		.pf0_pci_type0_device_id                             (0),
		.pf0_pci_type0_vendor_id                             (4466),
		.pf0_revision_id                                     (1),
		.pf0_base_class_code                                 (255),
		.pf0_subclass_code                                   (0),
		.pf0_program_interface                               (0),
		.pf0_subsys_vendor_id                                (0),
		.pf0_subsys_dev_id                                   (0),
		.pf0_sriov_vf_device_id                              (0),
		.exvf_subsysid_pf0                                   (0),
		.pf1_pci_type0_vendor_id                             (0),
		.pf1_pci_type0_device_id                             (0),
		.pf1_revision_id                                     (0),
		.pf1_base_class_code                                 (0),
		.pf1_subclass_code                                   (0),
		.pf1_program_interface                               (0),
		.pf1_subsys_vendor_id                                (0),
		.pf1_subsys_dev_id                                   (0),
		.pf1_sriov_vf_device_id                              (0),
		.exvf_subsysid_pf1                                   (0),
		.pf2_pci_type0_vendor_id                             (0),
		.pf2_pci_type0_device_id                             (0),
		.pf2_revision_id                                     (0),
		.pf2_base_class_code                                 (0),
		.pf2_subclass_code                                   (0),
		.pf2_program_interface                               (0),
		.pf2_subsys_vendor_id                                (0),
		.pf2_subsys_dev_id                                   (0),
		.pf2_sriov_vf_device_id                              (0),
		.exvf_subsysid_pf2                                   (0),
		.pf3_pci_type0_vendor_id                             (0),
		.pf3_pci_type0_device_id                             (0),
		.pf3_revision_id                                     (0),
		.pf3_base_class_code                                 (0),
		.pf3_subclass_code                                   (0),
		.pf3_program_interface                               (0),
		.pf3_subsys_vendor_id                                (0),
		.pf3_subsys_dev_id                                   (0),
		.pf3_sriov_vf_device_id                              (0),
		.exvf_subsysid_pf3                                   (0),
		.vsec_select                                         ("false"),
		.pf0_user_vsec_cap_enable                            ("PF0_USER_VSEC_CAP_ENABLE_DISABLED"),
		.pf1_user_vsec_cap_enable                            ("PF1_USER_VSEC_CAP_ENABLE_DISABLED"),
		.pf2_user_vsec_cap_enable                            ("PF2_USER_VSEC_CAP_ENABLE_DISABLED"),
		.pf3_user_vsec_cap_enable                            ("PF3_USER_VSEC_CAP_ENABLE_DISABLED"),
		.vsec_next_offset                                    (0),
		.pf1_user_vsec_offset                                (0),
		.pf2_user_vsec_offset                                (0),
		.pf3_user_vsec_offset                                (0),
		.cvp_vendor_specific_header_id                       (0),
		.drop_vendor0_msg                                    ("FALSE"),
		.drop_vendor1_msg                                    ("FALSE"),
		.pf0_int_pin                                         ("PF0_INT_PIN_NO_INT"),
		.pf1_int_pin                                         ("PF1_INT_PIN_NO_INT"),
		.pf2_int_pin                                         ("PF2_INT_PIN_NO_INT"),
		.pf3_int_pin                                         ("PF3_INT_PIN_NO_INT"),
		.dtk_mode_en                                         ("DTK_MODE_EN_ENABLE"),
		.hrc_arb_sel                                         ("HRC_ARB_SEL_LOCAL_QUAD_ARB"),
		.num_arb_ip                                          (1),
		.pcie_hrc_pulse_sel                                  (0),
		.pf0_port_logic_fast_link_mode                       ("PF0_PORT_LOGIC_FAST_LINK_MODE_DISABLE"),
		.pf0_prefetch_decode                                 ("PF0_PREFETCH_DECODE_PREF64"),
		.usb_hrc_pulse_sel                                   (0),
		.pcie_pcs_mode                                       ("PCIE_PCS_MODE_PCIE"),
		.sm_hssi_pcie_pcs_clk_mux_0_sel                      ("SEL_SAME_QUAD_PCLK0"),
		.sm_hssi_pcie_pcs_clk_mux_1_sel                      ("SEL_SAME_QUAD_PCLK0"),
		.sm_hssi_pcie_pcs_clk_mux_2_sel                      ("SEL_SAME_QUAD_PCLK0"),
		.sm_hssi_pcie_pcs_clk_mux_3_sel                      ("SEL_SAME_QUAD_PCLK0"),
		.sm_hssi_pcie_pcs_hps_clkmux_0_sel                   ("SEL_HPS_PCS1_ENABLED"),
		.sm_hssi_pcie_pcs_rst_mux_0_sel                      ("SEL_SAME_QUAD_PCS_RST"),
		.sm_hssi_pcie_pcs_rst_mux_1_sel                      ("SEL_SAME_QUAD_PCS_RST"),
		.sm_hssi_pcie_pcs_rst_mux_2_sel                      ("SEL_SAME_QUAD_PCS_RST"),
		.sm_hssi_pcie_pcs_rst_mux_3_sel                      ("SEL_SAME_QUAD_PCS_RST"),
		.sm_hssi_pcie_pcs_tx_mux_0_sel                       ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_tx_mux_1_sel                       ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_tx_mux_2_sel                       ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_tx_mux_3_sel                       ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_hps_demux_0_sel                    ("SEL_HPS_PCS1_ENABLED"),
		.sm_hssi_pcie_pcs_hps_mux_0_sel                      ("SEL_HPS_PCS1_ENABLED"),
		.sm_hssi_pcie_pcs_rx_demux_0_sel                     ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_rx_demux_1_sel                     ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_rx_demux_2_sel                     ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_pcs_rx_demux_3_sel                     ("SEL_SAME_QUAD_PCIE_CTRL"),
		.sm_hssi_pcie_clk_mux_0_sel                          ("SEL_MIDDLE"),
		.sm_hssi_pcie_data_mux_0_sel                         ("SEL_MIDDLE"),
		.sm_hssi_pld_chnl_dp_0_dr_enabled                    ("DR_ENABLED_DR_DISABLED"),
		.sm_hssi_pld_chnl_dp_0_duplex_mode                   ("DUPLEX_MODE_DUPLEX"),
		.sm_hssi_pld_chnl_dp_0_pld_channel_identifier        ("PLD_CHANNEL_IDENTIFIER_PHIP"),
		.sm_hssi_pld_chnl_dp_0_rx_clkout1_divider            ("RX_CLKOUT1_DIVIDER_DIV1"),
		.sm_hssi_pld_chnl_dp_0_rx_clkout2_divider            ("RX_CLKOUT2_DIVIDER_DIV1"),
		.sm_hssi_pld_chnl_dp_0_rx_en                         ("TRUE"),
		.sm_hssi_pld_chnl_dp_0_rx_fifo_mode                  ("RX_FIFO_MODE_PHASE_COMP"),
		.sm_hssi_pld_chnl_dp_0_rx_fifo_width                 ("RX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH"),
		.sm_hssi_pld_chnl_dp_0_rx_fifo_wr_clk_hz             (36'b000000010001111000011010001100000000),
		.sm_hssi_pld_chnl_dp_0_rx_user1_clk_dynamic_mux      ("RX_USER1_CLK_DYNAMIC_MUX_C2"),
		.sm_hssi_pld_chnl_dp_0_rx_user2_clk_dynamic_mux      ("RX_USER2_CLK_DYNAMIC_MUX_UX"),
		.sm_hssi_pld_chnl_dp_0_sup_mode                      ("SUP_MODE_USER_MODE"),
		.sm_hssi_pld_chnl_dp_0_tx_clkout1_divider            ("TX_CLKOUT1_DIVIDER_DIV1"),
		.sm_hssi_pld_chnl_dp_0_tx_clkout2_divider            ("TX_CLKOUT2_DIVIDER_DIV1"),
		.sm_hssi_pld_chnl_dp_0_tx_en                         ("TRUE"),
		.sm_hssi_pld_chnl_dp_0_tx_fifo_mode                  ("TX_FIFO_MODE_PHASE_COMP"),
		.sm_hssi_pld_chnl_dp_0_tx_fifo_rd_clk_hz             (36'b000000010001111000011010001100000000),
		.sm_hssi_pld_chnl_dp_0_tx_fifo_width                 ("TX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH"),
		.sm_hssi_pld_chnl_dp_0_tx_user1_clk_dynamic_mux      ("TX_USER1_CLK_DYNAMIC_MUX_C1"),
		.sm_hssi_pld_chnl_dp_0_tx_user2_clk_dynamic_mux      ("TX_USER2_CLK_DYNAMIC_MUX_UNUSED"),
		.sm_hssi_pld_chnl_dp_0_vc_rx_pldif_wm_en             ("VC_RX_PLDIF_WM_EN_DISABLE"),
		.sm_pld_rx_mux_0_sel                                 ("SEL_PCIE"),
		.sm_pld_tx_demux_0_sel                               ("SEL_PCIE"),
		.sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_sel           ("SEL_PCIE"),
		.sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_sel           ("SEL_PCIE")
	) pcie_hal_top (
		.i_hio_txdata                                (i_hio_txdata),                                                                         //   input,  width = 400,                           i_hio_txdata.data
		.i_hio_txdata_extra                          (i_hio_txdata_extra),                                                                   //   input,   width = 50,                     i_hio_txdata_extra.data
		.i_hio_txdata_fifo_wr_en                     (i_hio_txdata_fifo_wr_en),                                                              //   input,    width = 5,                i_hio_txdata_fifo_wr_en.data
		.i_hio_rxdata_fifo_rd_en                     (i_hio_rxdata_fifo_rd_en),                                                              //   input,    width = 5,                i_hio_rxdata_fifo_rd_en.data
		.i_hio_ptp_rst_n                             (i_hio_ptp_rst_n),                                                                      //   input,    width = 5,                        i_hio_ptp_rst_n.reset
		.i_hio_ehip_rx_rst_n                         (i_hio_ehip_rx_rst_n),                                                                  //   input,    width = 5,                    i_hio_ehip_rx_rst_n.reset
		.i_hio_ehip_tx_rst_n                         (i_hio_ehip_tx_rst_n),                                                                  //   input,    width = 5,                    i_hio_ehip_tx_rst_n.reset
		.i_hio_ehip_signal_ok                        (i_hio_ehip_signal_ok),                                                                 //   input,    width = 5,                   i_hio_ehip_signal_ok.reset
		.i_hio_sfreeze_2_r03f_rx_mac_srfz_n          (i_hio_sfreeze_2_r03f_rx_mac_srfz_n),                                                   //   input,    width = 5,     i_hio_sfreeze_2_r03f_rx_mac_srfz_n.reset
		.i_hio_sfreeze_3_c2f_tx_deskew_srfz_n        (i_hio_sfreeze_3_c2f_tx_deskew_srfz_n),                                                 //   input,    width = 5,   i_hio_sfreeze_3_c2f_tx_deskew_srfz_n.reset
		.i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n          (i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n),                                                   //   input,    width = 5,     i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n.reset
		.i_hio_rstfec_fec_rx_rst_n                   (i_hio_rstfec_fec_rx_rst_n),                                                            //   input,    width = 5,              i_hio_rstfec_fec_rx_rst_n.reset
		.i_hio_rstfec_fec_tx_rst_n                   (i_hio_rstfec_fec_tx_rst_n),                                                            //   input,    width = 5,              i_hio_rstfec_fec_tx_rst_n.reset
		.i_hio_rstfec_fec_csr_ret                    (i_hio_rstfec_fec_csr_ret),                                                             //   input,    width = 5,               i_hio_rstfec_fec_csr_ret.reset
		.i_hio_rstfec_rx_fec_sfrz_n                  (i_hio_rstfec_rx_fec_sfrz_n),                                                           //   input,    width = 5,             i_hio_rstfec_rx_fec_sfrz_n.reset
		.i_hio_rstfec_tx_fec_sfrz_n                  (i_hio_rstfec_tx_fec_sfrz_n),                                                           //   input,    width = 5,             i_hio_rstfec_tx_fec_sfrz_n.reset
		.i_hio_rstxcvrif_xcvrif_rx_rst_n             (i_hio_rstxcvrif_xcvrif_rx_rst_n),                                                      //   input,    width = 5,        i_hio_rstxcvrif_xcvrif_rx_rst_n.reset
		.i_hio_rstxcvrif_xcvrif_tx_rst_n             (i_hio_rstxcvrif_xcvrif_tx_rst_n),                                                      //   input,    width = 5,        i_hio_rstxcvrif_xcvrif_tx_rst_n.reset
		.i_hio_rstxcvrif_xcvrif_signal_ok            (i_hio_rstxcvrif_xcvrif_signal_ok),                                                     //   input,    width = 5,       i_hio_rstxcvrif_xcvrif_signal_ok.reset
		.i_hio_rstxcvrif_rx_xcvrif_sfrz_n            (i_hio_rstxcvrif_rx_xcvrif_sfrz_n),                                                     //   input,    width = 5,       i_hio_rstxcvrif_rx_xcvrif_sfrz_n.reset
		.i_hio_rstxcvrif_tx_xcvrif_sfrz_n            (i_hio_rstxcvrif_tx_xcvrif_sfrz_n),                                                     //   input,    width = 5,       i_hio_rstxcvrif_tx_xcvrif_sfrz_n.reset
		.i_hio_rst_pld_clrhip                        (i_hio_rst_pld_clrhip),                                                                 //   input,    width = 5,                   i_hio_rst_pld_clrhip.reset
		.i_hio_rst_pld_clrpcs                        (i_hio_rst_pld_clrpcs),                                                                 //   input,    width = 5,                   i_hio_rst_pld_clrpcs.reset
		.i_hio_rst_pld_perstn                        (i_hio_rst_pld_perstn),                                                                 //   input,    width = 5,                   i_hio_rst_pld_perstn.reset
		.i_hio_rst_pld_ready                         (i_hio_rst_pld_ready),                                                                  //   input,    width = 5,                    i_hio_rst_pld_ready.reset
		.i_hio_rst_pld_adapter_rx_pld_rst_n          (i_hio_rst_pld_adapter_rx_pld_rst_n),                                                   //   input,    width = 5,     i_hio_rst_pld_adapter_rx_pld_rst_n.reset
		.i_hio_rst_pld_adapter_tx_pld_rst_n          (i_hio_rst_pld_adapter_tx_pld_rst_n),                                                   //   input,    width = 5,     i_hio_rst_pld_adapter_tx_pld_rst_n.reset
		.i_hio_rst_ux_rx_pma_rst_n                   (i_hio_rst_ux_rx_pma_rst_n),                                                            //   input,    width = 5,              i_hio_rst_ux_rx_pma_rst_n.reset
		.i_hio_rst_ux_rx_sfrz                        (i_hio_rst_ux_rx_sfrz),                                                                 //   input,    width = 5,                   i_hio_rst_ux_rx_sfrz.reset
		.i_hio_rst_ux_tx_pma_rst_n                   (i_hio_rst_ux_tx_pma_rst_n),                                                            //   input,    width = 5,              i_hio_rst_ux_tx_pma_rst_n.reset
		.i_hio_pld_reset_clk_row                     (i_hio_pld_reset_clk_row),                                                              //   input,    width = 5,                i_hio_pld_reset_clk_row.reset
		.i_hio_uxquad_async                          (i_hio_uxquad_async),                                                                   //   input,  width = 400,                     i_hio_uxquad_async.data
		.i_hio_uxquad_async_pcie_mux                 (i_hio_uxquad_async_pcie_mux),                                                          //   input,  width = 400,            i_hio_uxquad_async_pcie_mux.data
		.rx_serial_n                                 (rx_serial_n),                                                                          //   input,    width = 4,                            rx_serial_n.data
		.rx_serial_p                                 (rx_serial_p),                                                                          //   input,    width = 4,                            rx_serial_p.data
		.o_hio_txdata_fifo_wr_empty                  (o_hio_txdata_fifo_wr_empty),                                                           //  output,    width = 5,             o_hio_txdata_fifo_wr_empty.data
		.o_hio_txdata_fifo_wr_pempty                 (o_hio_txdata_fifo_wr_pempty),                                                          //  output,    width = 5,            o_hio_txdata_fifo_wr_pempty.data
		.o_hio_txdata_fifo_wr_full                   (o_hio_txdata_fifo_wr_full),                                                            //  output,    width = 5,              o_hio_txdata_fifo_wr_full.data
		.o_hio_txdata_fifo_wr_pfull                  (o_hio_txdata_fifo_wr_pfull),                                                           //  output,    width = 5,             o_hio_txdata_fifo_wr_pfull.data
		.o_hio_rxdata                                (o_hio_rxdata),                                                                         //  output,  width = 400,                           o_hio_rxdata.data
		.o_hio_rxdata_extra                          (o_hio_rxdata_extra),                                                                   //  output,   width = 50,                     o_hio_rxdata_extra.data
		.o_hio_rxdata_fifo_rd_empty                  (o_hio_rxdata_fifo_rd_empty),                                                           //  output,    width = 5,             o_hio_rxdata_fifo_rd_empty.data
		.o_hio_rxdata_fifo_rd_pempty                 (o_hio_rxdata_fifo_rd_pempty),                                                          //  output,    width = 5,            o_hio_rxdata_fifo_rd_pempty.data
		.o_hio_rxdata_fifo_rd_full                   (o_hio_rxdata_fifo_rd_full),                                                            //  output,    width = 5,              o_hio_rxdata_fifo_rd_full.data
		.o_hio_rxdata_fifo_rd_pfull                  (o_hio_rxdata_fifo_rd_pfull),                                                           //  output,    width = 5,             o_hio_rxdata_fifo_rd_pfull.data
		.o_hio_rstepcs_rx_pcs_fully_aligned          (o_hio_rstepcs_rx_pcs_fully_aligned),                                                   //  output,    width = 5,     o_hio_rstepcs_rx_pcs_fully_aligned.reset
		.o_hio_rstfec_fec_rx_rdy_n                   (o_hio_rstfec_fec_rx_rdy_n),                                                            //  output,    width = 5,              o_hio_rstfec_fec_rx_rdy_n.reset
		.o_hio_rst_flux0_cpi_cmn_busy                (o_hio_rst_flux0_cpi_cmn_busy),                                                         //  output,    width = 5,           o_hio_rst_flux0_cpi_cmn_busy.reset
		.o_hio_rst_oflux_rx_srds_rdy                 (o_hio_rst_oflux_rx_srds_rdy),                                                          //  output,    width = 5,            o_hio_rst_oflux_rx_srds_rdy.reset
		.o_hio_rst_ux_all_synthlockstatus            (o_hio_rst_ux_all_synthlockstatus),                                                     //  output,    width = 5,       o_hio_rst_ux_all_synthlockstatus.reset
		.o_hio_rst_ux_octl_pcs_rxstatus              (o_hio_rst_ux_octl_pcs_rxstatus),                                                       //  output,    width = 5,         o_hio_rst_ux_octl_pcs_rxstatus.reset
		.o_hio_rst_ux_octl_pcs_txstatus              (o_hio_rst_ux_octl_pcs_txstatus),                                                       //  output,    width = 5,         o_hio_rst_ux_octl_pcs_txstatus.reset
		.o_hio_rst_ux_rxcdrlock2data                 (o_hio_rst_ux_rxcdrlock2data),                                                          //  output,    width = 5,            o_hio_rst_ux_rxcdrlock2data.reset
		.o_hio_rst_ux_rxcdrlockstatus                (o_hio_rst_ux_rxcdrlockstatus),                                                         //  output,    width = 5,           o_hio_rst_ux_rxcdrlockstatus.reset
		.o_hio_uxquad_async                          (o_hio_uxquad_async),                                                                   //  output,  width = 250,                     o_hio_uxquad_async.data
		.tx_serial_p                                 (tx_serial_p),                                                                          //  output,    width = 4,                            tx_serial_p.data
		.tx_serial_n                                 (tx_serial_n),                                                                          //  output,    width = 4,                            tx_serial_n.data
		.i_hio_txdata_async                          (i_hio_txdata_async),                                                                   //   input,  width = 500,                     i_hio_txdata_async.data
		.i_hio_txdata_direct                         (i_hio_txdata_direct),                                                                  //   input,   width = 50,                    i_hio_txdata_direct.data
		.o_hio_rxdata_async                          (o_hio_rxdata_async),                                                                   //  output,  width = 500,                     o_hio_rxdata_async.data
		.o_hio_rxdata_direct                         (o_hio_rxdata_direct),                                                                  //  output,   width = 50,                    o_hio_rxdata_direct.data
		.ioack_cdrdiv_left_ux_bidir_out              (ioack_cdrdiv_left_ux_bidir_out),                                                       //  output,    width = 4,         ioack_cdrdiv_left_ux_bidir_out.data
		.i_refclk_tx_p                               (i_refclk_tx_p),                                                                        //   input,    width = 1,                          i_refclk_tx_p.clk
		.i_syspll_c0_clk                             (i_syspll_c0_clk),                                                                      //   input,    width = 1,                        i_syspll_c0_clk.clk
		.i_syspll_c1_clk                             (i_syspll_c1_clk),                                                                      //   input,    width = 1,                        i_syspll_c1_clk.clk
		.i_syspll_c2_clk                             (i_syspll_c2_clk),                                                                      //   input,    width = 1,                        i_syspll_c2_clk.clk
		.i_flux_clk                                  (i_flux_clk),                                                                           //   input,    width = 1,                             i_flux_clk.clk
		.i_flux_clk_1                                (i_flux_clk_1),                                                                         //   input,    width = 1,                           i_flux_clk_1.clk
		.i_refclk_rx_p                               (i_refclk_rx_p),                                                                        //   input,    width = 1,                          i_refclk_rx_p.clk
		.i_ss_vccl_syspll_locked                     (i_ss_vccl_syspll_locked),                                                              //   input,    width = 1,                i_ss_vccl_syspll_locked.clk
		.o_hio_pcie_user_rx_clk1_clk                 (o_hio_pcie_user_rx_clk1_clk),                                                          //  output,    width = 1,            o_hio_pcie_user_rx_clk1_clk.clk
		.o_hio_pcie_user_rx_clk2_clk                 (o_hio_pcie_user_rx_clk2_clk),                                                          //  output,    width = 1,            o_hio_pcie_user_rx_clk2_clk.clk
		.o_hio_pcie_user_tx_clk1_clk                 (o_hio_pcie_user_tx_clk1_clk),                                                          //  output,    width = 1,            o_hio_pcie_user_tx_clk1_clk.clk
		.o_hio_pcie_user_tx_clk2_clk                 (o_hio_pcie_user_tx_clk2_clk),                                                          //  output,    width = 1,            o_hio_pcie_user_tx_clk2_clk.clk
		.o_pcs4_pipe_rst_n                           (o_pcs4_pipe_rst_n),                                                                    //  output,    width = 1,                               phip_hal.o_pcs4_pipe_rst_n
		.i_rxpipe4_dirfeedback                       (i_rxpipe4_dirfeedback),                                                                //   input,    width = 6,                                       .i_rxpipe4_dirfeedback
		.i_rxpipe4_linkevaluationfeedbackfiguremerit (i_rxpipe4_linkevaluationfeedbackfiguremerit),                                          //   input,    width = 8,                                       .i_rxpipe4_linkevaluationfeedbackfiguremerit
		.i_rxpipe4_localfs                           (i_rxpipe4_localfs),                                                                    //   input,    width = 6,                                       .i_rxpipe4_localfs
		.i_rxpipe4_locallf                           (i_rxpipe4_locallf),                                                                    //   input,    width = 6,                                       .i_rxpipe4_locallf
		.i_rxpipe4_localtxcoefficientsvalid          (i_rxpipe4_localtxcoefficientsvalid),                                                   //   input,    width = 1,                                       .i_rxpipe4_localtxcoefficientsvalid
		.i_rxpipe4_localtxpresetcoefficients         (i_rxpipe4_localtxpresetcoefficients),                                                  //   input,   width = 18,                                       .i_rxpipe4_localtxpresetcoefficients
		.i_rxpipe4_p2m_bus                           (i_rxpipe4_p2m_bus),                                                                    //   input,    width = 8,                                       .i_rxpipe4_p2m_bus
		.i_rxpipe4_pclkchangeok                      (i_rxpipe4_pclkchangeok),                                                               //   input,    width = 1,                                       .i_rxpipe4_pclkchangeok
		.i_rxpipe4_phystatus                         (i_rxpipe4_phystatus),                                                                  //   input,    width = 1,                                       .i_rxpipe4_phystatus
		.i_rxpipe4_rxdata                            (i_rxpipe4_rxdata),                                                                     //   input,   width = 40,                                       .i_rxpipe4_rxdata
		.i_rxpipe4_rxdatak                           (i_rxpipe4_rxdatak),                                                                    //   input,    width = 4,                                       .i_rxpipe4_rxdatak
		.i_rxpipe4_rxdatavalid                       (i_rxpipe4_rxdatavalid),                                                                //   input,    width = 1,                                       .i_rxpipe4_rxdatavalid
		.i_rxpipe4_rxelecidlea                       (i_rxpipe4_rxelecidlea),                                                                //   input,    width = 1,                                       .i_rxpipe4_rxelecidlea
		.i_rxpipe4_rxstandbystatus                   (i_rxpipe4_rxstandbystatus),                                                            //   input,    width = 1,                                       .i_rxpipe4_rxstandbystatus
		.i_rxpipe4_rxstartblock                      (i_rxpipe4_rxstartblock),                                                               //   input,    width = 1,                                       .i_rxpipe4_rxstartblock
		.i_rxpipe4_rxstatus                          (i_rxpipe4_rxstatus),                                                                   //   input,    width = 3,                                       .i_rxpipe4_rxstatus
		.i_rxpipe4_rxsyncheader                      (i_rxpipe4_rxsyncheader),                                                               //   input,    width = 4,                                       .i_rxpipe4_rxsyncheader
		.i_rxpipe4_rxvalid                           (i_rxpipe4_rxvalid),                                                                    //   input,    width = 1,                                       .i_rxpipe4_rxvalid
		.o_txpipe4_asyncpowerchangeack               (o_txpipe4_asyncpowerchangeack),                                                        //  output,    width = 1,                                       .o_txpipe4_asyncpowerchangeack
		.o_txpipe4_blockaligncontrol                 (o_txpipe4_blockaligncontrol),                                                          //  output,    width = 1,                                       .o_txpipe4_blockaligncontrol
		.o_txpipe4_cfg_hw_auto_sp_dis                (o_txpipe4_cfg_hw_auto_sp_dis),                                                         //  output,    width = 1,                                       .o_txpipe4_cfg_hw_auto_sp_dis
		.o_txpipe4_dirchange                         (o_txpipe4_dirchange),                                                                  //  output,    width = 1,                                       .o_txpipe4_dirchange
		.o_txpipe4_ebuf_mode                         (o_txpipe4_ebuf_mode),                                                                  //  output,    width = 1,                                       .o_txpipe4_ebuf_mode
		.o_txpipe4_encodedecodebypass                (o_txpipe4_encodedecodebypass),                                                         //  output,    width = 1,                                       .o_txpipe4_encodedecodebypass
		.o_txpipe4_fs                                (o_txpipe4_fs),                                                                         //  output,    width = 6,                                       .o_txpipe4_fs
		.o_txpipe4_getlocalpresetcoefficients        (o_txpipe4_getlocalpresetcoefficients),                                                 //  output,    width = 1,                                       .o_txpipe4_getlocalpresetcoefficients
		.o_txpipe4_invalidrequest                    (o_txpipe4_invalidrequest),                                                             //  output,    width = 1,                                       .o_txpipe4_invalidrequest
		.o_txpipe4_lf                                (o_txpipe4_lf),                                                                         //  output,    width = 6,                                       .o_txpipe4_lf
		.o_txpipe4_localpresetindex                  (o_txpipe4_localpresetindex),                                                           //  output,    width = 5,                                       .o_txpipe4_localpresetindex
		.o_txpipe4_lowpin_nt                         (o_txpipe4_lowpin_nt),                                                                  //  output,    width = 1,                                       .o_txpipe4_lowpin_nt
		.o_txpipe4_m2p_bus                           (o_txpipe4_m2p_bus),                                                                    //  output,    width = 8,                                       .o_txpipe4_m2p_bus
		.o_txpipe4_pclk_rate                         (o_txpipe4_pclk_rate),                                                                  //  output,    width = 3,                                       .o_txpipe4_pclk_rate
		.o_txpipe4_pclkchangeack                     (o_txpipe4_pclkchangeack),                                                              //  output,    width = 1,                                       .o_txpipe4_pclkchangeack
		.o_txpipe4_phy_mode_nt                       (o_txpipe4_phy_mode_nt),                                                                //  output,    width = 4,                                       .o_txpipe4_phy_mode_nt
		.o_txpipe4_powerdown                         (o_txpipe4_powerdown),                                                                  //  output,    width = 4,                                       .o_txpipe4_powerdown
		.o_txpipe4_rate                              (o_txpipe4_rate),                                                                       //  output,    width = 3,                                       .o_txpipe4_rate
		.o_txpipe4_rxelecidle_disable_a              (o_txpipe4_rxelecidle_disable_a),                                                       //  output,    width = 1,                                       .o_txpipe4_rxelecidle_disable_a
		.o_txpipe4_rxeqclr                           (o_txpipe4_rxeqclr),                                                                    //  output,    width = 1,                                       .o_txpipe4_rxeqclr
		.o_txpipe4_rxeqeval                          (o_txpipe4_rxeqeval),                                                                   //  output,    width = 1,                                       .o_txpipe4_rxeqeval
		.o_txpipe4_rxeqinprogress                    (o_txpipe4_rxeqinprogress),                                                             //  output,    width = 1,                                       .o_txpipe4_rxeqinprogress
		.o_txpipe4_rxeqtraining                      (o_txpipe4_rxeqtraining),                                                               //  output,    width = 1,                                       .o_txpipe4_rxeqtraining
		.o_txpipe4_rxpolarity                        (o_txpipe4_rxpolarity),                                                                 //  output,    width = 1,                                       .o_txpipe4_rxpolarity
		.o_txpipe4_rxpresethint                      (o_txpipe4_rxpresethint),                                                               //  output,    width = 3,                                       .o_txpipe4_rxpresethint
		.o_txpipe4_rxstandby                         (o_txpipe4_rxstandby),                                                                  //  output,    width = 1,                                       .o_txpipe4_rxstandby
		.o_txpipe4_rxtermination                     (o_txpipe4_rxtermination),                                                              //  output,    width = 1,                                       .o_txpipe4_rxtermination
		.o_txpipe4_srisenable                        (o_txpipe4_srisenable),                                                                 //  output,    width = 1,                                       .o_txpipe4_srisenable
		.o_txpipe4_txcmnmode_disable_a               (o_txpipe4_txcmnmode_disable_a),                                                        //  output,    width = 1,                                       .o_txpipe4_txcmnmode_disable_a
		.o_txpipe4_txcompliance                      (o_txpipe4_txcompliance),                                                               //  output,    width = 1,                                       .o_txpipe4_txcompliance
		.o_txpipe4_txdata                            (o_txpipe4_txdata),                                                                     //  output,   width = 40,                                       .o_txpipe4_txdata
		.o_txpipe4_txdatak                           (o_txpipe4_txdatak),                                                                    //  output,    width = 4,                                       .o_txpipe4_txdatak
		.o_txpipe4_txdatavalid                       (o_txpipe4_txdatavalid),                                                                //  output,    width = 1,                                       .o_txpipe4_txdatavalid
		.o_txpipe4_txdeemph                          (o_txpipe4_txdeemph),                                                                   //  output,   width = 18,                                       .o_txpipe4_txdeemph
		.o_txpipe4_txdtctrx_lb                       (o_txpipe4_txdtctrx_lb),                                                                //  output,    width = 1,                                       .o_txpipe4_txdtctrx_lb
		.o_txpipe4_txelecidle                        (o_txpipe4_txelecidle),                                                                 //  output,    width = 1,                                       .o_txpipe4_txelecidle
		.o_txpipe4_txmargin                          (o_txpipe4_txmargin),                                                                   //  output,    width = 3,                                       .o_txpipe4_txmargin
		.o_txpipe4_txoneszeros                       (o_txpipe4_txoneszeros),                                                                //  output,    width = 1,                                       .o_txpipe4_txoneszeros
		.o_txpipe4_txstartblock                      (o_txpipe4_txstartblock),                                                               //  output,    width = 1,                                       .o_txpipe4_txstartblock
		.o_txpipe4_txswing                           (o_txpipe4_txswing),                                                                    //  output,    width = 1,                                       .o_txpipe4_txswing
		.o_txpipe4_txsyncheader                      (o_txpipe4_txsyncheader),                                                               //  output,    width = 4,                                       .o_txpipe4_txsyncheader
		.o_txpipe4_width                             (o_txpipe4_width),                                                                      //  output,    width = 3,                                       .o_txpipe4_width
		.o_pcs5_pipe_rst_n                           (o_pcs5_pipe_rst_n),                                                                    //  output,    width = 1,                                       .o_pcs5_pipe_rst_n
		.i_rxpipe5_dirfeedback                       (i_rxpipe5_dirfeedback),                                                                //   input,    width = 6,                                       .i_rxpipe5_dirfeedback
		.i_rxpipe5_linkevaluationfeedbackfiguremerit (i_rxpipe5_linkevaluationfeedbackfiguremerit),                                          //   input,    width = 8,                                       .i_rxpipe5_linkevaluationfeedbackfiguremerit
		.i_rxpipe5_localfs                           (i_rxpipe5_localfs),                                                                    //   input,    width = 6,                                       .i_rxpipe5_localfs
		.i_rxpipe5_locallf                           (i_rxpipe5_locallf),                                                                    //   input,    width = 6,                                       .i_rxpipe5_locallf
		.i_rxpipe5_localtxcoefficientsvalid          (i_rxpipe5_localtxcoefficientsvalid),                                                   //   input,    width = 1,                                       .i_rxpipe5_localtxcoefficientsvalid
		.i_rxpipe5_localtxpresetcoefficients         (i_rxpipe5_localtxpresetcoefficients),                                                  //   input,   width = 18,                                       .i_rxpipe5_localtxpresetcoefficients
		.i_rxpipe5_p2m_bus                           (i_rxpipe5_p2m_bus),                                                                    //   input,    width = 8,                                       .i_rxpipe5_p2m_bus
		.i_rxpipe5_pclkchangeok                      (i_rxpipe5_pclkchangeok),                                                               //   input,    width = 1,                                       .i_rxpipe5_pclkchangeok
		.i_rxpipe5_phystatus                         (i_rxpipe5_phystatus),                                                                  //   input,    width = 1,                                       .i_rxpipe5_phystatus
		.i_rxpipe5_rxdata                            (i_rxpipe5_rxdata),                                                                     //   input,   width = 40,                                       .i_rxpipe5_rxdata
		.i_rxpipe5_rxdatak                           (i_rxpipe5_rxdatak),                                                                    //   input,    width = 4,                                       .i_rxpipe5_rxdatak
		.i_rxpipe5_rxdatavalid                       (i_rxpipe5_rxdatavalid),                                                                //   input,    width = 1,                                       .i_rxpipe5_rxdatavalid
		.i_rxpipe5_rxelecidlea                       (i_rxpipe5_rxelecidlea),                                                                //   input,    width = 1,                                       .i_rxpipe5_rxelecidlea
		.i_rxpipe5_rxstandbystatus                   (i_rxpipe5_rxstandbystatus),                                                            //   input,    width = 1,                                       .i_rxpipe5_rxstandbystatus
		.i_rxpipe5_rxstartblock                      (i_rxpipe5_rxstartblock),                                                               //   input,    width = 1,                                       .i_rxpipe5_rxstartblock
		.i_rxpipe5_rxstatus                          (i_rxpipe5_rxstatus),                                                                   //   input,    width = 3,                                       .i_rxpipe5_rxstatus
		.i_rxpipe5_rxsyncheader                      (i_rxpipe5_rxsyncheader),                                                               //   input,    width = 4,                                       .i_rxpipe5_rxsyncheader
		.i_rxpipe5_rxvalid                           (i_rxpipe5_rxvalid),                                                                    //   input,    width = 1,                                       .i_rxpipe5_rxvalid
		.o_txpipe5_asyncpowerchangeack               (o_txpipe5_asyncpowerchangeack),                                                        //  output,    width = 1,                                       .o_txpipe5_asyncpowerchangeack
		.o_txpipe5_blockaligncontrol                 (o_txpipe5_blockaligncontrol),                                                          //  output,    width = 1,                                       .o_txpipe5_blockaligncontrol
		.o_txpipe5_cfg_hw_auto_sp_dis                (o_txpipe5_cfg_hw_auto_sp_dis),                                                         //  output,    width = 1,                                       .o_txpipe5_cfg_hw_auto_sp_dis
		.o_txpipe5_dirchange                         (o_txpipe5_dirchange),                                                                  //  output,    width = 1,                                       .o_txpipe5_dirchange
		.o_txpipe5_ebuf_mode                         (o_txpipe5_ebuf_mode),                                                                  //  output,    width = 1,                                       .o_txpipe5_ebuf_mode
		.o_txpipe5_encodedecodebypass                (o_txpipe5_encodedecodebypass),                                                         //  output,    width = 1,                                       .o_txpipe5_encodedecodebypass
		.o_txpipe5_fs                                (o_txpipe5_fs),                                                                         //  output,    width = 6,                                       .o_txpipe5_fs
		.o_txpipe5_getlocalpresetcoefficients        (o_txpipe5_getlocalpresetcoefficients),                                                 //  output,    width = 1,                                       .o_txpipe5_getlocalpresetcoefficients
		.o_txpipe5_invalidrequest                    (o_txpipe5_invalidrequest),                                                             //  output,    width = 1,                                       .o_txpipe5_invalidrequest
		.o_txpipe5_lf                                (o_txpipe5_lf),                                                                         //  output,    width = 6,                                       .o_txpipe5_lf
		.o_txpipe5_localpresetindex                  (o_txpipe5_localpresetindex),                                                           //  output,    width = 5,                                       .o_txpipe5_localpresetindex
		.o_txpipe5_lowpin_nt                         (o_txpipe5_lowpin_nt),                                                                  //  output,    width = 1,                                       .o_txpipe5_lowpin_nt
		.o_txpipe5_m2p_bus                           (o_txpipe5_m2p_bus),                                                                    //  output,    width = 8,                                       .o_txpipe5_m2p_bus
		.o_txpipe5_pclk_rate                         (o_txpipe5_pclk_rate),                                                                  //  output,    width = 3,                                       .o_txpipe5_pclk_rate
		.o_txpipe5_pclkchangeack                     (o_txpipe5_pclkchangeack),                                                              //  output,    width = 1,                                       .o_txpipe5_pclkchangeack
		.o_txpipe5_phy_mode_nt                       (o_txpipe5_phy_mode_nt),                                                                //  output,    width = 4,                                       .o_txpipe5_phy_mode_nt
		.o_txpipe5_powerdown                         (o_txpipe5_powerdown),                                                                  //  output,    width = 4,                                       .o_txpipe5_powerdown
		.o_txpipe5_rate                              (o_txpipe5_rate),                                                                       //  output,    width = 3,                                       .o_txpipe5_rate
		.o_txpipe5_rxelecidle_disable_a              (o_txpipe5_rxelecidle_disable_a),                                                       //  output,    width = 1,                                       .o_txpipe5_rxelecidle_disable_a
		.o_txpipe5_rxeqclr                           (o_txpipe5_rxeqclr),                                                                    //  output,    width = 1,                                       .o_txpipe5_rxeqclr
		.o_txpipe5_rxeqeval                          (o_txpipe5_rxeqeval),                                                                   //  output,    width = 1,                                       .o_txpipe5_rxeqeval
		.o_txpipe5_rxeqinprogress                    (o_txpipe5_rxeqinprogress),                                                             //  output,    width = 1,                                       .o_txpipe5_rxeqinprogress
		.o_txpipe5_rxeqtraining                      (o_txpipe5_rxeqtraining),                                                               //  output,    width = 1,                                       .o_txpipe5_rxeqtraining
		.o_txpipe5_rxpolarity                        (o_txpipe5_rxpolarity),                                                                 //  output,    width = 1,                                       .o_txpipe5_rxpolarity
		.o_txpipe5_rxpresethint                      (o_txpipe5_rxpresethint),                                                               //  output,    width = 3,                                       .o_txpipe5_rxpresethint
		.o_txpipe5_rxstandby                         (o_txpipe5_rxstandby),                                                                  //  output,    width = 1,                                       .o_txpipe5_rxstandby
		.o_txpipe5_rxtermination                     (o_txpipe5_rxtermination),                                                              //  output,    width = 1,                                       .o_txpipe5_rxtermination
		.o_txpipe5_srisenable                        (o_txpipe5_srisenable),                                                                 //  output,    width = 1,                                       .o_txpipe5_srisenable
		.o_txpipe5_txcmnmode_disable_a               (o_txpipe5_txcmnmode_disable_a),                                                        //  output,    width = 1,                                       .o_txpipe5_txcmnmode_disable_a
		.o_txpipe5_txcompliance                      (o_txpipe5_txcompliance),                                                               //  output,    width = 1,                                       .o_txpipe5_txcompliance
		.o_txpipe5_txdata                            (o_txpipe5_txdata),                                                                     //  output,   width = 40,                                       .o_txpipe5_txdata
		.o_txpipe5_txdatak                           (o_txpipe5_txdatak),                                                                    //  output,    width = 4,                                       .o_txpipe5_txdatak
		.o_txpipe5_txdatavalid                       (o_txpipe5_txdatavalid),                                                                //  output,    width = 1,                                       .o_txpipe5_txdatavalid
		.o_txpipe5_txdeemph                          (o_txpipe5_txdeemph),                                                                   //  output,   width = 18,                                       .o_txpipe5_txdeemph
		.o_txpipe5_txdtctrx_lb                       (o_txpipe5_txdtctrx_lb),                                                                //  output,    width = 1,                                       .o_txpipe5_txdtctrx_lb
		.o_txpipe5_txelecidle                        (o_txpipe5_txelecidle),                                                                 //  output,    width = 1,                                       .o_txpipe5_txelecidle
		.o_txpipe5_txmargin                          (o_txpipe5_txmargin),                                                                   //  output,    width = 3,                                       .o_txpipe5_txmargin
		.o_txpipe5_txoneszeros                       (o_txpipe5_txoneszeros),                                                                //  output,    width = 1,                                       .o_txpipe5_txoneszeros
		.o_txpipe5_txstartblock                      (o_txpipe5_txstartblock),                                                               //  output,    width = 1,                                       .o_txpipe5_txstartblock
		.o_txpipe5_txswing                           (o_txpipe5_txswing),                                                                    //  output,    width = 1,                                       .o_txpipe5_txswing
		.o_txpipe5_txsyncheader                      (o_txpipe5_txsyncheader),                                                               //  output,    width = 4,                                       .o_txpipe5_txsyncheader
		.o_txpipe5_width                             (o_txpipe5_width),                                                                      //  output,    width = 3,                                       .o_txpipe5_width
		.o_pcs6_pipe_rst_n                           (o_pcs6_pipe_rst_n),                                                                    //  output,    width = 1,                                       .o_pcs6_pipe_rst_n
		.i_rxpipe6_dirfeedback                       (i_rxpipe6_dirfeedback),                                                                //   input,    width = 6,                                       .i_rxpipe6_dirfeedback
		.i_rxpipe6_linkevaluationfeedbackfiguremerit (i_rxpipe6_linkevaluationfeedbackfiguremerit),                                          //   input,    width = 8,                                       .i_rxpipe6_linkevaluationfeedbackfiguremerit
		.i_rxpipe6_localfs                           (i_rxpipe6_localfs),                                                                    //   input,    width = 6,                                       .i_rxpipe6_localfs
		.i_rxpipe6_locallf                           (i_rxpipe6_locallf),                                                                    //   input,    width = 6,                                       .i_rxpipe6_locallf
		.i_rxpipe6_localtxcoefficientsvalid          (i_rxpipe6_localtxcoefficientsvalid),                                                   //   input,    width = 1,                                       .i_rxpipe6_localtxcoefficientsvalid
		.i_rxpipe6_localtxpresetcoefficients         (i_rxpipe6_localtxpresetcoefficients),                                                  //   input,   width = 18,                                       .i_rxpipe6_localtxpresetcoefficients
		.i_rxpipe6_p2m_bus                           (i_rxpipe6_p2m_bus),                                                                    //   input,    width = 8,                                       .i_rxpipe6_p2m_bus
		.i_rxpipe6_pclkchangeok                      (i_rxpipe6_pclkchangeok),                                                               //   input,    width = 1,                                       .i_rxpipe6_pclkchangeok
		.i_rxpipe6_phystatus                         (i_rxpipe6_phystatus),                                                                  //   input,    width = 1,                                       .i_rxpipe6_phystatus
		.i_rxpipe6_rxdata                            (i_rxpipe6_rxdata),                                                                     //   input,   width = 40,                                       .i_rxpipe6_rxdata
		.i_rxpipe6_rxdatak                           (i_rxpipe6_rxdatak),                                                                    //   input,    width = 4,                                       .i_rxpipe6_rxdatak
		.i_rxpipe6_rxdatavalid                       (i_rxpipe6_rxdatavalid),                                                                //   input,    width = 1,                                       .i_rxpipe6_rxdatavalid
		.i_rxpipe6_rxelecidlea                       (i_rxpipe6_rxelecidlea),                                                                //   input,    width = 1,                                       .i_rxpipe6_rxelecidlea
		.i_rxpipe6_rxstandbystatus                   (i_rxpipe6_rxstandbystatus),                                                            //   input,    width = 1,                                       .i_rxpipe6_rxstandbystatus
		.i_rxpipe6_rxstartblock                      (i_rxpipe6_rxstartblock),                                                               //   input,    width = 1,                                       .i_rxpipe6_rxstartblock
		.i_rxpipe6_rxstatus                          (i_rxpipe6_rxstatus),                                                                   //   input,    width = 3,                                       .i_rxpipe6_rxstatus
		.i_rxpipe6_rxsyncheader                      (i_rxpipe6_rxsyncheader),                                                               //   input,    width = 4,                                       .i_rxpipe6_rxsyncheader
		.i_rxpipe6_rxvalid                           (i_rxpipe6_rxvalid),                                                                    //   input,    width = 1,                                       .i_rxpipe6_rxvalid
		.o_txpipe6_asyncpowerchangeack               (o_txpipe6_asyncpowerchangeack),                                                        //  output,    width = 1,                                       .o_txpipe6_asyncpowerchangeack
		.o_txpipe6_blockaligncontrol                 (o_txpipe6_blockaligncontrol),                                                          //  output,    width = 1,                                       .o_txpipe6_blockaligncontrol
		.o_txpipe6_cfg_hw_auto_sp_dis                (o_txpipe6_cfg_hw_auto_sp_dis),                                                         //  output,    width = 1,                                       .o_txpipe6_cfg_hw_auto_sp_dis
		.o_txpipe6_dirchange                         (o_txpipe6_dirchange),                                                                  //  output,    width = 1,                                       .o_txpipe6_dirchange
		.o_txpipe6_ebuf_mode                         (o_txpipe6_ebuf_mode),                                                                  //  output,    width = 1,                                       .o_txpipe6_ebuf_mode
		.o_txpipe6_encodedecodebypass                (o_txpipe6_encodedecodebypass),                                                         //  output,    width = 1,                                       .o_txpipe6_encodedecodebypass
		.o_txpipe6_fs                                (o_txpipe6_fs),                                                                         //  output,    width = 6,                                       .o_txpipe6_fs
		.o_txpipe6_getlocalpresetcoefficients        (o_txpipe6_getlocalpresetcoefficients),                                                 //  output,    width = 1,                                       .o_txpipe6_getlocalpresetcoefficients
		.o_txpipe6_invalidrequest                    (o_txpipe6_invalidrequest),                                                             //  output,    width = 1,                                       .o_txpipe6_invalidrequest
		.o_txpipe6_lf                                (o_txpipe6_lf),                                                                         //  output,    width = 6,                                       .o_txpipe6_lf
		.o_txpipe6_localpresetindex                  (o_txpipe6_localpresetindex),                                                           //  output,    width = 5,                                       .o_txpipe6_localpresetindex
		.o_txpipe6_lowpin_nt                         (o_txpipe6_lowpin_nt),                                                                  //  output,    width = 1,                                       .o_txpipe6_lowpin_nt
		.o_txpipe6_m2p_bus                           (o_txpipe6_m2p_bus),                                                                    //  output,    width = 8,                                       .o_txpipe6_m2p_bus
		.o_txpipe6_pclk_rate                         (o_txpipe6_pclk_rate),                                                                  //  output,    width = 3,                                       .o_txpipe6_pclk_rate
		.o_txpipe6_pclkchangeack                     (o_txpipe6_pclkchangeack),                                                              //  output,    width = 1,                                       .o_txpipe6_pclkchangeack
		.o_txpipe6_phy_mode_nt                       (o_txpipe6_phy_mode_nt),                                                                //  output,    width = 4,                                       .o_txpipe6_phy_mode_nt
		.o_txpipe6_powerdown                         (o_txpipe6_powerdown),                                                                  //  output,    width = 4,                                       .o_txpipe6_powerdown
		.o_txpipe6_rate                              (o_txpipe6_rate),                                                                       //  output,    width = 3,                                       .o_txpipe6_rate
		.o_txpipe6_rxelecidle_disable_a              (o_txpipe6_rxelecidle_disable_a),                                                       //  output,    width = 1,                                       .o_txpipe6_rxelecidle_disable_a
		.o_txpipe6_rxeqclr                           (o_txpipe6_rxeqclr),                                                                    //  output,    width = 1,                                       .o_txpipe6_rxeqclr
		.o_txpipe6_rxeqeval                          (o_txpipe6_rxeqeval),                                                                   //  output,    width = 1,                                       .o_txpipe6_rxeqeval
		.o_txpipe6_rxeqinprogress                    (o_txpipe6_rxeqinprogress),                                                             //  output,    width = 1,                                       .o_txpipe6_rxeqinprogress
		.o_txpipe6_rxeqtraining                      (o_txpipe6_rxeqtraining),                                                               //  output,    width = 1,                                       .o_txpipe6_rxeqtraining
		.o_txpipe6_rxpolarity                        (o_txpipe6_rxpolarity),                                                                 //  output,    width = 1,                                       .o_txpipe6_rxpolarity
		.o_txpipe6_rxpresethint                      (o_txpipe6_rxpresethint),                                                               //  output,    width = 3,                                       .o_txpipe6_rxpresethint
		.o_txpipe6_rxstandby                         (o_txpipe6_rxstandby),                                                                  //  output,    width = 1,                                       .o_txpipe6_rxstandby
		.o_txpipe6_rxtermination                     (o_txpipe6_rxtermination),                                                              //  output,    width = 1,                                       .o_txpipe6_rxtermination
		.o_txpipe6_srisenable                        (o_txpipe6_srisenable),                                                                 //  output,    width = 1,                                       .o_txpipe6_srisenable
		.o_txpipe6_txcmnmode_disable_a               (o_txpipe6_txcmnmode_disable_a),                                                        //  output,    width = 1,                                       .o_txpipe6_txcmnmode_disable_a
		.o_txpipe6_txcompliance                      (o_txpipe6_txcompliance),                                                               //  output,    width = 1,                                       .o_txpipe6_txcompliance
		.o_txpipe6_txdata                            (o_txpipe6_txdata),                                                                     //  output,   width = 40,                                       .o_txpipe6_txdata
		.o_txpipe6_txdatak                           (o_txpipe6_txdatak),                                                                    //  output,    width = 4,                                       .o_txpipe6_txdatak
		.o_txpipe6_txdatavalid                       (o_txpipe6_txdatavalid),                                                                //  output,    width = 1,                                       .o_txpipe6_txdatavalid
		.o_txpipe6_txdeemph                          (o_txpipe6_txdeemph),                                                                   //  output,   width = 18,                                       .o_txpipe6_txdeemph
		.o_txpipe6_txdtctrx_lb                       (o_txpipe6_txdtctrx_lb),                                                                //  output,    width = 1,                                       .o_txpipe6_txdtctrx_lb
		.o_txpipe6_txelecidle                        (o_txpipe6_txelecidle),                                                                 //  output,    width = 1,                                       .o_txpipe6_txelecidle
		.o_txpipe6_txmargin                          (o_txpipe6_txmargin),                                                                   //  output,    width = 3,                                       .o_txpipe6_txmargin
		.o_txpipe6_txoneszeros                       (o_txpipe6_txoneszeros),                                                                //  output,    width = 1,                                       .o_txpipe6_txoneszeros
		.o_txpipe6_txstartblock                      (o_txpipe6_txstartblock),                                                               //  output,    width = 1,                                       .o_txpipe6_txstartblock
		.o_txpipe6_txswing                           (o_txpipe6_txswing),                                                                    //  output,    width = 1,                                       .o_txpipe6_txswing
		.o_txpipe6_txsyncheader                      (o_txpipe6_txsyncheader),                                                               //  output,    width = 4,                                       .o_txpipe6_txsyncheader
		.o_txpipe6_width                             (o_txpipe6_width),                                                                      //  output,    width = 3,                                       .o_txpipe6_width
		.o_pcs7_pipe_rst_n                           (o_pcs7_pipe_rst_n),                                                                    //  output,    width = 1,                                       .o_pcs7_pipe_rst_n
		.i_rxpipe7_dirfeedback                       (i_rxpipe7_dirfeedback),                                                                //   input,    width = 6,                                       .i_rxpipe7_dirfeedback
		.i_rxpipe7_linkevaluationfeedbackfiguremerit (i_rxpipe7_linkevaluationfeedbackfiguremerit),                                          //   input,    width = 8,                                       .i_rxpipe7_linkevaluationfeedbackfiguremerit
		.i_rxpipe7_localfs                           (i_rxpipe7_localfs),                                                                    //   input,    width = 6,                                       .i_rxpipe7_localfs
		.i_rxpipe7_locallf                           (i_rxpipe7_locallf),                                                                    //   input,    width = 6,                                       .i_rxpipe7_locallf
		.i_rxpipe7_localtxcoefficientsvalid          (i_rxpipe7_localtxcoefficientsvalid),                                                   //   input,    width = 1,                                       .i_rxpipe7_localtxcoefficientsvalid
		.i_rxpipe7_localtxpresetcoefficients         (i_rxpipe7_localtxpresetcoefficients),                                                  //   input,   width = 18,                                       .i_rxpipe7_localtxpresetcoefficients
		.i_rxpipe7_p2m_bus                           (i_rxpipe7_p2m_bus),                                                                    //   input,    width = 8,                                       .i_rxpipe7_p2m_bus
		.i_rxpipe7_pclkchangeok                      (i_rxpipe7_pclkchangeok),                                                               //   input,    width = 1,                                       .i_rxpipe7_pclkchangeok
		.i_rxpipe7_phystatus                         (i_rxpipe7_phystatus),                                                                  //   input,    width = 1,                                       .i_rxpipe7_phystatus
		.i_rxpipe7_rxdata                            (i_rxpipe7_rxdata),                                                                     //   input,   width = 40,                                       .i_rxpipe7_rxdata
		.i_rxpipe7_rxdatak                           (i_rxpipe7_rxdatak),                                                                    //   input,    width = 4,                                       .i_rxpipe7_rxdatak
		.i_rxpipe7_rxdatavalid                       (i_rxpipe7_rxdatavalid),                                                                //   input,    width = 1,                                       .i_rxpipe7_rxdatavalid
		.i_rxpipe7_rxelecidlea                       (i_rxpipe7_rxelecidlea),                                                                //   input,    width = 1,                                       .i_rxpipe7_rxelecidlea
		.i_rxpipe7_rxstandbystatus                   (i_rxpipe7_rxstandbystatus),                                                            //   input,    width = 1,                                       .i_rxpipe7_rxstandbystatus
		.i_rxpipe7_rxstartblock                      (i_rxpipe7_rxstartblock),                                                               //   input,    width = 1,                                       .i_rxpipe7_rxstartblock
		.i_rxpipe7_rxstatus                          (i_rxpipe7_rxstatus),                                                                   //   input,    width = 3,                                       .i_rxpipe7_rxstatus
		.i_rxpipe7_rxsyncheader                      (i_rxpipe7_rxsyncheader),                                                               //   input,    width = 4,                                       .i_rxpipe7_rxsyncheader
		.i_rxpipe7_rxvalid                           (i_rxpipe7_rxvalid),                                                                    //   input,    width = 1,                                       .i_rxpipe7_rxvalid
		.o_txpipe7_asyncpowerchangeack               (o_txpipe7_asyncpowerchangeack),                                                        //  output,    width = 1,                                       .o_txpipe7_asyncpowerchangeack
		.o_txpipe7_blockaligncontrol                 (o_txpipe7_blockaligncontrol),                                                          //  output,    width = 1,                                       .o_txpipe7_blockaligncontrol
		.o_txpipe7_cfg_hw_auto_sp_dis                (o_txpipe7_cfg_hw_auto_sp_dis),                                                         //  output,    width = 1,                                       .o_txpipe7_cfg_hw_auto_sp_dis
		.o_txpipe7_dirchange                         (o_txpipe7_dirchange),                                                                  //  output,    width = 1,                                       .o_txpipe7_dirchange
		.o_txpipe7_ebuf_mode                         (o_txpipe7_ebuf_mode),                                                                  //  output,    width = 1,                                       .o_txpipe7_ebuf_mode
		.o_txpipe7_encodedecodebypass                (o_txpipe7_encodedecodebypass),                                                         //  output,    width = 1,                                       .o_txpipe7_encodedecodebypass
		.o_txpipe7_fs                                (o_txpipe7_fs),                                                                         //  output,    width = 6,                                       .o_txpipe7_fs
		.o_txpipe7_getlocalpresetcoefficients        (o_txpipe7_getlocalpresetcoefficients),                                                 //  output,    width = 1,                                       .o_txpipe7_getlocalpresetcoefficients
		.o_txpipe7_invalidrequest                    (o_txpipe7_invalidrequest),                                                             //  output,    width = 1,                                       .o_txpipe7_invalidrequest
		.o_txpipe7_lf                                (o_txpipe7_lf),                                                                         //  output,    width = 6,                                       .o_txpipe7_lf
		.o_txpipe7_localpresetindex                  (o_txpipe7_localpresetindex),                                                           //  output,    width = 5,                                       .o_txpipe7_localpresetindex
		.o_txpipe7_lowpin_nt                         (o_txpipe7_lowpin_nt),                                                                  //  output,    width = 1,                                       .o_txpipe7_lowpin_nt
		.o_txpipe7_m2p_bus                           (o_txpipe7_m2p_bus),                                                                    //  output,    width = 8,                                       .o_txpipe7_m2p_bus
		.o_txpipe7_pclk_rate                         (o_txpipe7_pclk_rate),                                                                  //  output,    width = 3,                                       .o_txpipe7_pclk_rate
		.o_txpipe7_pclkchangeack                     (o_txpipe7_pclkchangeack),                                                              //  output,    width = 1,                                       .o_txpipe7_pclkchangeack
		.o_txpipe7_phy_mode_nt                       (o_txpipe7_phy_mode_nt),                                                                //  output,    width = 4,                                       .o_txpipe7_phy_mode_nt
		.o_txpipe7_powerdown                         (o_txpipe7_powerdown),                                                                  //  output,    width = 4,                                       .o_txpipe7_powerdown
		.o_txpipe7_rate                              (o_txpipe7_rate),                                                                       //  output,    width = 3,                                       .o_txpipe7_rate
		.o_txpipe7_rxelecidle_disable_a              (o_txpipe7_rxelecidle_disable_a),                                                       //  output,    width = 1,                                       .o_txpipe7_rxelecidle_disable_a
		.o_txpipe7_rxeqclr                           (o_txpipe7_rxeqclr),                                                                    //  output,    width = 1,                                       .o_txpipe7_rxeqclr
		.o_txpipe7_rxeqeval                          (o_txpipe7_rxeqeval),                                                                   //  output,    width = 1,                                       .o_txpipe7_rxeqeval
		.o_txpipe7_rxeqinprogress                    (o_txpipe7_rxeqinprogress),                                                             //  output,    width = 1,                                       .o_txpipe7_rxeqinprogress
		.o_txpipe7_rxeqtraining                      (o_txpipe7_rxeqtraining),                                                               //  output,    width = 1,                                       .o_txpipe7_rxeqtraining
		.o_txpipe7_rxpolarity                        (o_txpipe7_rxpolarity),                                                                 //  output,    width = 1,                                       .o_txpipe7_rxpolarity
		.o_txpipe7_rxpresethint                      (o_txpipe7_rxpresethint),                                                               //  output,    width = 3,                                       .o_txpipe7_rxpresethint
		.o_txpipe7_rxstandby                         (o_txpipe7_rxstandby),                                                                  //  output,    width = 1,                                       .o_txpipe7_rxstandby
		.o_txpipe7_rxtermination                     (o_txpipe7_rxtermination),                                                              //  output,    width = 1,                                       .o_txpipe7_rxtermination
		.o_txpipe7_srisenable                        (o_txpipe7_srisenable),                                                                 //  output,    width = 1,                                       .o_txpipe7_srisenable
		.o_txpipe7_txcmnmode_disable_a               (o_txpipe7_txcmnmode_disable_a),                                                        //  output,    width = 1,                                       .o_txpipe7_txcmnmode_disable_a
		.o_txpipe7_txcompliance                      (o_txpipe7_txcompliance),                                                               //  output,    width = 1,                                       .o_txpipe7_txcompliance
		.o_txpipe7_txdata                            (o_txpipe7_txdata),                                                                     //  output,   width = 40,                                       .o_txpipe7_txdata
		.o_txpipe7_txdatak                           (o_txpipe7_txdatak),                                                                    //  output,    width = 4,                                       .o_txpipe7_txdatak
		.o_txpipe7_txdatavalid                       (o_txpipe7_txdatavalid),                                                                //  output,    width = 1,                                       .o_txpipe7_txdatavalid
		.o_txpipe7_txdeemph                          (o_txpipe7_txdeemph),                                                                   //  output,   width = 18,                                       .o_txpipe7_txdeemph
		.o_txpipe7_txdtctrx_lb                       (o_txpipe7_txdtctrx_lb),                                                                //  output,    width = 1,                                       .o_txpipe7_txdtctrx_lb
		.o_txpipe7_txelecidle                        (o_txpipe7_txelecidle),                                                                 //  output,    width = 1,                                       .o_txpipe7_txelecidle
		.o_txpipe7_txmargin                          (o_txpipe7_txmargin),                                                                   //  output,    width = 3,                                       .o_txpipe7_txmargin
		.o_txpipe7_txoneszeros                       (o_txpipe7_txoneszeros),                                                                //  output,    width = 1,                                       .o_txpipe7_txoneszeros
		.o_txpipe7_txstartblock                      (o_txpipe7_txstartblock),                                                               //  output,    width = 1,                                       .o_txpipe7_txstartblock
		.o_txpipe7_txswing                           (o_txpipe7_txswing),                                                                    //  output,    width = 1,                                       .o_txpipe7_txswing
		.o_txpipe7_txsyncheader                      (o_txpipe7_txsyncheader),                                                               //  output,    width = 4,                                       .o_txpipe7_txsyncheader
		.o_txpipe7_width                             (o_txpipe7_width),                                                                      //  output,    width = 3,                                       .o_txpipe7_width
		.i_pin_perst_n                               (i_pin_perst_n),                                                                        //   input,    width = 1,                                       .i_pin_perst_n
		.i_hio_ch0_lavmm_clk                         (i_hio_ch0_lavmm_clk),                                                                  //   input,    width = 1,                    i_hio_ch0_lavmm_clk.clk
		.i_hio_ch0_lavmm_rstn                        (i_hio_ch0_lavmm_rstn),                                                                 //   input,    width = 1,                   i_hio_ch0_lavmm_rstn.reset
		.i_hio_ch0_lavmm_addr                        (i_hio_ch0_lavmm_addr),                                                                 //   input,   width = 21,                          hio_ch0_lavmm.address
		.i_hio_ch0_lavmm_be                          (i_hio_ch0_lavmm_be),                                                                   //   input,    width = 4,                                       .byteenable
		.o_hio_ch0_lavmm_rdata_valid                 (o_hio_ch0_lavmm_rdata_valid),                                                          //  output,    width = 1,                                       .readdatavalid
		.i_hio_ch0_lavmm_read                        (i_hio_ch0_lavmm_read),                                                                 //   input,    width = 1,                                       .read
		.i_hio_ch0_lavmm_write                       (i_hio_ch0_lavmm_write),                                                                //   input,    width = 1,                                       .write
		.o_hio_ch0_lavmm_rdata                       (o_hio_ch0_lavmm_rdata),                                                                //  output,   width = 32,                                       .readdata
		.i_hio_ch0_lavmm_wdata                       (i_hio_ch0_lavmm_wdata),                                                                //   input,   width = 32,                                       .writedata
		.o_hio_ch0_lavmm_waitreq                     (o_hio_ch0_lavmm_waitreq),                                                              //  output,    width = 1,                                       .waitrequest
		.i_hio_ch0_pld_rx_clk_in_row_clk             (i_hio_ch0_pld_rx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch0_pld_rx_clk_in_row_clk.clk
		.i_hio_ch0_pld_tx_clk_in_row_clk             (i_hio_ch0_pld_tx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch0_pld_tx_clk_in_row_clk.clk
		.i_hio_ch0_det_lat_rx_dl_clk                 (i_hio_ch0_det_lat_rx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch0_det_lat_rx_dl_clk.clk
		.i_hio_ch0_det_lat_rx_mux_select             (i_hio_ch0_det_lat_rx_mux_select),                                                      //   input,    width = 1,        i_hio_ch0_det_lat_rx_mux_select.clk
		.i_hio_ch0_det_lat_rx_sclk_flop              (i_hio_ch0_det_lat_rx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch0_det_lat_rx_sclk_flop.clk
		.i_hio_ch0_det_lat_rx_sclk_gen_clk           (i_hio_ch0_det_lat_rx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch0_det_lat_rx_sclk_gen_clk.clk
		.i_hio_ch0_det_lat_rx_trig_flop              (i_hio_ch0_det_lat_rx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch0_det_lat_rx_trig_flop.clk
		.i_hio_ch0_det_lat_sampling_clk              (i_hio_ch0_det_lat_sampling_clk),                                                       //   input,    width = 1,         i_hio_ch0_det_lat_sampling_clk.clk
		.i_hio_ch0_det_lat_tx_dl_clk                 (i_hio_ch0_det_lat_tx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch0_det_lat_tx_dl_clk.clk
		.i_hio_ch0_det_lat_tx_mux_select             (i_hio_ch0_det_lat_tx_mux_select),                                                      //   input,    width = 1,        i_hio_ch0_det_lat_tx_mux_select.clk
		.i_hio_ch0_det_lat_tx_sclk_flop              (i_hio_ch0_det_lat_tx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch0_det_lat_tx_sclk_flop.clk
		.i_hio_ch0_det_lat_tx_sclk_gen_clk           (i_hio_ch0_det_lat_tx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch0_det_lat_tx_sclk_gen_clk.clk
		.i_hio_ch0_det_lat_tx_trig_flop              (i_hio_ch0_det_lat_tx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch0_det_lat_tx_trig_flop.clk
		.o_hio_ch0_user_rx_clk1_clk                  (o_hio_ch0_user_rx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch0_user_rx_clk1_clk.clk
		.o_hio_ch0_user_rx_clk2_clk                  (o_hio_ch0_user_rx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch0_user_rx_clk2_clk.clk
		.o_hio_ch0_user_tx_clk1_clk                  (o_hio_ch0_user_tx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch0_user_tx_clk1_clk.clk
		.o_hio_ch0_user_tx_clk2_clk                  (o_hio_ch0_user_tx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch0_user_tx_clk2_clk.clk
		.o_hio_ch0_ux_chnl_refclk_mux                (o_hio_ch0_ux_chnl_refclk_mux),                                                         //  output,    width = 1,           o_hio_ch0_ux_chnl_refclk_mux.clk
		.o_hio_ch0_det_lat_rx_async_dl_sync          (o_hio_ch0_det_lat_rx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch0_det_lat_rx_async_dl_sync.clk
		.o_hio_ch0_det_lat_rx_async_pulse            (o_hio_ch0_det_lat_rx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch0_det_lat_rx_async_pulse.clk
		.o_hio_ch0_det_lat_rx_async_sample_sync      (o_hio_ch0_det_lat_rx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch0_det_lat_rx_async_sample_sync.clk
		.o_hio_ch0_det_lat_rx_sclk_sample_sync       (o_hio_ch0_det_lat_rx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch0_det_lat_rx_sclk_sample_sync.clk
		.o_hio_ch0_det_lat_rx_trig_sample_sync       (o_hio_ch0_det_lat_rx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch0_det_lat_rx_trig_sample_sync.clk
		.o_hio_ch0_det_lat_tx_async_dl_sync          (o_hio_ch0_det_lat_tx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch0_det_lat_tx_async_dl_sync.clk
		.o_hio_ch0_det_lat_tx_async_pulse            (o_hio_ch0_det_lat_tx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch0_det_lat_tx_async_pulse.clk
		.o_hio_ch0_det_lat_tx_async_sample_sync      (o_hio_ch0_det_lat_tx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch0_det_lat_tx_async_sample_sync.clk
		.o_hio_ch0_det_lat_tx_sclk_sample_sync       (o_hio_ch0_det_lat_tx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch0_det_lat_tx_sclk_sample_sync.clk
		.o_hio_ch0_det_lat_tx_trig_sample_sync       (o_hio_ch0_det_lat_tx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch0_det_lat_tx_trig_sample_sync.clk
		.o_hio_ch0_xcvrif_rx_latency_pulse           (o_hio_ch0_xcvrif_rx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch0_xcvrif_rx_latency_pulse.clk
		.o_hio_ch0_xcvrif_tx_latency_pulse           (o_hio_ch0_xcvrif_tx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch0_xcvrif_tx_latency_pulse.clk
		.i_hio_ch1_lavmm_clk                         (i_hio_ch1_lavmm_clk),                                                                  //   input,    width = 1,                    i_hio_ch1_lavmm_clk.clk
		.i_hio_ch1_lavmm_rstn                        (i_hio_ch1_lavmm_rstn),                                                                 //   input,    width = 1,                   i_hio_ch1_lavmm_rstn.reset
		.i_hio_ch1_lavmm_addr                        (i_hio_ch1_lavmm_addr),                                                                 //   input,   width = 21,                          hio_ch1_lavmm.address
		.i_hio_ch1_lavmm_be                          (i_hio_ch1_lavmm_be),                                                                   //   input,    width = 4,                                       .byteenable
		.o_hio_ch1_lavmm_rdata_valid                 (o_hio_ch1_lavmm_rdata_valid),                                                          //  output,    width = 1,                                       .readdatavalid
		.i_hio_ch1_lavmm_read                        (i_hio_ch1_lavmm_read),                                                                 //   input,    width = 1,                                       .read
		.i_hio_ch1_lavmm_write                       (i_hio_ch1_lavmm_write),                                                                //   input,    width = 1,                                       .write
		.o_hio_ch1_lavmm_rdata                       (o_hio_ch1_lavmm_rdata),                                                                //  output,   width = 32,                                       .readdata
		.i_hio_ch1_lavmm_wdata                       (i_hio_ch1_lavmm_wdata),                                                                //   input,   width = 32,                                       .writedata
		.o_hio_ch1_lavmm_waitreq                     (o_hio_ch1_lavmm_waitreq),                                                              //  output,    width = 1,                                       .waitrequest
		.i_hio_ch1_pld_rx_clk_in_row_clk             (i_hio_ch1_pld_rx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch1_pld_rx_clk_in_row_clk.clk
		.i_hio_ch1_pld_tx_clk_in_row_clk             (i_hio_ch1_pld_tx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch1_pld_tx_clk_in_row_clk.clk
		.i_hio_ch1_det_lat_rx_dl_clk                 (i_hio_ch1_det_lat_rx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch1_det_lat_rx_dl_clk.clk
		.i_hio_ch1_det_lat_rx_mux_select             (i_hio_ch1_det_lat_rx_mux_select),                                                      //   input,    width = 1,        i_hio_ch1_det_lat_rx_mux_select.clk
		.i_hio_ch1_det_lat_rx_sclk_flop              (i_hio_ch1_det_lat_rx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch1_det_lat_rx_sclk_flop.clk
		.i_hio_ch1_det_lat_rx_sclk_gen_clk           (i_hio_ch1_det_lat_rx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch1_det_lat_rx_sclk_gen_clk.clk
		.i_hio_ch1_det_lat_rx_trig_flop              (i_hio_ch1_det_lat_rx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch1_det_lat_rx_trig_flop.clk
		.i_hio_ch1_det_lat_sampling_clk              (i_hio_ch1_det_lat_sampling_clk),                                                       //   input,    width = 1,         i_hio_ch1_det_lat_sampling_clk.clk
		.i_hio_ch1_det_lat_tx_dl_clk                 (i_hio_ch1_det_lat_tx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch1_det_lat_tx_dl_clk.clk
		.i_hio_ch1_det_lat_tx_mux_select             (i_hio_ch1_det_lat_tx_mux_select),                                                      //   input,    width = 1,        i_hio_ch1_det_lat_tx_mux_select.clk
		.i_hio_ch1_det_lat_tx_sclk_flop              (i_hio_ch1_det_lat_tx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch1_det_lat_tx_sclk_flop.clk
		.i_hio_ch1_det_lat_tx_sclk_gen_clk           (i_hio_ch1_det_lat_tx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch1_det_lat_tx_sclk_gen_clk.clk
		.i_hio_ch1_det_lat_tx_trig_flop              (i_hio_ch1_det_lat_tx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch1_det_lat_tx_trig_flop.clk
		.o_hio_ch1_user_rx_clk1_clk                  (o_hio_ch1_user_rx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch1_user_rx_clk1_clk.clk
		.o_hio_ch1_user_rx_clk2_clk                  (o_hio_ch1_user_rx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch1_user_rx_clk2_clk.clk
		.o_hio_ch1_user_tx_clk1_clk                  (o_hio_ch1_user_tx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch1_user_tx_clk1_clk.clk
		.o_hio_ch1_user_tx_clk2_clk                  (o_hio_ch1_user_tx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch1_user_tx_clk2_clk.clk
		.o_hio_ch1_ux_chnl_refclk_mux                (o_hio_ch1_ux_chnl_refclk_mux),                                                         //  output,    width = 1,           o_hio_ch1_ux_chnl_refclk_mux.clk
		.o_hio_ch1_det_lat_rx_async_dl_sync          (o_hio_ch1_det_lat_rx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch1_det_lat_rx_async_dl_sync.clk
		.o_hio_ch1_det_lat_rx_async_pulse            (o_hio_ch1_det_lat_rx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch1_det_lat_rx_async_pulse.clk
		.o_hio_ch1_det_lat_rx_async_sample_sync      (o_hio_ch1_det_lat_rx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch1_det_lat_rx_async_sample_sync.clk
		.o_hio_ch1_det_lat_rx_sclk_sample_sync       (o_hio_ch1_det_lat_rx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch1_det_lat_rx_sclk_sample_sync.clk
		.o_hio_ch1_det_lat_rx_trig_sample_sync       (o_hio_ch1_det_lat_rx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch1_det_lat_rx_trig_sample_sync.clk
		.o_hio_ch1_det_lat_tx_async_dl_sync          (o_hio_ch1_det_lat_tx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch1_det_lat_tx_async_dl_sync.clk
		.o_hio_ch1_det_lat_tx_async_pulse            (o_hio_ch1_det_lat_tx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch1_det_lat_tx_async_pulse.clk
		.o_hio_ch1_det_lat_tx_async_sample_sync      (o_hio_ch1_det_lat_tx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch1_det_lat_tx_async_sample_sync.clk
		.o_hio_ch1_det_lat_tx_sclk_sample_sync       (o_hio_ch1_det_lat_tx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch1_det_lat_tx_sclk_sample_sync.clk
		.o_hio_ch1_det_lat_tx_trig_sample_sync       (o_hio_ch1_det_lat_tx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch1_det_lat_tx_trig_sample_sync.clk
		.o_hio_ch1_xcvrif_rx_latency_pulse           (o_hio_ch1_xcvrif_rx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch1_xcvrif_rx_latency_pulse.clk
		.o_hio_ch1_xcvrif_tx_latency_pulse           (o_hio_ch1_xcvrif_tx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch1_xcvrif_tx_latency_pulse.clk
		.i_hio_ch2_lavmm_clk                         (i_hio_ch2_lavmm_clk),                                                                  //   input,    width = 1,                    i_hio_ch2_lavmm_clk.clk
		.i_hio_ch2_lavmm_rstn                        (i_hio_ch2_lavmm_rstn),                                                                 //   input,    width = 1,                   i_hio_ch2_lavmm_rstn.reset
		.i_hio_ch2_lavmm_addr                        (i_hio_ch2_lavmm_addr),                                                                 //   input,   width = 21,                          hio_ch2_lavmm.address
		.i_hio_ch2_lavmm_be                          (i_hio_ch2_lavmm_be),                                                                   //   input,    width = 4,                                       .byteenable
		.o_hio_ch2_lavmm_rdata_valid                 (o_hio_ch2_lavmm_rdata_valid),                                                          //  output,    width = 1,                                       .readdatavalid
		.i_hio_ch2_lavmm_read                        (i_hio_ch2_lavmm_read),                                                                 //   input,    width = 1,                                       .read
		.i_hio_ch2_lavmm_write                       (i_hio_ch2_lavmm_write),                                                                //   input,    width = 1,                                       .write
		.o_hio_ch2_lavmm_rdata                       (o_hio_ch2_lavmm_rdata),                                                                //  output,   width = 32,                                       .readdata
		.i_hio_ch2_lavmm_wdata                       (i_hio_ch2_lavmm_wdata),                                                                //   input,   width = 32,                                       .writedata
		.o_hio_ch2_lavmm_waitreq                     (o_hio_ch2_lavmm_waitreq),                                                              //  output,    width = 1,                                       .waitrequest
		.i_hio_ch2_pld_rx_clk_in_row_clk             (i_hio_ch2_pld_rx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch2_pld_rx_clk_in_row_clk.clk
		.i_hio_ch2_pld_tx_clk_in_row_clk             (i_hio_ch2_pld_tx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch2_pld_tx_clk_in_row_clk.clk
		.i_hio_ch2_det_lat_rx_dl_clk                 (i_hio_ch2_det_lat_rx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch2_det_lat_rx_dl_clk.clk
		.i_hio_ch2_det_lat_rx_mux_select             (i_hio_ch2_det_lat_rx_mux_select),                                                      //   input,    width = 1,        i_hio_ch2_det_lat_rx_mux_select.clk
		.i_hio_ch2_det_lat_rx_sclk_flop              (i_hio_ch2_det_lat_rx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch2_det_lat_rx_sclk_flop.clk
		.i_hio_ch2_det_lat_rx_sclk_gen_clk           (i_hio_ch2_det_lat_rx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch2_det_lat_rx_sclk_gen_clk.clk
		.i_hio_ch2_det_lat_rx_trig_flop              (i_hio_ch2_det_lat_rx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch2_det_lat_rx_trig_flop.clk
		.i_hio_ch2_det_lat_sampling_clk              (i_hio_ch2_det_lat_sampling_clk),                                                       //   input,    width = 1,         i_hio_ch2_det_lat_sampling_clk.clk
		.i_hio_ch2_det_lat_tx_dl_clk                 (i_hio_ch2_det_lat_tx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch2_det_lat_tx_dl_clk.clk
		.i_hio_ch2_det_lat_tx_mux_select             (i_hio_ch2_det_lat_tx_mux_select),                                                      //   input,    width = 1,        i_hio_ch2_det_lat_tx_mux_select.clk
		.i_hio_ch2_det_lat_tx_sclk_flop              (i_hio_ch2_det_lat_tx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch2_det_lat_tx_sclk_flop.clk
		.i_hio_ch2_det_lat_tx_sclk_gen_clk           (i_hio_ch2_det_lat_tx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch2_det_lat_tx_sclk_gen_clk.clk
		.i_hio_ch2_det_lat_tx_trig_flop              (i_hio_ch2_det_lat_tx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch2_det_lat_tx_trig_flop.clk
		.o_hio_ch2_user_rx_clk1_clk                  (o_hio_ch2_user_rx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch2_user_rx_clk1_clk.clk
		.o_hio_ch2_user_rx_clk2_clk                  (o_hio_ch2_user_rx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch2_user_rx_clk2_clk.clk
		.o_hio_ch2_user_tx_clk1_clk                  (o_hio_ch2_user_tx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch2_user_tx_clk1_clk.clk
		.o_hio_ch2_user_tx_clk2_clk                  (o_hio_ch2_user_tx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch2_user_tx_clk2_clk.clk
		.o_hio_ch2_ux_chnl_refclk_mux                (o_hio_ch2_ux_chnl_refclk_mux),                                                         //  output,    width = 1,           o_hio_ch2_ux_chnl_refclk_mux.clk
		.o_hio_ch2_det_lat_rx_async_dl_sync          (o_hio_ch2_det_lat_rx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch2_det_lat_rx_async_dl_sync.clk
		.o_hio_ch2_det_lat_rx_async_pulse            (o_hio_ch2_det_lat_rx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch2_det_lat_rx_async_pulse.clk
		.o_hio_ch2_det_lat_rx_async_sample_sync      (o_hio_ch2_det_lat_rx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch2_det_lat_rx_async_sample_sync.clk
		.o_hio_ch2_det_lat_rx_sclk_sample_sync       (o_hio_ch2_det_lat_rx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch2_det_lat_rx_sclk_sample_sync.clk
		.o_hio_ch2_det_lat_rx_trig_sample_sync       (o_hio_ch2_det_lat_rx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch2_det_lat_rx_trig_sample_sync.clk
		.o_hio_ch2_det_lat_tx_async_dl_sync          (o_hio_ch2_det_lat_tx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch2_det_lat_tx_async_dl_sync.clk
		.o_hio_ch2_det_lat_tx_async_pulse            (o_hio_ch2_det_lat_tx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch2_det_lat_tx_async_pulse.clk
		.o_hio_ch2_det_lat_tx_async_sample_sync      (o_hio_ch2_det_lat_tx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch2_det_lat_tx_async_sample_sync.clk
		.o_hio_ch2_det_lat_tx_sclk_sample_sync       (o_hio_ch2_det_lat_tx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch2_det_lat_tx_sclk_sample_sync.clk
		.o_hio_ch2_det_lat_tx_trig_sample_sync       (o_hio_ch2_det_lat_tx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch2_det_lat_tx_trig_sample_sync.clk
		.o_hio_ch2_xcvrif_rx_latency_pulse           (o_hio_ch2_xcvrif_rx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch2_xcvrif_rx_latency_pulse.clk
		.o_hio_ch2_xcvrif_tx_latency_pulse           (o_hio_ch2_xcvrif_tx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch2_xcvrif_tx_latency_pulse.clk
		.i_hio_ch3_lavmm_clk                         (i_hio_ch3_lavmm_clk),                                                                  //   input,    width = 1,                    i_hio_ch3_lavmm_clk.clk
		.i_hio_ch3_lavmm_rstn                        (i_hio_ch3_lavmm_rstn),                                                                 //   input,    width = 1,                   i_hio_ch3_lavmm_rstn.reset
		.i_hio_ch3_lavmm_addr                        (i_hio_ch3_lavmm_addr),                                                                 //   input,   width = 21,                          hio_ch3_lavmm.address
		.i_hio_ch3_lavmm_be                          (i_hio_ch3_lavmm_be),                                                                   //   input,    width = 4,                                       .byteenable
		.o_hio_ch3_lavmm_rdata_valid                 (o_hio_ch3_lavmm_rdata_valid),                                                          //  output,    width = 1,                                       .readdatavalid
		.i_hio_ch3_lavmm_read                        (i_hio_ch3_lavmm_read),                                                                 //   input,    width = 1,                                       .read
		.i_hio_ch3_lavmm_write                       (i_hio_ch3_lavmm_write),                                                                //   input,    width = 1,                                       .write
		.o_hio_ch3_lavmm_rdata                       (o_hio_ch3_lavmm_rdata),                                                                //  output,   width = 32,                                       .readdata
		.i_hio_ch3_lavmm_wdata                       (i_hio_ch3_lavmm_wdata),                                                                //   input,   width = 32,                                       .writedata
		.o_hio_ch3_lavmm_waitreq                     (o_hio_ch3_lavmm_waitreq),                                                              //  output,    width = 1,                                       .waitrequest
		.i_hio_ch3_pld_rx_clk_in_row_clk             (i_hio_ch3_pld_rx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch3_pld_rx_clk_in_row_clk.clk
		.i_hio_ch3_pld_tx_clk_in_row_clk             (i_hio_ch3_pld_tx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch3_pld_tx_clk_in_row_clk.clk
		.i_hio_ch3_det_lat_rx_dl_clk                 (i_hio_ch3_det_lat_rx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch3_det_lat_rx_dl_clk.clk
		.i_hio_ch3_det_lat_rx_mux_select             (i_hio_ch3_det_lat_rx_mux_select),                                                      //   input,    width = 1,        i_hio_ch3_det_lat_rx_mux_select.clk
		.i_hio_ch3_det_lat_rx_sclk_flop              (i_hio_ch3_det_lat_rx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch3_det_lat_rx_sclk_flop.clk
		.i_hio_ch3_det_lat_rx_sclk_gen_clk           (i_hio_ch3_det_lat_rx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch3_det_lat_rx_sclk_gen_clk.clk
		.i_hio_ch3_det_lat_rx_trig_flop              (i_hio_ch3_det_lat_rx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch3_det_lat_rx_trig_flop.clk
		.i_hio_ch3_det_lat_sampling_clk              (i_hio_ch3_det_lat_sampling_clk),                                                       //   input,    width = 1,         i_hio_ch3_det_lat_sampling_clk.clk
		.i_hio_ch3_det_lat_tx_dl_clk                 (i_hio_ch3_det_lat_tx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch3_det_lat_tx_dl_clk.clk
		.i_hio_ch3_det_lat_tx_mux_select             (i_hio_ch3_det_lat_tx_mux_select),                                                      //   input,    width = 1,        i_hio_ch3_det_lat_tx_mux_select.clk
		.i_hio_ch3_det_lat_tx_sclk_flop              (i_hio_ch3_det_lat_tx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch3_det_lat_tx_sclk_flop.clk
		.i_hio_ch3_det_lat_tx_sclk_gen_clk           (i_hio_ch3_det_lat_tx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch3_det_lat_tx_sclk_gen_clk.clk
		.i_hio_ch3_det_lat_tx_trig_flop              (i_hio_ch3_det_lat_tx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch3_det_lat_tx_trig_flop.clk
		.o_hio_ch3_user_rx_clk1_clk                  (o_hio_ch3_user_rx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch3_user_rx_clk1_clk.clk
		.o_hio_ch3_user_rx_clk2_clk                  (o_hio_ch3_user_rx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch3_user_rx_clk2_clk.clk
		.o_hio_ch3_user_tx_clk1_clk                  (o_hio_ch3_user_tx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch3_user_tx_clk1_clk.clk
		.o_hio_ch3_user_tx_clk2_clk                  (o_hio_ch3_user_tx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch3_user_tx_clk2_clk.clk
		.o_hio_ch3_ux_chnl_refclk_mux                (o_hio_ch3_ux_chnl_refclk_mux),                                                         //  output,    width = 1,           o_hio_ch3_ux_chnl_refclk_mux.clk
		.o_hio_ch3_det_lat_rx_async_dl_sync          (o_hio_ch3_det_lat_rx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch3_det_lat_rx_async_dl_sync.clk
		.o_hio_ch3_det_lat_rx_async_pulse            (o_hio_ch3_det_lat_rx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch3_det_lat_rx_async_pulse.clk
		.o_hio_ch3_det_lat_rx_async_sample_sync      (o_hio_ch3_det_lat_rx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch3_det_lat_rx_async_sample_sync.clk
		.o_hio_ch3_det_lat_rx_sclk_sample_sync       (o_hio_ch3_det_lat_rx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch3_det_lat_rx_sclk_sample_sync.clk
		.o_hio_ch3_det_lat_rx_trig_sample_sync       (o_hio_ch3_det_lat_rx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch3_det_lat_rx_trig_sample_sync.clk
		.o_hio_ch3_det_lat_tx_async_dl_sync          (o_hio_ch3_det_lat_tx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch3_det_lat_tx_async_dl_sync.clk
		.o_hio_ch3_det_lat_tx_async_pulse            (o_hio_ch3_det_lat_tx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch3_det_lat_tx_async_pulse.clk
		.o_hio_ch3_det_lat_tx_async_sample_sync      (o_hio_ch3_det_lat_tx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch3_det_lat_tx_async_sample_sync.clk
		.o_hio_ch3_det_lat_tx_sclk_sample_sync       (o_hio_ch3_det_lat_tx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch3_det_lat_tx_sclk_sample_sync.clk
		.o_hio_ch3_det_lat_tx_trig_sample_sync       (o_hio_ch3_det_lat_tx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch3_det_lat_tx_trig_sample_sync.clk
		.o_hio_ch3_xcvrif_rx_latency_pulse           (o_hio_ch3_xcvrif_rx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch3_xcvrif_rx_latency_pulse.clk
		.o_hio_ch3_xcvrif_tx_latency_pulse           (o_hio_ch3_xcvrif_tx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch3_xcvrif_tx_latency_pulse.clk
		.i_hio_ch4_lavmm_clk                         (i_hio_ch4_lavmm_clk),                                                                  //   input,    width = 1,                    i_hio_ch4_lavmm_clk.clk
		.i_hio_ch4_lavmm_rstn                        (i_hio_ch4_lavmm_rstn),                                                                 //   input,    width = 1,                   i_hio_ch4_lavmm_rstn.reset
		.i_hio_ch4_lavmm_addr                        (i_hio_ch4_lavmm_addr),                                                                 //   input,   width = 21,                          hio_ch4_lavmm.address
		.i_hio_ch4_lavmm_be                          (i_hio_ch4_lavmm_be),                                                                   //   input,    width = 4,                                       .byteenable
		.o_hio_ch4_lavmm_rdata_valid                 (o_hio_ch4_lavmm_rdata_valid),                                                          //  output,    width = 1,                                       .readdatavalid
		.i_hio_ch4_lavmm_read                        (i_hio_ch4_lavmm_read),                                                                 //   input,    width = 1,                                       .read
		.i_hio_ch4_lavmm_write                       (i_hio_ch4_lavmm_write),                                                                //   input,    width = 1,                                       .write
		.o_hio_ch4_lavmm_rdata                       (o_hio_ch4_lavmm_rdata),                                                                //  output,   width = 32,                                       .readdata
		.i_hio_ch4_lavmm_wdata                       (i_hio_ch4_lavmm_wdata),                                                                //   input,   width = 32,                                       .writedata
		.o_hio_ch4_lavmm_waitreq                     (o_hio_ch4_lavmm_waitreq),                                                              //  output,    width = 1,                                       .waitrequest
		.i_hio_ch4_pld_rx_clk_in_row_clk             (i_hio_ch4_pld_rx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch4_pld_rx_clk_in_row_clk.clk
		.i_hio_ch4_pld_tx_clk_in_row_clk             (i_hio_ch4_pld_tx_clk_in_row_clk),                                                      //   input,    width = 1,        i_hio_ch4_pld_tx_clk_in_row_clk.clk
		.i_hio_ch4_det_lat_rx_dl_clk                 (i_hio_ch4_det_lat_rx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch4_det_lat_rx_dl_clk.clk
		.i_hio_ch4_det_lat_rx_mux_select             (i_hio_ch4_det_lat_rx_mux_select),                                                      //   input,    width = 1,        i_hio_ch4_det_lat_rx_mux_select.clk
		.i_hio_ch4_det_lat_rx_sclk_flop              (i_hio_ch4_det_lat_rx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch4_det_lat_rx_sclk_flop.clk
		.i_hio_ch4_det_lat_rx_sclk_gen_clk           (i_hio_ch4_det_lat_rx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch4_det_lat_rx_sclk_gen_clk.clk
		.i_hio_ch4_det_lat_rx_trig_flop              (i_hio_ch4_det_lat_rx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch4_det_lat_rx_trig_flop.clk
		.i_hio_ch4_det_lat_sampling_clk              (i_hio_ch4_det_lat_sampling_clk),                                                       //   input,    width = 1,         i_hio_ch4_det_lat_sampling_clk.clk
		.i_hio_ch4_det_lat_tx_dl_clk                 (i_hio_ch4_det_lat_tx_dl_clk),                                                          //   input,    width = 1,            i_hio_ch4_det_lat_tx_dl_clk.clk
		.i_hio_ch4_det_lat_tx_mux_select             (i_hio_ch4_det_lat_tx_mux_select),                                                      //   input,    width = 1,        i_hio_ch4_det_lat_tx_mux_select.clk
		.i_hio_ch4_det_lat_tx_sclk_flop              (i_hio_ch4_det_lat_tx_sclk_flop),                                                       //   input,    width = 1,         i_hio_ch4_det_lat_tx_sclk_flop.clk
		.i_hio_ch4_det_lat_tx_sclk_gen_clk           (i_hio_ch4_det_lat_tx_sclk_gen_clk),                                                    //   input,    width = 1,      i_hio_ch4_det_lat_tx_sclk_gen_clk.clk
		.i_hio_ch4_det_lat_tx_trig_flop              (i_hio_ch4_det_lat_tx_trig_flop),                                                       //   input,    width = 1,         i_hio_ch4_det_lat_tx_trig_flop.clk
		.o_hio_ch4_user_rx_clk1_clk                  (o_hio_ch4_user_rx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch4_user_rx_clk1_clk.clk
		.o_hio_ch4_user_rx_clk2_clk                  (o_hio_ch4_user_rx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch4_user_rx_clk2_clk.clk
		.o_hio_ch4_user_tx_clk1_clk                  (o_hio_ch4_user_tx_clk1_clk),                                                           //  output,    width = 1,             o_hio_ch4_user_tx_clk1_clk.clk
		.o_hio_ch4_user_tx_clk2_clk                  (o_hio_ch4_user_tx_clk2_clk),                                                           //  output,    width = 1,             o_hio_ch4_user_tx_clk2_clk.clk
		.o_hio_ch4_ux_chnl_refclk_mux                (o_hio_ch4_ux_chnl_refclk_mux),                                                         //  output,    width = 1,           o_hio_ch4_ux_chnl_refclk_mux.clk
		.o_hio_ch4_det_lat_rx_async_dl_sync          (o_hio_ch4_det_lat_rx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch4_det_lat_rx_async_dl_sync.clk
		.o_hio_ch4_det_lat_rx_async_pulse            (o_hio_ch4_det_lat_rx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch4_det_lat_rx_async_pulse.clk
		.o_hio_ch4_det_lat_rx_async_sample_sync      (o_hio_ch4_det_lat_rx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch4_det_lat_rx_async_sample_sync.clk
		.o_hio_ch4_det_lat_rx_sclk_sample_sync       (o_hio_ch4_det_lat_rx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch4_det_lat_rx_sclk_sample_sync.clk
		.o_hio_ch4_det_lat_rx_trig_sample_sync       (o_hio_ch4_det_lat_rx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch4_det_lat_rx_trig_sample_sync.clk
		.o_hio_ch4_det_lat_tx_async_dl_sync          (o_hio_ch4_det_lat_tx_async_dl_sync),                                                   //  output,    width = 1,     o_hio_ch4_det_lat_tx_async_dl_sync.clk
		.o_hio_ch4_det_lat_tx_async_pulse            (o_hio_ch4_det_lat_tx_async_pulse),                                                     //  output,    width = 1,       o_hio_ch4_det_lat_tx_async_pulse.clk
		.o_hio_ch4_det_lat_tx_async_sample_sync      (o_hio_ch4_det_lat_tx_async_sample_sync),                                               //  output,    width = 1, o_hio_ch4_det_lat_tx_async_sample_sync.clk
		.o_hio_ch4_det_lat_tx_sclk_sample_sync       (o_hio_ch4_det_lat_tx_sclk_sample_sync),                                                //  output,    width = 1,  o_hio_ch4_det_lat_tx_sclk_sample_sync.clk
		.o_hio_ch4_det_lat_tx_trig_sample_sync       (o_hio_ch4_det_lat_tx_trig_sample_sync),                                                //  output,    width = 1,  o_hio_ch4_det_lat_tx_trig_sample_sync.clk
		.o_hio_ch4_xcvrif_rx_latency_pulse           (o_hio_ch4_xcvrif_rx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch4_xcvrif_rx_latency_pulse.clk
		.o_hio_ch4_xcvrif_tx_latency_pulse           (o_hio_ch4_xcvrif_tx_latency_pulse),                                                    //  output,    width = 1,      o_hio_ch4_xcvrif_tx_latency_pulse.clk
		.i_ch5_tx_data                               (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                                      
		.i_ch6_tx_data                               (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                                      
		.i_ch7_tx_data                               (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                                      
		.i_ch8_tx_data                               (80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                                      
		.o_ch5_rx_data                               (),                                                                                     // (terminated),                                                      
		.o_ch6_rx_data                               (),                                                                                     // (terminated),                                                      
		.o_ch7_rx_data                               (),                                                                                     // (terminated),                                                      
		.o_ch8_rx_data                               ()                                                                                      // (terminated),                                                      
	);

endmodule
