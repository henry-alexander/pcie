//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ors+7tAvFPlva1iUO2arrnEH/zOFS9iWvAJgOSc3r4d/71pnnDDVjIC2B3Co
Fxvt0IikT18F/BgjIK6JHv7xgsaaMb1rfs++YBVoPAUvsHFqxk3xN8GQuHTP
UbZlr0ERQ22ZJGs7KLt0keG/D3OzESf5B9+29DJ8oxD1NQqK9hpGioBKYdX7
UIDd2yXFmSBGQZuoBsW4fGWDSmYs3p+bVc+XbncDPoi6SP4aqQEv8MLszHEE
1QUENUfeHmz6eJmGKmc5PvUOYXAf1yP7EocWU/3dQL5wMTbL7i0+imjN9spj
PKyL+S0EiaYw87ZO9v5xvN964N10Pr0g7NMTNqgEQw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c9qGgbgt3/buF1Q+XNsnTWTytEgc4dz7cDvHDr0Y/9PEkjw+UOaW6UrKghk/
GpBZLthCbBcYq9xxI1Ecbi0vBwbw8wqzQVVvwTIA2pc/9WrcH7PyGWO+AMp8
AThAZYv5ePp55LVcTplvYNJuypty9BvUDgad0QG0B8btOqd+gA0zauzoG7YA
N9rxjMjbTq86xr1+a7o9rkcHiqEX6QL/mUFqtEokbm/JYl04Hf/Nhvmg3yz7
xviSjlcK+bgqAT9HwfHjs/fWVmEIbRi5qBG0h5HDzKUnorM/O9qI08b8RNTh
BgQ/PCnBBBuueKY1wjtmvVMlOiJClJGO9puM8qjpzQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Dg6op5zk8n+HkcYRiooIu2Uq7U8Tq7eoPLdeZjGAklZTHe0brqpkrDu8PKZu
ZqxZQ2e6bca+HmRNQtYBC37gqo6PcKsMGxmtjUIufZKwgBf6OQBk9UM8P/qy
eZFtNVVw99VOlyCHuC32SrHUnrMmRT+b81vPWeEAuf+9gAboCkc1u1oByQl8
mSZCsx5Ni+KxCWcquBGcO8cSo5a+XOPDaf11qUtKjBAzSV3EHad7i5DZY+J1
/wvVMn42yzpCrrK0wMjGIvrzuYUgWo03hitlQe8QpIOWZjxTPVZMBSyImqes
vBetH9IQHVl7xsRg3ZvGCKuvv4neEXJyJlAVTT5xQw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Kp0r68vYbg+RT2eyVQR7VQoM4Y+YCBvnNlc1JwHQzVZ0QWVS8q2ICLZIHil3
gzq8Kde+tWSdxwvtAMZszHKD+++02QhLwx664f7RnE10LcLIpRNjJL5GI3j1
bNU9njCwtDEiorY1lE9wGmpEUgQjLhnYOiB3XLZOUT+axecYTCE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
mFHd/fuJmptkgZTtIE4Kj9a4OXrHd6yukWSgd0skbz0ftAqOrXsbO8ibN7jG
RfLr+2u8K831/8vy84h7e20OCJgXFc0mYvWdycrLb97S+Ph7mJyZU/8Zeenc
1XdW+WGssUDEhv4SIUPXrauIbsWygXNxD7fXHrijZUnjYUujIpuZx/pK50Pi
gIlRSL7zxHUI81FLe+uVMudAIxSkDP/bclILhokB9knWYhPJNZgBwKrebSpc
ef6Kp2+t+l50NvJVAqmoiMcBK9fV7atO+5FuNDwtEr5SRpKXqqOsE2jwGESE
g7paLi3lfMqNnb3uicsEa+Tq3/eJ3H9JA4oS+flFwB8Mb0Is3S5CC20lxxrg
XbHsUMydX4aNWaMCUxRIBYD2p+cREHI43rqQezCWSaZnE/XPjAjsWRoZ6qnl
niSFR/VZ8knhiWJTmdCb4hFJPdoMZkxmfr7gyMarqOpnG5RD7r7GCqCWdKU6
aOKCSqIH9BBHoaV5nAsWFgKIXbBTXal6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SYwqZvligtQ5iQcQLT+ukk2ofZtkMeXJyhiPzIj3CoRZPzegyOPP61qGNJPf
cDY48JvqF2gf7ugSuZkgdU2DVsSJZo11B9fqkOvd+DonUnoEH995lhluya2Q
YisZPdFScpbvzkSBYCZ15BsyCTqXOTVj/lDvGN+sS9WEAWiy2Hg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WDB9NkxZWtCKVlhfXLFKu1LGXWeDMkHKBQHhKW82WUAJH12ku2n3CZoYXKM4
nekIjAX/oxN14UbQ18zBtr1V+UJ3lmHPfnBXdHroC54aQNvNYT/uvB/2kn7I
PbNsHkoAjiGj2IU4BfyvfCWDdcxeuJtcbEVonTkA0WmRBWHDr4Y=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 46864)
`pragma protect data_block
hxLAcs8MRBXurQyIjqDiO7nIe9SOzUg56lAZ7a0sBsFTggmVYt/IA/AEHNOk
++2mBtvELpnRULc6G4XQGUBdxP9cIu7+SI5c5v0kvZp+5Zng5GV5nEiJXAtj
G0ATff6PBPLhQwWVXgdFzOI02/ImpftcRPCH5dT4t5Wuo0jTjtVV9j8yuq9k
bQg6eekB+ycH3L/4hQp7Qa6F5cC6YkJ52qm6OZoc4JoD+fIwUkCJeWjt/eDA
IkLKZcNbdKniAdD8/x+x+cFfkNFWWDGkaxMB0kdMrxoDDR8k6rZfIolPGMZI
1hJ4peJshRhYwpMmy6Bv2sQPYeseMl0t32/SbvN1s9lacjJb0DnzMkwYamYP
BReRqFFee2DSRu/9k2RD2cp9uT3AQ2Xx7kkK/yvC57ONJFNf+KN+Hycc/Cs+
cInEUeK34sW6xw3Qu9JcZbJHhDSVSOEOJZ913mNaCRNyuCtacPyd76qTbj7W
Wh7PjkXV6JmkhzO2wbBgLPfqfxtYoprlWvZzep5X0cchFAje5uKgIgvagbz4
e1ocZdwgUYeSDRZBOTTv16BfI55lHjvAf7faQqBW0rMhjdcRA2Pl9+zayUGe
aqG/SX1IBV/pIzSGX5jp8sjbWD8Ps9v++8ZEe0meizePybiPoPIG3LSOu4LP
lL6nPp5P3/vALYPECbNdDhrHSMZFF4lCMB5wrVS5/7kgQRaujR0wV0P77vRJ
W+HKD8sCYDkP0cs333W7+QUW4JjxJ7WW3jjqAI1CtUi5rF10pK50TfcNt1Zh
2njsniElGrYQeon2jQ7M/JvCr2z/RJCzNo+IaT85AhecQ5j/FWN5YI26JCbD
cRJQMG37P8ENB1WRzt4jS02i9KU+fCyYAcO5KVuyB9e95YPxwXhREZuxGANp
wcACljkPugfBILZW2fCXMuP5kQ/q6+4qA4bSfkzo7NJSAjmwgMqrjY4hbk5w
TxsWTipadDBPJrdRbalAKIubcMxY28WR6uU8L9fa7hhiDb6GDolt+z9XYFxG
oGHnEjI/rA0p6vO7Vt9t/mASemOwm7fXiyiOMPbIrdvXX/XxDkgPrPqUcVeO
s4QhGddIpjAxPcF92mBryeItYyKc+hOVuzn+UwbrhasBYCul5uWW9aIwsAb9
Xg8TGE8IoVg/PcCw5e+kbLq5GkvNfvaIgcQIz7CqmsLivfbWfm3ocFspvpmQ
Lw9QlPxZVmOQPJa4pbhVbfh4Fpp+zSy8YvCL3cCM7BxzxW07gfuc9i6sLgpm
grm9AvgpzEZethvymXmeyO+BZXsjkes0S/OkzkHKSaLw94iMapcqpzqqa102
HzTcZQihYJWqPoXibSlklrOylcU7nb/nQv58VSecyEwsm/Iu3CPaaT4NMLxM
UWmnu6vSEDssjm9JkyKvlWzoEiPTR8eJ2CkubXQV7IsH/4iIJ7wrrDIuzJrh
Vo9wq4MugV52noFppVoGovx+DQkjY3oskNavjrH1HdG0ziswTry1BX8+RtTT
2TYvxpIkJKNkINSi9ifgyA6aTK+J3F6Gk3we/yam32ZlthSDTD6y1+m2cin9
IiCdmCOqG1Xl+CQPYDz93dS0gliYEAE6O8cG+4Vdl1gIlh7xUcWG2Nljndjl
ZtmPHAWbDk+uz9wR77+Iv/3FmbM2TlJM7joa7YnrNCIt3r5NNRMpdzsKV0um
BIE5VTb5vWrIRWal5Sv6a1PlQSLSSM2pTAUIRvzfG8ajsb8kkcQoM8Wtkk6R
ApjEgpq8N2QijEpiXZsXtIBgkOJ5bwecX59tzsGx4HdfszCYBS6+HFa8/Av/
jiuueN/k6zLF8Lge/z8mr/yKtk9+jq3G/aUbQw1GNazTyuBQ5+/Lhfo/4a5X
8810yTD0AfZ5O1Vj2lLE6PbrMi2fjjR4RNMSyb3CsJa4f3DEZj2kvSeT87/P
9G/ofkaWGz7t8Rm8UGxRv3/mRGmTg+hNy9Pdzo+f+dzjFRASbb/+OIW70q6t
iMwmUs2cyENxydkypUZbOfLU7NIdyDBp1u15QbyfmTJ20glRFnJdaGRhvdgA
y3XesMJb6OHXEqBUwsGSsYg73EqEFQbJsAItZ9nc4ql0L7ZmSNduqdxloBRq
9WR+CYLNdKdsvDs/Ezqv7yv7ISyiojXZqWnfcLm3OyIPLYdwbSoemqmPO7Fq
AMXyr1nelbpIR4i4zkBvbOwr/9fktlUqygSF4hQIQKpin8QRpqBmfC25kZZX
L+owhNy01wEFvcOt2k/Xn/1sZwLfMJSCb0/DFP2KlpxyggK89k4hRzNaEPr7
wGMK4PoiFR7BBaqLcXJfCNrDWf2b9XeREIijKPoJG5pLyjWdQjLsGJwDeZiN
uGl0YahZJUQVJ0M+a20yMo7WI9ObyAvBRZE/rASzVlhcxplN5+PLp++hVfL2
xsii0ye7A1LzimcrJ4Ue8HhqUNo4alH9IQNC5D02QjU0/xa//96hAwVjhgC8
56CzCHmgfypGovnQhyG6KBDDb06jRz7HoTaRKT8JY1I8GA5ia8esFij2dVvw
CAvV2wL6pdarlfBOb1fqB9OFgrvtaOV5UxEINcNHvBSqcvLYppxDgA5R8Q66
nrSgMMX3MPLXUgtMWZBRb2yHK3EiI0Y7DUAmhAox8wI88BqGTStjJM5g96h5
IsMfJxKPxAPvUxnOlBUKvw6gG3zr/D/EKveOlbrQG+RogfT5KEnUI6c0hIwd
SYQQlMm0qBwxMALqmcH9ZoCaTyH8jZ9zdAHHAhAXDHF74/Ui27KSkCo1lGJM
zRW4/azR/+DOUudSUGOpgbKLB0IQkWKsdDJ/QmCHvGA4qYDFTVbkd/Z0z/ma
4chotrXypucVglluXABFKyfVCkqQbX1FkhkN4XFCZdOtogDf23xjOTRHfS32
esZRJ3JczKI92LZEkz15j44MI37CnXXV0o6pImOfL3Xpl4w0jbLxBEJh6H7O
T+ga1moyEgFHl8LcNXU5jr8h8TwkRWLfJ/EkYRaXe+N1nZdt7wepBGjGfutW
wboXPdJM2w5G2ZSPdrSUHXW0tH3dgRI/rx3v4IWDBHU62KRRdiXRo2Vd4IkU
eSZ8ewyEKPLMKgidjjBG5dB8X1d71teTXc1Jj1O69PDvJ/biY6M5qkUGqNa6
ylcXJ9493YkQjN8siOHVuUzbIEdTZVJx786dEDrs2mqGR7PIQrWVwqvwT2g/
IKx965hbsTueXQ9Szmkjj/f4kCba+/BZwS90oGsQtFOfjddxx4SMALOZOvBZ
7nyomIEBi6SttLDKJiyHV5eiE9ZnN3hL0QlrAHRi29h1bdYMPTljPxZHLfQl
fwzzzh/7Ut5A3pzH2/U6IAr3JZQ/ZYfRkQgJghkHHDSbDZi8Iq/b8MEN03nW
fj/yFT+YAyr3+VVTr4BMPuraV+q4D07do4wp0Df6U++QRNHfPe24pWqtzylB
vWBFGH8Wu00PsFXWojlhnq4mVuVzrWHTMXoofzDBfHcs/lg1bllqVWN23VEz
dNkJXd/ocjbj9aJJdM6/wEoMgBFA7LdSTVQcwG7QWmlhhIxMr3+BAGvFV3YS
VFG0gvX/5DxQ3rBMNaW8ZQwvQCtUfEf2vmjUvMhjSjpqfUHDfxJkQ6whrjRk
iC4YijBlcFIgQqE9UIW3z/I25ffrh5Mxt7S67nPMJ3exbFT4iredT+Uw0eSn
pcCBZyoyssnB2+GDxSStVXSx7P842B3xaUpqjj0qlT1uVlmjWjvSmwIV9t8S
hHW7zTHbB1293cgGEbhVl2JWxTkSf+PQYBbWEQDgNTCnmOFjd0jkcCYcqhFB
SmbYLk1Cmsl+6flMQ7OZ79WRR1h+FutTXswS6xH6qV6UBksMccTZJVKjhx+L
muoz6W9CmuAXoEINXvUvPPayLrgOMHKYztSx6hNsUdo8k+qMMAw6tue9DwUd
bT0FMrE4ExsMhmffZq5MTwDdbI1ibw6r/I6gCGu/AEj1jwFLbr+qezHA2GZY
7NN+Jd3kQo1sKsmxnwYIYx6fHSlCQA2k8dvWLOIJIwzHel+lRIYsV3v7gUSw
U33meC6b3iEVuOecpcmZ8fpMQ6El9WtUpmqisAR35RYbhYKNaad993971na6
++4TPqkwhj4DA+h6iZ6k4Vv5YD5TbrG1Mr2sBmGlPWShTf5igqYN8pDi0KN0
tX8Xevk8RUZIklUTAchkXvh/ot1gvJRprwTBpsxoA9Havrgg/o0G0W7G5yZH
gvFlSbuVHcR+MmCyxMGrtviJBwx77P/FK+c4ebUb60pTTruFqWwB2yUwbouJ
jmfBR2mBREQHcGYyGMSLimZOrIjHwrzhePGA7lvmucZrQaKRjizlwf3hm+JE
Ik2C9Se4BuNpHU9OcfMcf+o2kG2J+t/CYE/c9o0BPz4A3NcIc4CHU45U9qF7
ubcKDKJf89B69RfSAiT3hWrkNPdUlSYxAMLajCixydCxqtMa/uvDl90vBByz
wcnPl/br3fsDSq7ZmJS/n4pKKvkn6o1kyDAFZLrjITmDHnysX5Y7spEgiDPI
22YV7fkznx84UAH94FuxerkuVfVTtgm7eIeutu3CYVK2ptQPfhoijLPuwwD4
U62pyOcl7YNCB0hrUxkGa53vi73yCStAkor4IUqKv9Ufrm6dQs/0zPNv6Ay7
5h4Vwso0UxHT2IZd3kCeGAUToIUCChfgBK7BJloYO6KOQHEwLi9Fa+/hcue3
qrRyQAi7mVK5zXHMgHR7jfiIsqaiFBOwerRyWa8AHsaHTxpyFSTh39yVqo1d
61vrRXubrIR2aSzQ9I+vz4h2ds0YLwXcS/b0kiPS5xJ7uGsp/HFqC6rUDapn
JzKFI2xv/9/wULG+Vlh34Q+ImM5kHgx89w5N7eGOrDG4x57FhH2Bzt5X5s5y
TATzjcU2AkJG2z0Tjy7KMMNuDxR8/yuPsJa5BoG7zBP4uLuBgY2hB2JRKF+t
dvuQEIR+rBm0CpnB8BM07vYVK7Cov/TQOSSUEOjCjyph1UW4QGle1R1AdcIz
sY5D/dbMpCSiEZ3R7qXEoPnbKIBg3hAWR316eg2vF54l6xMfKVaonVFrc6ge
N1bZGum/h9K7f4meSTITzQkv3AJ7x2Em5kWc4Tr66KCoXDBGn0gZSCkAwpZn
TXrJ5F4msik7kf1NdM0yusH4hZlpzJoG2MrqDU5TSoWtPWT1QfYPoxGb/PD5
g0SK0k6HeT+9xwWeC6+Xje5HN/g5NPa5UG3cqVGX24G5+s/xpYbiR8zAdmux
cZ+Wj1uhkRW41jXkl8a3tueWZZHpjzVWHklK/NfyeJeQOEzoK22b3ao38vRZ
ZvndCiP3KwouhlHaHoI8R3vh9uDw2nOr9DLXWHIHPGqC3i1R5F0Or6Pk8h/X
1q6BE3xQDeGIiXYA7GkdU2wlsu7eF65FhybVAH61qLIiOFH9Ni0rmGXuy5CR
mMuZD/keJy9DCPXw7yIqzgjrJy05uaLGiPKuICyHYUTI+Rh7jPH+bY3jVjc8
CsrJxmJfAh3p9Gxm+uM5iLd1evBlas2YfEzTYfkFvxNzYf96Fjb7f+tY8jqW
SzjV0syPxPPO4XpzuDGu7WoO8htylMCvP8I50IbPXmETX7c9vFwr0FhCTpjz
Rsjx7dZzy/L9rC38q41hHxQaQrxJx2hDpN1pdQNsWsd3B1hSpk1qEhAPFYh7
5ik/8aMh6OgXI+7NJKig9nFBbWbrXuN9KYTm2g451o9Rkn0ooEcGAS7NI+sk
d4MlKcRt0QCc4aUalYbmwI8+OFpXPYoApGza3HsFJu5gY1MdOLeAwRMTC8+r
+JeUh90CaBVsCgbDUrikfrs5r8bKYiI2AymDXncRK+z+HiC727Nl00c7aXxe
zL5jxUOTLJ2OJS0REDbL5KgC0CuNrIvPvIHYYAM08J0i6rXqFZzTUTiUrOBU
+ke+O5EmISJNo2w2Xprcuk1Kr6m+IZNmp7Whh+duy3fQ5vhiMN4c+lTiFIaa
3XtOogkTsQ8BG3eWCLonJcRoXyVqRtLdpKbeQgiBf69WAl0s927R5142IWiG
wWTctnvvDW6UaMm3ACPJyROdRKwtPbFOk2pFdE58FVJ/kcKGA0ojPup55/Do
XuZhkEH34RjQIUKEEEOp8bNzHT7B+AUYE9VRGOi11/ywzte/ScoWkDQ8Rydu
ffa92FZ6aZzx7+PBnXoMig4TH94ZBSIC8y33Tcc7ixzGiYXDtrJMJ4OJfR0M
HJZrXMKffU3r2gfZXqp6LE7yW/IAab9GaeGMyJ3sunjPXqy4lCFZieMu2yI8
Whxwcs7ADHuUPF4A9JyXQ8XnlV8MfZeJ97WAPqDL9Z7VhTQK/PSSWsXEjjMt
dy5oy7fiv8bb3cMIXOrrFeDlPkAlWeTjVzjwdmK97Sj49GomOfn/+VMik/aF
e/E8gYweV2VdK97dchgdGhS5M2WUAJoIW5yoIOfocsqUVWCJbBisyq0+JhF3
/dluh48GmJtNoAaEJOjYk93NTNLuzp+RcrnYzXaWgpd1aNuY7CPgjtw7IYzm
OFYf/xseqEyWiwx0sgf5o6wUidBt3Df4gOIBNXJf57hwgAZ9Mu0nEvfnJJwc
WoxCaBk5WeUpk96Oedw8/DykqVU6VTFN7O2rVOrQ6UgqSB3veIDfUM/c7/jS
5odpqLLkXZ69ElN7VlN09/FeSR2tN18e4i5WYq/huNpevNmUXIPaTKAra1J9
TP4GaQ0sHjLlSrPKRxxlzv4EoeQXAUo0vCtQb3BstpUBVXcEKR3J3gFOp2kg
KkxSct3y8opFRUKXOsmidKZvMIdDRqKsjoo36XdTPptXCGFt6IjK7cbiDEnU
pB1fML/HX+5yEoiC865lbWFX+gvFVJvyQOwioDSU0SSC6V8JfWEMq/9AacfQ
EUKaJuzmbV06nmqsTia1IpvuAKfk7LsPuFJcC5C7okBwqlbVAwC/BK7W+xEA
zIho2df0f2VmtUM019e8bKXVKOXiY1iOGuKqZPOWpFIIZcTOpCMAGp3jvRvS
9atZ8HZgQgrs64vApom0ilA4L5NQakuluZpKtDXLSEWI+V7s7DLNvC34NXib
m6yhmZrc+gLApjEXleLhi2E86IgiHnRfD3VIA99+GVmDWk2Vwut3eRd5ZG41
/lF5c8PEr4zuNg9F5Np1bRRR3CdqC480lLD+4FQloPq45G6NrdiPZLsOk8Ks
u84HQag/95qvVx7YJji9EGPXvcS6O34uR/rCB1vQy2LMNHK687qXeeAVYH+Q
voi8CZOwWz/BVdGswzWPU6HRgRbfvybRMP5pH9QkFk0hmCANiJGgnJmFAi1N
iRDHJBjX3DwcPKfBY25HihegYAlgAxqH7s1eMBMraa6mJTKF+ViKu+HdKxCz
8uW3XL1fjLmqPf1ee8IRk640mQTln4zRlBFce7Q/PDiR3RPYypnRA7oNaFT6
HgUG4aTxRAqdfUfuyUhZZv5e1en4rENyQYuHJH6ma6R5E5G4DCTqJdC9/OqW
tORUSmhOfk55xR3wgVp5ysOCCiBRr0e+GB8b/G7pB4Na+xR+0n6R/B0GUIvS
ZLVK18NpMbwLwSvARKf0H9mB7NkPBnnR32DmWbP+xrVxQOy/DvAUUqHd16O5
eJhIViTCijqsugx12u0EeBnysnekEXnZAnG224cOR/NrgqzR0i8XEuPVvcO2
pOqjyHH8xwqxbFwnmI50och3FPjXOf96Fdfxw+whuwGue91IxyWuQMggp60W
Prcnrk5l6JUzSidL3IR4HcXvXMLjkeYTnMbZ5u9mpWDeC+oIOtffbRl2gchi
puzbeG7+kXpzPHkXl19uWzp7wa5rL0aE8Oe/qYaFNcYkHQhU7W5SLuchZHMd
UvnpyWE1rny9iI4+MYHeX02Dk8aXrDbhCV+0uZ7HnnskZ/D2ihYSaFoI81KB
6WHNm5iJo9XP6SMqUa5XyJP4L2dgaVRV8qYfmCYo0ktVZwehFNljDi94AIgt
9vhWmyRzn8ZSS/5bZeNRRIVMU7W16qH+pTyj2O/CSulGkpO9cLLc6Tz7G/Eg
emllpv+fCLNJwj2TauYxGgZLl5FGLk2THaz8iNAYcajhRhZUxVx0WspGomfr
j63KOrYB83g9QMs6xOVhDy1hhADp0ILmOYvk/mAF3GYNvAK5Azck2YVWbaAV
swIsDmjrYriJFX1/kx2YkerFPWC/BivJspeElfAElBBKMy0VMWwn52+81xe6
ClAgNLZRVexsI5kgCUZwMdK88kki0DxUju2rCYfdQz+VpIWpTt5Eyn+b9lXX
x0vX/OF/nhseN7H1IE6xuErIaC2+jYPp5GQeRQ0DKQonogAZk44Pg5YBYfhc
guUw2YI4Nzlb3ggCz5Y3aCblJ+lXDd1a9/xMfmNmxgfcyyY/q7YmcEd8rvMw
tqXgeM2No6I5wfCuED2bPTfn5UtE+nJcx/VuIH828E5n8U2teL6DrwRXwMJC
Cu+doywojNdCETQdKV/Ce7h4vil2/vRlGHsRKSHDpJqeWuzRodrIH5jEj8Gt
pWZAUHIRXuis0ug4zc52Kf2h5RHgnYXqjWzAfkduHJrCLqWjNAMm01eVVidS
MG/vGNEqpPJZWBR9Fg6jRYiR/5ZDeYSI7iF6t/S5gCGnddXLpKJYVVttKZxh
uObPvp1/k648j2fqPNB3+FwlgL2zBug1un+ePO/NPfWApTmWJAxCkhy8NSmT
OEjveLxPdoRqhlCrPlfoQCBi53O0Cp/X0YyFue7c0/5IHiWHXY4CODY31UmM
GsP+9ONdc+WMi+botalWoOgnKD7BI1CFyGW2HYgaRLrQYbZPu3ELrB81rELw
UAOTV9OC5etTrX/Oe2dVjOSlye/CkXskkBpPPZwj4SqqoZS4E2gKrtBf8ORQ
a+lDysQQyRraBsNmbAEsIYt+rJh+/YSqVT3Kzte7pLNesHCl9mvhoaEVCVvt
VeSGMz0/kZNzUDs5QfWlcAOS5iScxLlypBONQItlKMcMJFpFDyaFIPY0lwi5
qh7N5ifW8rvfFyn65dEIJwP9q2oBYbwn7+h3tbVzN62717baIkyOegMfWkxM
0tBc1QgWQC2HAW+eYbanJqrQXajMjxDJ90VUbsYBer+DQAg1PVWoZ58VcC+u
bzUhIQolOq872pi191jbYwyd0p5Mwn8xBlIUVfqhLNK5ERYrAOHZYU7/6xQ9
bzpI48+Hn3a4a9shNBWu15BHK1mGcPakXfUJK1E1x87IPeGlqbRg4d1TemMQ
hN3XUYzJkQm9icoEYyVwGqEnjXvlWTcpvgeT8XBLkcHPp6dRGlM+3z2KfPai
fRvjJ+vsJDwTI1K9UJ3rzdb8tFM8hymR/qruH05K/sV2gCDt499G1WCwxHnz
Ssg6v9Kx0H/tFbmOLRzmPj0o+BnDCpjhyuT0t2JMEeQCtcEgeA0FEU5MkhHX
LUGUyYWayQAusYtisjcJZP1VCfcCZz86zuQOoSTK9HEFfAATE27AgY/GCGBG
+G5ghAM0xpoWPt87p4iGB4slIW/xXfL8TlFjUVrrHjmcNPYTwynqPQBMynU8
SmmFRRU109dCgrbmWJkd5JCSWBE1+oWB98wO/Qgunwm04SjZ2aPda54N87W5
ymdFK5Zh4q+uE+NMKGczIbLIRA96Rd+JuxDB1ichMMYhABHDytwFaCXNJXDO
bYhSv+ZPWlp5diWu3aZksfNUspd0m3zMgD9NPqBPD2aoD9Pxz50EbnKi+XN2
JZlQMl7sE/ZESKb2Y3tHsUb5qZTmubCFLRoRxKVEoOvT8AsGQnnlZ79P9e43
G8w0ohy/IP3cy7FCEZWzPPn9wo9cAMpyEWZvEkCr4bsD8OHlMykCGddnHacm
pL49jo856bmzOMO8usNEbmJD/CTaTaOA0l89qxBkZydtBN4mGxStyuNmkKxQ
B9QKMKpXNaCdUWR76GCDTlhqjHihNipg6yJVhH5/0eDCTNTIRAh1j/XAy2LN
pezHztRkx1oDb4Bsj+yZoavmJQi/aLohilUusG7ztV4Sg+qSonPBKgQOgDoA
1KiZ3P2fFUkGJnw1E8KbQX3UXqMoVRXx5N/TF9rpRgWTOjYtcDkD8aOu+miv
8Dio8wAMrKRc+YgBSMCsrYmbO5nLWps48bqDyxgAC4CptRKQnP2xDjYVaSJX
usdtH+aEJMCQNwEKCo/sk8diuutgb7Ru+IrRRaMu/PDZwVcs36e67hC6+43I
NYYjFkp42k/UGzi8rmpZ5v93U6eDutxBq1dgmBQrR8wJAnsw0cHGp5oHyqIk
kH85BE4y0jhn08aPgNzDt8uAWFu/Ifxu8AS5+PzGgLVPs8ZVS0F/H6oKsEB1
aW7lfEyVEs6IyPOGGdIxHXlNL5TfXNLxL4mw50waQp1sSxvqGUh79TJ8Fdz3
VEJ9X9oko3jGS4z+1ppSU4kg5U0FXVY7lUd1WvazQOxQCqqbU+g6k7ogY5gz
kyh/JwpXGPzUlXvt9bcJLv+J9a6eJbnQwu0HdVqvHeNJmG1E9sgxG0++oi/a
GWoY1A8bcYKbbtn4JOrCpaAT+6+oXv8qIZ/t49xtPKW/S2y3vz0uuAofeqBk
ee9XTkdTL2LkVCuGcypyrs8HDY6hwQlrMIujjXzSa1PwMhyHtzXArbBssGnK
U1qCeuLQ6tuhxdGXywiPKSqcxkeZvnLXo+Qm4SGMebwy/4pBYY3mrKKb5m/A
uUXywTYle+ZgMiH3dk+pcXcs8RfWD+pLEQN++ZWdzmgItSM/ETmu+sHZtNUN
yN/NMshfSroSyvplc6deJ6NYghJGsB3IbBqObpF/YoBMXh+2A8QpKccHO8g1
dJJMBNc3A8FuSpbaUqJ8O45fQud0pJ0WYJSHdSxpOBbpP1GUh/N7ZD3vAR/M
umusataYWlZCRaeG9DR0A2loyYUMbzcPxBZWvyy6AAIqZhOAkKbO6Fh1hgq1
bq1THWo7F8a7i35QkwF76QwBuHp44buO4LFfAbgbUS6wJBO250c3uRX9J7+3
oK7dQ9LQa8BnYDlxlU0Lf95eVD0nWlVvXEhqJCDeUgKmKZbP/vYwK+oC655r
SBtpqEc429DwO6jron6Fv6evpFss9SrWphjri0QCLkeRPb/kbAUMXsWJ0oJE
8l9h5gmy0Ruc6Tzl1G3G9CyO/TzFfc0rb5VClP8VKrYKqhU0pjrFXDvM4JnI
VLh1DyW1o3y0yPntEcj7h3uhLYbyxD1/rRicmLEXy/zBaajOkZyBruytbBlP
JKnqmYvi3MaN3+pA7UrAhiupH4T1bF/qrT7WPI6EZ6V1UwJXNDUYUQfxGoja
/AAxKz0G99SXDI3eN0H9UtvJREQsxiQtlCO51EI/i2zSF3Pn6B7bLKYf/cwM
N9o8lujnIFtpGSWRS/xmM9nKCDa9IWvUDJq64rhKqJaei9noF0bW+ixdJbMo
WXbQRVrpk17E+bTP9mW05zq38pBu7tzzwWKs02MNRoTwFcNLmrLViYj2ILA/
JU2GIyLcUyTXsDf2iZ5SQn+7piNK/nHmWWl9SJvqNFD1P/NBlKnAsrIvztOD
TWBmQQ2ALwMdXbZr1PPUE2H8vHIbfkcZjVuCJzofxh8JN67fsvL+JV75yB/H
v7ZktAt98G/UlzgJiMA3KMrwB1rw+zfQsZlK7wM3JdID0BZeGspRVxhqIKmL
+LTOjC4eT9oNnKy7LFPXlnZEofAj+b7ENcZAPDK/k20y/0SLIxVv6yjbJYvE
IOUaYGlCSBQCZPL1YUKSPXfg3Bulero+3sIfSQ98US+F1wRQEgs2YnlbrJPV
iozJaow//i7HY8PbDrE8g2OgtCXznUvOWUKU11FloS41/l9tIIjOXLweO5Xh
o8PiiyW56skNLup5hjhpsgrT5wYv8pFnn5myBPc8YU5YB7u/T10faw/gH/Y7
evCHs7Oe4g4kY2UNozYFocF2ZUkMWNqeCgeM2WigGi+oqbdybVUOoPcy/ZKj
q29BwYFeWb3fCdO/n+QVhC4sfZYpmcRZO0QIXE7nLXIpngoCs85fULKqMBO7
8Nddw0BFa9TFPNV6TQk+5qt+Oj4YnFC+zOx5RiUPCCtRmuK+107TXGNwNYM2
ohe17yqKufNwI4+C3gFCyGpvy/Mmgj34DCipO7vFd6RoFxqtaDeC8T5mbiwH
AXnJ3WK4oE55LECSWlKKaUvSXKHjHFf6heX0BxLGCQnO4fVK6ryhXh2sHj/x
M3S/7+ul6DZTnLP3ACXAo9ouAOfquefUVptOOBecS80OMQ1B56bSqzRyz+m0
zgquUV61+dfPQJGZONuzyaLwIWoZ4hPmKkVXqeHzM/GOHG+P+7y3iNNio4O3
d3l+HB9Se8dS7uaRSVKbuiEeJ956ULl5Zq4Z0tI4Hg+RFJlISXcf0NWMiRIT
Pl5R+WE3fE49KsjZ5JrVoMfepNTaFgunONNgzD7MMRvAdYPW9c0lFel5iYFj
O9gLRWhuELN3uJSkm6tcgIZ2H3CYLlloeqZiU+kf4/LdBeTjdP1mJtBEYrme
pcHNPkfU3yFfn2otzc9uPRGtOgtIAaGKWMldmY4blDNpmZL5GYK1TifJQiV1
UXgwgp/b6lkCXbcdcx5gjHZeA9MGBHeBRxjVrgzcpHaxaZCPhGX/LnmhPio6
0uBDY/xkRMB53QKqxwEAVvHJPWa0dLnuoI/PQqcQY5sVK5esOG0JmNZa8hyS
rtMpC20m5ZsenR0+nT6UMwa0v7sJjQQhmnbYM72jf4ag8mwYm5acF7JNW9lL
w8F6YNF4E3cKtWidpzap0LkI11Tvydk9C3N2+uR+n5u1jofwjxjig/Sw3FfD
gB2gHn9HXaMmksHgTFApGHlMrvDFMKHBBufnBK6VW98wKj7Rwtwppd2lO5dP
Frr6Uip2tq/zQqbLkszIWe23eT5aVMKHmo4Yg/cn19GVwz46MuKoiU4n1uOV
ajdK5OETqKuAZ3sdYroPLjaw+KvOepwC7aRQjfu6DUAXXZpS7DCqCBHY04MB
IgeSzL46wjL8T4VTXNp7ZkrXM7cbWUlO6c2fsAbYRnTeeGZ1cGRcDcxlbPfM
3CAy7uKfJiucp9X6LMMjtFjYkeHArmpkL4diEl4Y7fBDDuuE5dECDB2aBMxP
9KZml0d/waFxkx7A+KMU1XfILXHsb7ODCteqikI6sV9QUZSPWrMo1sup+4XO
hsYyehFpknA68EePPKzqGpjRoKhajc8PrZZhdaTKyTBx9t3biG7+8sDZCzRr
iigLytayFySsZAdfoODQXj/EDrg+XZ9Aw5WZrkfAFKbtShs6As9dqsOvSGXi
UQMrAvPX4fitPk6Ja8qjLi8rfz2OkquCsbOpto2gXuFF77Og9OQPWn1N69i5
p6qWMDe4q9gMsuL2b3k5V2ttJIQPPlkomAURVEKqLN+o4EyGyeWFkeZrZuWm
ZjdO921ZHdvFQmJAUfzJEVoW77ZEMdDGLg+zMHbtM4N7rr+cAVKvfjSGqKI9
PBl9PHs6FizzgTpyPBgbIEvGBhhPMPdNfazAUOyT6vxmQc26TbyurBNtVclU
t0VJg4Gux7keM4nFVd4LifDbz8u1gywE0CA1i/jSeXF6WH7SgzvrKA/Fvm4X
jwcPmePQwp1w/hMemkTsRPdFY0HEhmHLxk/CEZvuMgJbmjfmK5Wker7kcpKv
F0rOxX2NF8yvArWQuz88E4AJ9oiRp3pRrRTzi7pW2Fb2D1aZTDCltznNcklA
QQWknLjir8drt5iEwaf4ulQM/7RzFA25vfIiyC4MeEZroHoC7VjQC4taVFl8
EqOdio2/cZ7D8CtqOnlUCRQUdozB9SH76TYKlVmczbDf7wKWlzjh1ReN4R4H
Z1jIh9iG95mCyE31ECQ9LVI5rwwwzh5XMCRT1lV/0i8gYa/POh3D+14D+cZ2
RabPbBZTNt5nQzWfuv89BHjr0d45C4JUWCUEFLEdJxDBHer4ayCXACaT9tWk
ZvttBapfyLXHIgyYe42KKp+3Suo9SpHPT7BZse1jVxkkJqNLB1oUW/WXnO5v
waNiW18zg4LvzZUwr2REH0Sh1FXzt3IrkS6SiYbFIqw6KOUpuiXQoAfbVSv+
Fj5etrBTvxgQjgou178egD/MHjspZjJJ+IGqYmQf6IVdrWB5mAtbW4qjrgOY
FkTXbYFYo8JUFnqYTKMc9wcWy4zIcnmoj2iwZrm9KNVAIJk6bhNFGXblHxbo
XfOevpYn0jTkOftuUTwu9S4NTmUVmEuzHg0rW2qqGJmVtvKwlJpx8kxMYyXE
0UB21cpUM38M28+Q8Jwn0ApZvqvf1ujaVYgXuYK/tfupFGnArnrzma1QgSXv
UtwryT99v7HfV+H4Gv2oFzri72VBIMuBzVBTmUHLqjJIyS6owcblxe46XLnp
H1kJd5vS+Y9oDjuaAc40NYz+CiLsafFSmC0Dse3/T5ciWGIRxTEE9dJ5J/G/
YzbjlpT/oG57V2uFLSoNUMO33OQ1Te8NKPZg0gBv6HouVQ2h2ugWSkNZO/HL
6Zd/jwSY1QebFrBeafHRVLb7xcKyzP0FE5+PUb33BfNnavT8x0o+Sbyuu2Ai
0i4pSZvEjEvUaLevg1/ITV+m9SF/hz6TUZRcadAwi6X3cE5j2EhclIXYWstN
6r5fqHZWqm+hnTXWEUJ090HJ1yd1xt9OqJhJRBX74JBZtsEo5CWRtX78CVvR
YitzcvuKkga7qH1d+SXVYuHFa7GZ0EcatTNcbR6FrYnKdRe0xYv6J0ou0Rpz
HN4PigNSSWMEn/BsLMg5KgWNosdS79vmRm83uuTOjlP5FdW5tW4z+F8rbdpG
nU8GBi5hqLiL3jQcHDKkKhGxltQfFrKmv37Ha1wxlnkj+77x/ZUPpxjXEhLr
434s3LbYJzn33cxIWCZfwajNZXKQr8ivaWHDEjehP5CspKhUw8bjUKSl80IE
mW+JRduPVajekFqad0hYw92DlnUNgp9MqYj9ZQWFE2C/IktBw1SiBRrhA+eM
NrFcz68RBvL+bSVCsEfCBLDTQYr4/8NCDVwe9P3rghxZuN9oTkyxKUm+rFhC
7Lvw9De2JyK797KI6TAtDXOXoosaB1DVYnIrI03fFHgW0Q0YouODxszZDd7K
vtiz0kvvzViEI1myeILHKcNqOj9eGqKzpEhJsj6ND/W4WR1RBFQH9cfi4pSG
2dx82+BschBeoe6JqhPxeYk2EwV4ZmW+sFZqcgSWl5wfmt/U8sw3rUNfv4b5
/CEHdLeYK7UUJWjrn/nXp0gXPYrwnvcEK274dAUoTxi2etyqnZVRfhEUuGTi
jtvB2nm+AdzGlaS9W/b59j9d2nJztx3DhTFOJFCxs1IR1JSO4s3wk95HJzcF
hhLJQbSvT8EkLJYf9EdCM3Dyn2/rVWGhmP52F5iwCZgIy8I8qjQf3OklDLB6
WO1eF9B48K9tR4VBMxWG7X1RltEoTyn0qDjhcXsbHE2+7YB+vOtWJy/4RvcJ
fO0CXL9jQ5eBRKs/5ySlnpsNIJ2G9MOBwrkRVWBF35Pl7GdorbWgd42Z3ii3
n8xjves4o035hjwEnKyf+YEWyFJ6oJJ2O9K5rPlDxUup6bdCezY+6TC0z3xs
8F6mReNKDFAx4aLkVPDPd9bm2IwoLmB5L17SM9EcdVKGx6jucAMx086jCcBb
pe66nnpkZ2dTopbkYHxInTrLYJ/KhXopJ5y8yjxz9RBN71QpKRJOkiWBtB9h
yEMpXiAeY05YS0uwQRDt1GfZyW2FMfJXYUnwT9eFVZhpD5FBU/1cJuWYjSOE
sKOvt9Wqoyc8gMqxC2WYE7TWTwBbfdAny4C3U4iv08SbB5U0jmOVonC+0v16
+HeiOiey/akfoTT8dUhJiGI5AMJTLhgNBxXcz2NL5alicHu9b3TrYnlxao6Q
qh4O6qGH1dhZpHZjHJ09lzQAPvyg6UQK3rJOJKb04162mKxHp76J/h/wi2Ae
oZoPVVCG/yGX3ztsB3j4aebTqBlj2AFfouGHCnqpWQJoz+Ulyk5n+1Z9S5Fo
U7vpMjP5jQfDds5qIwOIgKUdOO3FiGwvvWxKZF0LstWn6gqGgLeve9K4b6Q3
2hhQ7MvgI7KC69i5t/AVv7Ph9t3CPGs5WrJ4qUxZF+ysGjTb0vxCxFJGUReK
Fwc5F4bEEUeRSwyr1dPoiQRbLxl+ulGCEoAfaT0KEOZpJDwhV2wx9uxpLTH0
ZDokocnEVPfbxqdhqTcWWOOEVi7E8P2v4e5XkQdvR2vtqWcqKKXfAuQKZVWB
yT3Pjvxw9iCybm2sfZNCNx/gf29bEIfskKx4juAOu+0rj8JkRxkykaUwU+Yd
nCHPPjE7rlGIPHjQXj3mGsTLCQrXhp5L9wn9i/5vKfr+06HaI3AYWZrHWvJt
1amXogIWDdU7PkO22wr+QNnzl8ATLlTArYL8cNkzWWplIWpbqIE/raecqZSq
q2hiZNAU+1PlX5wFmVSmhmcmAkBhJfXgP8vb98tLqMNNlY37M/isEDtwrhLe
pzS7afZkiSN5rJz1s7EIYIcIEZY3okWAN2qhMbCVUnhKJ7s4XdzomK+4TBeI
7SS72qDJ29DGE8ZHdfm9NXvTLkevdWl8H1HsEq8W84IJmlyE7qmFzPW+VQMb
XZrXjZxcf8qBc5KOgdnSQ9cNOGzkddsONgQD/vqmc5/a0DmsXpTPFoOwgqV4
/qjJyr0ZmK01S/keOGxm9qd0SCeZobF6ryntS9IXb36oUYeqS+WkXS13Ex6f
4BkRBTRaAPPjv7puLe24IZk/P1FW7tYC7QVn5NSMdZ8XhFY/RNh3g7jen2HV
BoCMf/8YHXf7ZsxPKWqTIaIvJ5TrWsLuz7JaftFfOoY6fWHVSO85J2JNPDED
daayK2WHDSFBR3+404xzHuhdLy/D7yrzCj74x8xl1x2+Mv6FSRPf1WKQPKyq
5w8foIXnI1AUknoPvn2gwJcd+srC+m/+U590wPDOBdpdYs42zwQUOsQO5xZQ
gEJZ1jmrXVHmRxNsOLbUaqIWZ3ykuZM/v+pRfF2JZXToafl27yhUa5+m7eCa
om6Op7JHYaSRHixNtJD/ryIgwji+Ww33VD/+r9d3pvY/eb5bL5ydapmOFwwt
+mddDj8lGE/zPWVPWnD3N55LAfsa3Yw8uDu61JTxHe+2rbY5wSzrb5kAR0Hc
Q5tuLVQWGJQSTkD28L+fLtFEid6bN9EUxggjhlWwhVeWEPOKu+DgVZTCr7c0
4zvXwYu90FUJz6B3h2D+FuuQ8uf2w2AJzAcJM5ncEDrjVrwT4o5mtRq7vCfY
Rg/kcQ4w8fglojdeX/NqIqjuh3V5l9AOaClpMnFf4Zre73MWAOMSesBA7Vp+
JlryOZyk95pcYXKAVUHtDt0r8fYSi57D2gKF8e25V+WrlHx8UdbgEAVKuMIt
03nLl3g85k+DdfXnTZC+7uZ+Oxv3CEEYgfH/RDM37+L+hsujGONCH4acO4D2
UTqhWOh7eqEZFOLnp5rfM5HHfkRYgtmycaRonGRl7xWaMUzT49nI4Q0rsWwF
ZK6S8a27Z5ewopu6wrVE8kdJ1LKba2e1M+5ir1M4T09W4Haf3Smuzo3VUOB8
2tsavC2yxQx7/OwDqgyr5raFGucbefu78UcIV9eYtMF4E5w2Lau5tzi1txY/
dKj00B6uo06ib4OPhYErvGIHImkCGasaYnLvQ5SWun0x4lGUci8fOBhIjGqA
BiuwccVZtuOJEd1gSsqQZ1XATkmnWpamBQzv+0MOlqgK+JSdMlQM3v4JEdCQ
AuS0ARBpljUYKtgj8f3mY2ul0kuTD8Q5T7Rfifi8bc2TklSNsxkyfA/C3hr6
bUeO0r0mlEP3X2OtNBms54YYHhwAiKfUIk/j2n2tm9KpXkcBqttqfNDYvsmN
6BNGCUdvkZtkB1gweLrajTazVaKYkQ2csCABIJ3e8fi1kjHsSHD8KLXB2Ip9
ogA3ewur0TIBhNwnjDVxsAH8eDbfRRn9wx3fRsytiEn42Qi5s5xRU7NrIuUj
LSNTfNRK0M5jMGYUwov5wGZtA+K8kbvDYyC4Pn2mYA5qZh+F1Xy7wzR9k8lf
SWh31YwgWFjs9fzdL2R8RPuHn0TJDIp/0D1dJIZuq+lMY2EwMpfBgGFYc6Iu
9hU1Hitur9vrp7q8lXhmCRW1O8yItn71Fr+kQwFszOlZiYB5Rb7IPGMXnP2y
SRABeTXX1IsQ577Tm6xcNM2BBAmn9ywM/Wt5kF9lA4eGAjRTK/Mc7SxHwVij
UG5Xgbh7aqx3YWoeuTdlrlqvmiV9Mf/PdgbVmqviyFe9kV/qYlSJyhUgs594
M7N71HnXgb0tXLcrpIB2kEcBxghEwCNRloiAj4Q0PCnAJ4JqWYOrcKk1D/Iy
RusJ2tz3H4Oz9qmGaRtqJwPQ8ty6ddyW1fF5IBscoMyLuF9869vg/exxBPvg
o26bBF1X8F5vIiH+Wdw4kNlQkxYaWOy9PmfhzImFd11RWeHzSlQmoJiykvzQ
MAa+qjvkvye9GEvAyW61Tb2+HJFPcerOploQnHCnKVhKAYfXLw2odDShdiGp
+2FoFUmuLjYqnhL/oGQLVGfWrOieSFKCVjgHx59zfo9FnGTosETtZAGNr1rk
5/vmOADRJyomuHPhUQC9NjpPFJCEQMrcnyXFmuIpuEsoicILoC3wViYFKeBK
bjLosKpBPCOmlkjR8DuS41KbXo4Vbj128NrDHlsp0GMibfKiG+eo4cIR0fGg
qYFEx7QcOPz/5LObRJgbcUN8psD98nOFjGQF/EiOe7sfUAgxVpXHvG97UuYk
19BwoJx547SxKCUG8ilcMU57yLSz4JvX7crbrfqP/Kg84ewtmrRbAN5WYKvb
FyoTHiQLGZKt23rLHrjM+Tij083n6bgUVAXYj6M0N2ZUS8VNe7iMXAo9hXgK
AlhlBBs8px7NX4qecCCuuWGdg09Ton2w9Oh3aSszK0oh3oigiEijHc9xPJtt
QeMqAOVHt6rcKt79oAHhykuVy591Mny2J2A9YpdrtT9BN9KMrMjB0qRmfNaQ
2V4AHIdEuBYK5hXZnHCzE29MSsUrtKAHJErHPIlr0YQz0G8/7MqCrfBhQ8J/
eeWAMzrrM1rir43qjbtK4IlEZGk5a0GNxr35/fCA2czcQTcke6v+eljiLeEZ
FWUAjQQqoqsp68RYJD0mQZCQTDgBmFYPy2/RlJ6WuOLalMGQ9zBJnw150H2v
Va1q5z9GFjiw0e18oj3qOhc9vHn+ClbTnLmTwHwfrORxsjAOFwBXfhSLPREE
YeoloufIgqZjoZZOnPiRX3fXPB035/kYTLUCpGlcg64YPlFP0nAF4PAsh5bk
rxyv8+UwpRKuZ9dmxWjVTNJ23weWjkijozFFaCWCqTpUU92Wz6CsUUef6KSk
1IiGFVbq/l8OxufcWTrSucf3sn6YdY2j4eh9+SZR/CzdPKZUSWUUKWhGa+qT
tfqntaq/TGTqf5pAxAmn5FE3CiQkmXQZ1eID8OdJt//x5xSJU+/AsFngTeHf
Z/QxZ4o3t9KNGrExLP0Kehnr0R7fRR4JeKMlv09B7r9e3WMGLlFPTXI9AorM
TZR7uVzc0pFdX9HBoUzXh8ePJxV9P+DkB2Xa9+lf210fG4B+T8YNq5c6Yrxs
SfKpTGD7xAZ17LFsBLe3VnWTiZez2y0A9rVjelIym8FUn5VWNCCtkfOkl/oA
WbJVd8ufyplAdmARZUBmwbnU7JKtOatMpPMmOLRAp3aY0kI21dPnGIK8rUAk
ZMV/CH4J7AUHZszYI4U+wEB2C4QNvzbiH3mAH1C6NmPeEnPj/+HDiujY6CN7
h/XnZePonDDpJpOq0dL+ykHT1M+OmWndOdyEj2IfTt6ayqwbDLfyRDZTSInZ
yIFBqU5cgsFpk3CkBiAG0Uz+iwrB+/B+XD5yS+y1XBSMXDwDeca13wYc4h22
zBmbd5yXy1YoeTcS22biXrqkTTqh2Id4BMVMPkGIN5XkfA1WxosD8S0yp9Sv
QZbKucEaaYamhgsCd/0yD9IYEuHGh9gPk6hGkrDpVssUhJWBYA4xY3/BrCiy
XsaoXQlFU8QuofkztK62LBlGyO8STyNA7H1lWyhe2dilfooac80Lzne8919I
EyB32SJpGamaOPrEH7YHd+jFUTfK18wGdgRJuElqPLuW4h6a07eWkzFa85WS
Lz/9E7MWIJt4qMZxDTljEovAyvp9cx36UOQsGCua7RSA0zh9+G2roxGY/7iZ
5d9EieOD6Ylk4muva8/KhrZDQSUd0Mz0eZA/xH7SbxVdQuGJVd3Qkb6J9i/a
merKewwH0DtQdbajjOGRseZ7QQ6lWS6wt46V6pP9dVvVVhVfarraL7KtkEo9
iiD66GrkvxxDi9hGrGEG3HP34KVYSK4eTYgwvAgTJFHvIDTYTkQ0g+PUKNT3
s+5qdbKg+Q2F16IxzGfJUJsDSWTVbuIzf/srW2xCQa3GSsG5aabT6zhlDZMI
+NBDfXV7sRIsGxCABYJbtl1ieufbWP+/hRF5libVWStwDhOS8ncL90EOeQBI
f7Iap9ftYuZHvzYALACDpCGM/A9nblF7srj5Z11I4XYrINcQOa73XGYVuvNA
h3n8AClqcLrjMHhRDxyeoZMsnSHBMa9EngMIPBkwXpCbr6nx8qDS2rBtXhJr
TQp5F82eLxTZJaLP7zXsetLqv3jKtnR6ygeIJtK7Hbw+EHvPEmdVDlk2HmZc
m88BzCUBRByBvKncO9gjbXUSptCqnq5LrLivO4BPHuL98TzcVjJUmzxOPtsJ
MZo/1vyhNdV74DNt6C7fcXpqDZXMlUcw4VySIcAliO1bmpw1wMe3u+KwCXr/
81mgcVuunViDvLfWgzkvGCyZRFPiMQgs65v9PDF8yMpXYS7Gyl4QI+rn4xng
wXWe2reMupS+4HIokDMbc5U6eTG0Af9a7crY3BKXXL2oPHYMd7lWDhWF2t2n
iVsGhteUnNICXAQbUfQux7cJiNympv37aAUVBQjpeyiPdT/pjEFT6TMlihVt
XH/z2t1+O4NCRGwzow+2QD9CU34PM/MqEvw+IWNbnl6BRm5gXC3DJx65ZyHa
+w8fTVW90OG28QobcYEQT2D1bKmhcyGKvLeBa7W2RTaerQts36fQt7f2xpy2
LOazdN+81lq+Ad5e5c+bNR0DdEKgOtHmqKZTRpkvqo1LnBWOF8ztuxWKOOCB
Qmgn4m54/pStDG8zJ4yZV4CPCw7FGoM4wpTkllabzaC/So0m+KfoiVhPi839
c/y20Cfsu8/Jt1kUj1V/KP+HDtQ0AYJly4GfuWWbk/KEbz5ymTzqclsu3+hn
389ZOXYbadeDNjbhLAqkqSpjd8gGXtkdvpwpLcMd4wnEHWShRj3Py876Kr6K
7aBHiG54b/q5QZIlnn0ARRDHpClFDO+aF0duYcSz2LDwIIpmHRvJuyMxKYZv
ET/gk3AO3tj9sfHl1PPfGcQcwfXa3SDqoWY1cNQp3N0JI7HxsF9fKvh68whS
GLIeHt3hWXpfo3nOSHiiURrD1Q7VCIFr34wTNjlcKqclCQyKsR7H4g8ujC3H
JBaRfEKljiznL/4H4KInQDFr4wZUu3ShBuoxUnQS0CAbra8Q0GbhUwOJWleX
kHxUee5TsUsJ6uYiR48am1HbcH6L6mGLG0Nvbwmda5T4lKOGAHgINxA1NaUP
XQl5vXJZjlR+Ga7Jy7LIwd7GUe9fH/a3jj6SO8sKhOQZqhivoncXafinNdrM
9o/y9mMzsY6Y5QxIdn1GCVMQzbf158pNRTkXXh+LsN/WC3gxYqfZVLHwMhgw
2WYApNKJCbr8GCds7KUWG86NGHYyJDXVyyRkcOpCeHvrcbdh10jOq+k/J2Qp
Y3bC8Pkn0M0gHvmk4arftjYOgqsgKqUUsoh0ts1bZHMhwsf1FY4KJgC1rKfA
nzrT2O7jNxQ4/wkBPQBAessN4Z2oZKAhznLdEEsrjbJ6JxgKBEXfliBZBBcL
mW6oFMf5Ae1MeF4eGCpGjlkxlFr6oeV6cI/ZO+2cs2C2AZSJo6SJJ8jYYlQV
VxP+ZY0YicCSAvPjOgZXN5+mpqmo3mItEIdTU9Bn7o44hWHagtM+6S5iZBmX
hX5f9cmfl1CRwqJXl569y+jUKRENf9xAvoMyT4qAk9mWQzhrK8U7B9mqoVFQ
GK5vH9rFGz1FRC9x72C7DguJOHGMag2W6NTjp3Uj9vRIYjbrfXqM34SgbOvQ
/76idA4NmqBXNBxzFjdrd8ZyQU/xlku0mM3Trde/B0P9rgAZgfkdlCSPgfA0
nyYJcwRuKNTF0tp2JNQcq3WuZ5YcZ/y2xZkztjQBZqBNaE1UqQB56xGDw26o
RqjCyUBSdOTMUrPjjEi88Us3dDrIpOYbeVwfET1htrk3jTnQZjJ7iUd0PYKJ
yhJPUSk2crKzQ8Sg7ZoU+Yqgwc6uXwVO2KeNi3IgpfHUZEc9FgTZWc7EFVhz
1NvMhCSQSdnooTJ2hnZshfq8LrlrX9U1/Z57jjMLxoHemAlL1XEwMV6hMxay
SGes/XnbcIkXoqQuP6EoZ1UZ6KflpCeyqBVV8i3NCGLf2a4sXNZC4ZMUzQBe
gMW/QM0wT2s+b8Ot/Ti8zrmjlwaZg6m5HvOgpMnfy9GuSZtHPV7eRh6wknoX
m3dFfOrMCNl3uAkFSCyrc3FSGilGVw8fFRZyBl1hcakCyyp425miu0trE3fB
ZhyNQlyLJcQS6Zf1BdIIKAdCZAO7/G8LPkrNjn6GUIUnGoOhXNRdusR7oToP
3rN/Urzft/dZr5bnI6BELJf+U/OYKL9w//zc0mbKlUtFNNGUjiUMaGHpyMLU
fRhbiVtGUoN7ACkMGcvBc82RjmOfhH4ImJaYrZamrZF6HJ4+4oja1ogjQvxF
+tgEPtJPRiuqtRM925BB91RIjgSLV2sMDqoajRjsQrk0eySFcsD0fDR88MfD
6nuuSihsenDYV/97GHjzFyrKa9+k3jTGgyIsblJ+APgcXWyVvLlEnohuPdCm
nxBMmIgSm9GxwIfP/lhnjeOegkyx64I3t8xmxk8zYIxi3df+TQh1Qz9tRdrM
SaQTvIxHvRHFTY3Tl5UAZm6VyuAUI2ANqq+yoAS4G3Ukl2kTO2oPg9exRFce
td3hxYZ4AqRz4ykutT3l5duCD1paXjrPtAYTPW4vK5P3vo0oriR5UOkKnK6y
hb1goMTtT0HNntilOtSO2j0kskaMX/0xINWV8KyEGXpHJ/+SVUWSy9oP1DM5
9ApKkBZdj14qRK17/VRhMc3EqPmHCqn/CihBt7wiWSlLyEKA1SHt/ttKd7ZD
uc2UqoEjRXoI8o+g1p4cHqI/XWQriWs5ARJe5ZWjLiTeaQqqWsPoPuobW1aE
6yYVB3ESYH9uHS/f5djHtW4iQY9FoiQ5AIUTII/Lpjz5+eFexHXOMd+KI9yX
5oFe/UnC2o5OKtCZZ46byTs8HKgZ3kUCw6E6+rFW00gYKjd8Cbnt2dYaaCmY
HZn5f3QZWolvJ/GoqTXhq63mm5IYcOtd9LGADYfWpSVuglnTaa0dNwLXWUFO
DWVLiqH5oFocWdWLchE2VCExz4rpDLn3UtPst6dr4mkmTannaVdkc5Nsmqj0
QYCSffhB2tB0FdhUsGUdm4TTqPCoFchEO0sUZTdoFGueqvVRAffWsbYQbb00
19p0qoaP/dpCtfH4LZZII6HZZZH4ni+RFCLjVtFWlm+1I8vZlrwL25nc3FjW
9R8hwUL+01Ott5yDPEiP/bzL+eFQefDb2cuJlQ1eDSt7KZ/of/kSDbEH6o5V
q5hteZsPsSRY/QnfMH6oxu2ZKu2wGgad/SoqD48IMohaUWMMM5TwBfnG8Ywv
ubPG/yaXZRV6hV51tbPKhoxgE4VMOxUYVCiuG8i1976wq4If87T32OqT3/mP
wJyjXYnPOebKAvehLyJBCJBDeJrBMhVwHVKwC7JPGPQ3RT5waugCQl4vPLmQ
bQ/AvyGP5GA3QQmiEm9qGWdlA+mIjh26inznNXIiXbENH9O162YHKbCk9Ex6
v6QJ0YT854BwNI6or6pidFE02tATw7QPH433Q+6R1ioifAucQ0rt+/nDw1Qj
1I8yUz2DAi3/1ZQmiymCyd56dKtMp5TtTyDOm4J8ZP4qmUQO7cJMIkW87pVX
dtspcsVsYYbs7ZZUnn1vDgk5FZy1L3zwkY0WdUYJ8gJuzX6tdWLr66zOBglE
sgjF8FlnCovWxyGmxnp/L+dM0JM/DmYgCKRZEZzEFkKUup4Map6tweQUKjsr
s2abUXf6kY8nd7ER2Mpkl4GIJbXxkgaae6zkJu4wF1APkN+S23VMz1xLxM+s
oPcxlI1O0U4finEmylCU5IWR//GyjSPP5q/n1pOtP7AK76R+q4dcBdqLomxD
wfQzNTQpDQkl0xr3w3PMZI/cuPzCGQSqwk/IETG+LtAqqE9I4Y2UWgviTXlZ
19StUF8VioL9h+1QYovbYzUuJvnEG2v9Ogu7jnVnqbRAP46YtMP2avBFTM9/
qVaW9ftnASjmBKC1GUjjz5iLq57XqWUdJe4B7ANE4ubW40YlNLxAn2wGN99M
6212huJDlMpSgAX30ABhG5o3OSAO47c9l9RH65bqHkvD1B0T+V6KfuhaAA1d
k7B88Cf+NNiY0OMCEvltOZbJlBd8ngQl8m5b18vs4Y+WX5yBq5MTAxHuNmsq
rKtOYU7xFy0RQYTTcEuZo1z+egH4TAZYGRhGwJ3jCmE9qIuzYby/3oljm+ZG
v81b8E11UkU07I08s1YwI2WJc2aODmxMnO2KpS7w/TkjeQQ+4330MANn1DRL
zGReQnxUdiM9cnS/kdwuuZuUNho5HFLMwgVrM7gJiBSnhMEuY5fQdQCy9tHp
Gi9g3meZUghvqfjJta1IUjR4J8l5Jt2Z7Hifw3faMLONEvGRFEijVmku6vZn
cmHx3haqIWJ2+0e/mAjK78DXn2kovqoIO+OtgQSIuH9cm7gMsC1GujHTWf7L
gHF5ZI39bdlBFHUUXdhbq11O9U9MEzj7L/g7EqD4J/xKozhN4YQq1/n5ZJTj
Vm71FbpQqmpPufgJ0mudTssEP/GFqE+mg8o4nKyWPMFyrP4HicCZsVWFWFTg
sJ9APiV5bqq7JF78GczMUMGQvqhlFWgj6p+8OcN7owe8KZtJieZlFhwF233+
zmaZeX6J9Hy5c+Ib+VYmCUew/R9Bpyq47Mml6TL/2z5oeSwl5KLQteyv+O3e
NzlsJxINVtkp5p1h+j4DQ9Yzg+OAMlPX8xZnEz9InYYRAX+PPein2bxkF/tg
oQ/pTIPEMbnu2er19g3Wd2IegyoN/fqKPS3WqrLQ8N8qqJdopgVfK6MAb3wn
f/vS0yATmf3Mm4eZiLD1ACMLMEI45DJQCU6Fnnp0Lk/roRNVOVAr9QSY1cyA
xqOQKcScxn0Uts5Y12wtEfMBMGBhk3IBfJEW3xZiP0OoXRvdGAdVaLZcGxe2
Bbr4nNVJBwN/SY+vxI/vLmW5gOjXuJmWZJTHQFA9IvjOeELpNSZ79ZMvuVd8
pY3Pc9XMdDseDNikrxZ45n7k3x7A+hzgIGR8N8B0F8xYXrJMp7/gxedeacFp
WXDInD1dn+Ev6rCI3isCVjaK0zU2GfwLBjfTWouBh0qy8DuuwV0xDnJ3umV+
P/ohNqnJ5/EBzP4CZgveicVawwOXcgJBomv4hn8TUYckaFfWfWsiUwxHVf1h
7Ee0n1+83FoUlDiQ1QetwaKPF94Sf9nU+Diyi+NHpzHTlkGy6VM0RxxwXiGA
JqYovYsn2iILVhMyQ+Ajd7BdXQdI3m82CdkXUm3UcI9Xcm9p3awDE9J2EJSL
l6xo4DcV0TN61aA6ZLeQdBa6zz1PIUxtd8w6iSsl5+YGTZMmr6Xl/oKh7mLW
qZ8p5FWmjU/02Ub/opOHjAPcVjQX0CcBTaTC/BiPDF7U4rsikWpFMf4GdkUQ
b0m5T5FsTZifaOJ39w0vamylOg57dQTOzDskT/iZcS8e4/YrY1Ao/r9XXGV/
Ww5pxBeXY0MWz9H2enWLkqsauq+me48/pDXZ6sFcmelxUBaA/3j9p4U9oegS
qTU8OVdSPwNliKEoLfZBL9Zl6csQHk1dykNHbfR7qKew+m2g/EoRYGaQNHI/
3kF0NIOXS2Lkz9WSiWQmKtreZ1TkaE1CbMp7gev5tZMJyoXxNNj4/IlNz9ST
Hel3P0FcrU8Xl5tJl0dIxnfEnGcP8wunoRpgO74FhEKn9QRF8oQDX/xIsIkp
KM8idFHDpZF80vBkuYqrE16wYb0+43XJUiVBGXooAua0uwGmacuNsfBobHXy
3VY9w6Gn13rkdNTL4fFna8+gLZDoTrIeZFuMjUjbUXF2otkU0/nKoDpEN/tL
8E7NarGT65TTGN6DwJkbB4KLUeUQ+3yodXZuf/GvfBLI2nYtqznVMekzYH+q
9ul5LPCQRDK9NDFD+WhQ2VmbQo11Hcm3cKRkUY+K9DbzFbX5GVja7QviuAtG
eP/svGuwP7bFjo6xh7Cl1eWDx0vEjvQNbDVp9IQKoFehqw0fFeKgHDXwSXfh
4bS/O5yIi9b7JBAztCXz2lYsaqIABPiwhKIEbhRTdSlcN9GmfJKEACug888h
97GzV3GbLx7VcAUx7m6U0OE+ADAI2+Nq8Xims/XLT3E2/33YCvbfaWuUkZQq
GjAUGrl4rPJCnPoNojxGrJyglcpnhknKuG1LZirn19efMcQ2bFyinPfTZ4/E
lyg0U8pb9I/nIOCFqhAMcVPaYkR2tJb+JlQUCAkqYc5W28nvHY0R4GGUCxvs
kC+fWsKVuGkQ5hr1Au2PibjzTZOqmdf6TPweCnOIinmzzd8/epmU+NzWTHCm
sP3t9JNFoQkwF/63gztOuUf8HEX5InGxEhNzv5k/qgaVhN3mfkF4d/8PpeY7
fl0jriERSZl3Qz5nn2zjbckyN8CTNFRDR6AWaotwYYUDgmR13+oImNZPzz6/
rMZUOqaN5kYfxUXd9qJT7mGlYcj+l8f0jVOs4jhYY36y/ARg+Is94Q+Iq2+S
oQflm+8u4b2ydlRU/0/YdwhoClYbB9EwLAYeE1UuPK/2ajTc9h3mS5EIXSsZ
TK7ZT84dKHPFHsT+mmRrTUj8OkEUXZ5pK2Ef3wBBF8LpRT9b7UfVrt629o9/
ci71zAM/VZ9yD0CZelafsTpbtHi/ttLVM01trGZXUhYGVCQR8X0UJ+AYO/gP
1D8oiSnjJ32/HPsWevfCTJxorxdLpPlhe0KsBlYTyX+kiK8+lHToU8cGlhJW
V9pVO3h5TSs7oNhs5spE4vQqw0bYPG4Gv58EWX0XkVjwlpw/7alOL8aMEvwI
Sizd/btEcHFCWGefWFscOVSC69TrY92bb/S8MU4Na3ecJeiu8pUDyW8cCXmt
TP27S514Yr0IeN5XZ45Gg9xXyerccnaxmI3BuJXbfpDAMLcs5/UplpfDEjPj
Rbuodbjx56f9cb/pmcjlWgKu1cpMmr8iKdIiqcZ3vE/1PYSv6/IlaQ2/G1wj
fxJ6zuGsaKeBOF6apeJD+CBrmrIa5HkEAfslIWE3y2k9lTyAAweKe9luv+U5
ha2msK8Kijtvp018m08mH/xnqI6/TNIJpSHW69TMztcZ95/yS/RHz2x3EaQ/
O0foiOAZVzKC7KmDapb3Zcx6ynsURHz3p3X24zmVYFifSEzL0unCGiSvSbxF
pGzqjgvuoV4VpFXG+yb2eIFJJBm4XGRLA3sBpmm09B8WpKL6X8sOoX4HLVSA
U3j+iSexBBiulQz2tig4n48ye7XfYrZpV5l111n5mSGcc18TaEXlJu7M2g5/
5TOurUyaHur4rD+pMjggm/sMrKohWlq9vbKlEEe6mAjBp1f6fUTxBbfd/fi7
j9X6yfDGUifLR6U9GPd4tsY9uJjtxD1K7/b86qD672gv1dOuPe41ZXo91udy
xfam1MCY4M2iWcCjWYUvra/KkBrXfaYBDW41RXh8aTqKuayTPf6PJaeflkKq
nA/MAScoPxnCKo1UfMNoG3abKcMKexvsAq4qFr+UV+ar6LfOU4gWh28le/3h
rGPkMNVJvX9p2LuftG3IpjtgOjfNDcUXxJ3Y0qoCZc7XCMHDNWEebVd9zwHX
Ssjy+e9z/0NT6DxALS2mygh486zkNrmxvu4GvJ2n6sL32QjztVCDEPHxB+Q4
tgcTVWlBxn6UVKthmwdfTCKqogsFt/UO6hpLqNg/pfpZTjgutI+DiwMD1Sg1
6QYRFFmLyvwFWN9rQlKKyXpcJkBFG4tKpqDd0SQiksDfnqBCoPI/VUY/Gt40
VaDpjG9srKFU8YKofAMsSHUVYLGZAKuDj6dwIETzymadD1ZRzrdMDrR+DetX
AMOwRiefyAwynyYtYoGpYPfPpuAhEsJFBbLtIrIVhRci4rhf96Ks6H3PSDsX
wG9VlpPpWlZYYkqNr6pLPXrHEhTYpHNRJF4I04lVk3Nid19q0pyHyd+0mGDv
pQcKHO4DPtwEOW9mNyhXES0+JL886vCB9EbrKewA0i9aS8qJ4lBldenGw0lm
v51hhNBxDadY+V6jUVHRRKNQg6Z7XO8gSwBUNH3HX/FM1dD/18czAY9OtPHE
dbyLVFJnKqe4hPrObYcnSYHjCV4maZTUhKsP+DiONulYLUIwbSSfSem6tleX
pZU6+rQ8abgN9VDLjT/Bq1LNTcqrDXNlcvN2224yZ9bOsmmCjawpUHzzaZiJ
+Mwdk7yXOhKlgFCgOnGwQjAN44hMi9yQGxDsprfGPI2jVy4ABFOqfkfK0sKO
bvYydSHpFoXpgCx/ZRQ9lx68UquEsVs1P/qkDQrTflILmPx/5ErUG/8YcBZl
mG0xSkhYM7f1n1z1yK6Yf7unkUz9JL7Lux6XPYju0kkTwPCuYza3ZzO6ICu9
n5UkbOIBf74KxXbJcDZrW2U5GX+X6q0U6QXap1mJGat6oM7h2za+TrgYU6uc
d+68wrPS+v9hsQ4KSzpS485+nzJPUP1s01B8fZo5YyaOP9cJc22UiOR8/dJ+
GunXIiURN5OFGbNfx/tTOtEubPAMHN6BQsXo1IO2gRqGp4PfL0247AJHko2g
KAx+lJ974doWGZghB0+k5jOX8x7Xzyv+zdzQvLu3R3GgfA9gUToYvN/2FkBn
KKfVIk44xHR7QPn1fpniC7S32z6TJSdPbzZk9AtDTpMRYhdd55GdkWJdrNpU
/cWtfadDtLpf4/qJw8k3zL17aLdHT1a7/7+h1hxJKKoLU4OrHZV1F4pnTHpw
2yrQOISEDlWN9LstA27NzBhWPam0wde/N89FLoN+6ab0JlAzxBkavmfr0GRR
hOLbUfP+kbUHNlFKIcTp9VFT9/BMwJ6PgUgCs9yd/8cWPCda7Z7uU9e9k1fD
Xfyv53vrbeBt71fzllf0EbQHXWmKGpKIW5Bp2c8tCXNLLQ5MseP3GacvsjbB
3qA4itaRFH5/16mh4zvUM1tNpDqOYs/0KIVDAZDurORanLIKjCSeeATD7yg9
zTWFQgs+9wB4OoA0Q3Ri0gJ4Jd3+jYIqGf+zjPAaJ60ckdV3FsiVxD/CVvlo
xxCrauj5M0TbKnU+tX76qBsrJhC+WPphFIyI9a8LlRtnp5iRCoNbxyNls4Em
X7OukVUF2w3MVPg4k35cpxANMM4ZLhfhSr9+NoEoN/p5pf7ewNRGqavhwXdX
F/aCFXrRhq9KjCMbhIHRAp6WJP6SpXWHuD8DZzuk+ruYTXobXRV92Apf2WzD
9+ocxYWr6nWRAewA8pJFuuC7DP9gIhpdXai303t32Tpu/AGYBp1VWeCy2fva
mdElYToaa1f4adplNosOapNnsYS6bLzd+92DHMQVtOfXQDuEtyxWshpZAn22
nEdlkAplIO3PmgMbUinEDolMf3N/cZkrqfNZV11yEqx+5i8lnyIBR0zCsdhF
bZKgrtZdYR5RLGCYmpg1GZ0RprPfWOVHerPSndtNB+i+At0Zu5zLiMk2UWYK
Im/iX1kduoEQF/scNztbidAJtPcI3OErPihXKdRxQ/g6ZjqbYu7BJ4AUuqiv
OxFTbHM1JDl6u3ueaMURFYJJvWn8l8ggeDqbn9xnMykXfcNtjADhvmcCYGxb
Pf9lbx8ImbXl0XHoec9PjRA2XptRwN48xyzdo2uEzccOVXedHldbBTfp6Xrw
xuuZBlpAXVQeU6klFyHV2E01FI9d+tjS7wTNmI3oWESojCVD9aQ11JymAR34
lYXufaQpwIz6Z5xQdFGsWjjZwmg6mEpxUDJXJqtCYuVX1MIGpjOx3jJdzozb
PojyRJ/5favVq93JGBgOGzY7dd2NarHHRKnaUHMuhOHS9Zt6pRbkHD2aY3H8
2acbh/EN/I39+S2hYbQhaqhBWIgQN3NpOlReBe1lDMXqz/GOnS6J6NuXM0C7
Zt6nULYSTfqPHZtqC9FaJPyBr2VUeQessN9o+IgZeR+fnYs+oC9nGV3ffz3z
Tv6KgY6Bl1qwn0kmVj95WdkneyYolQPfBRx2hKdYJcq0fS1cJh8Ln82fLD8r
BjzjskyBuEmYifOwES/4ymqGZw4OEQKFaZ6O7yj9Ef0EJ0+igjyPoT4yjkTo
G+kju/oYQ6IubNZsF0xkQ3FBeKiqtk8nmBxAKnaRrdU15HWnmYwaaaI7Jriu
jzSZG1ZoRU9R4OdDJ0tdsNOUJMpkwZk8t9GswLwt1E4QDvSNP51FRjOPNskd
KmfakWiBlawBiM6M6+CxTM++pyUNaa1Et/N8drxLjWIEVLqAW74PKJ5j0Ep7
tv+V4ncyYyNrXso8RhhbEJGy2CmlKnjG9B00wOmbHCG8dQMkM9v9M4lgoiPQ
tmmGi3pL/JK2XV8iE5FXQxVzdV0UbNADcg5kBqRysX+IsVhovevx9rI112Dw
71yBirAxf8kO7ZUy47Xnv2yRSBAcPlGUWH9IJUwplE4yvX2OCRAjt6I3TRBo
FLZNqhAF6Cv1nRv+ADF5Wvu1n+iTcqWzzyJj9Wj1tmOT1K9VRQ+klBaOdBrP
DO2OEMCjyDGZ2t6mZwKJaHCAdAc4bCqGB/qx4H76jPVsX9nnaU81BNBTNIiU
zVt6S8C+x+YTpv/MNVBpKEDsspGpl+XqYjoxNvxpJiRCM7MaRM4pS8LSi/jg
g1qL26mPnThzPG37cHHztzRNDnNIGv0N3YsvdgCdd2UN5lkSzbL6VXsnNPK9
bg+48VRMyY4JoD8wb8zlvlxXwr1AQOrxGt3OUnm6Gysz4tc46FFq2h4DOsaP
r4W/zaxTIvo9ieRqUpB7HFOQgQT6Q94a+j2HuIsGcl53ASjl8ohXfEwS6sdS
/zZvr1Z5ggLgBG+ICM7nN1EH0tFLQ+iGY6rEqygiMG6lg8PU7XHwchzHxjeX
zPk6a1MxPzT+s+ctgHY+aaUd0xJkPkAzoaISxDCEumGB5/jWwQd+Ab+VL5oT
Y0ifiIedIeSoCR/MVo4WzR+8KCS5K1DSIZne/XzLXnC2ILtwmzF2mq7wBMDW
2wr6qwCso/NqQINPKXZjivCrS29nr4iSL9p5+AuxWiHy0xDHsCJ59F/WdQ+G
7bd9JLKgTxZ/b7wVL0M/M+l2K94DgjE3RWhnBFX5rIg9uNxj6sql9XHnVvB4
ZJLAU2dFTflG8j2kgHi89d4eznmo0db/FzLL94/nXsgXOBJr6eC5aCUVB83E
/IAuGyQ9v+lF7JFS6Qhh6JvKKY371Cw4Ynf5ioNrWFjTe5OAasxJMRHcycJ6
YysSJYcP++PAyR3OEVzkEsM3FHVz0CZb1uRqpVaXsNwXQCoeRuADYjBaXakQ
bB9xuU7Y9kdzFww5oeEayNMFvNdwFe7JhrZqWN7EjOQGS7pjeWx6T/MZk7tG
e4nr+9VKfdI3Pm2Jkgx+Q1hJGOP6tqglUwyi/0eEGAszD4G31U8XiPkB8H8z
IF2WpAMFIPgWoaYmb5tbsL0yFsSGildwIrYu9Cy3N4M8jqvAYoZ21Bopi4Be
uG2J1f9Uf17Omo7+LBS2JmqaLXixB2QL+UmcX8+rWigvVOgjlpyL7tUu1Qvw
5zdXoCvKJa4rRMv7rqzRdgzYhiVp92iEBQmAW/y9r3o9CGwZanxMI6B1ir5R
tyXvUQ0IsKMv02lohwpnaHNWbno/E5TJrF/qfHfhyCXdxdcLY3bFWDkiIfYj
rt2t209637hoyxe1hqbGHAHHXQp/p0WgeaFYZIbHPoi0qcLZlJDM4ztaYtu6
HfZKVkm7cC5w2fdyQtROa8/pe3GUuzCoTExBcQHXsst+UUexRwplEt/2tD67
W/Rgt96WjPBnaL/r3GL83DCHwDWBRuatd6IBlXkRJFh2JyEO0AIX57XLZ7rC
tgNjNQsqRqgccVtoVAHhCfhibkNXNYvM9lZ+yTPMI4MKaiVBZ4zFXw72OFi1
0iumftSKM+sfzgGZPCOT5aADLezCEm5oTqdbI9T4bMf1qgXAXabpVUd5Gmul
K0ME9IfTtRu3ZPYEbOeAByUWQMDWD9VV8t2xX2f/3u+Bqp5YiH+jGNGAZQOI
RE5f4Z4rEnalJEUWMPY+K52hhZrbDxv6rb8SxxKcXgFvEK2sJe6mvPQNRNit
iPFdZAU6dn0T5Owfvjymb27VA7THlcNQ0rDwyL//mQZe7znxM6H48j9vr1mu
zOk4CBOJ7wJuFKD8MuVMUO9+11lRXMjxm8REFMJ2vTJLc7M3LkpRfyJeibmp
0ycVhYOAEK1bb7yQLuamSUbLvz8Mey9V536WgD1nFEJwa4V+EfZQQ7iGx0uT
s5QXI4/EdmslY9mvB5Tg8NbdeYP0RIXCSSMlepOtLTpNUiuyxoGZuZPkdQxO
NB3jhj1yfOA6/ddlKntj/LkKh//SxeA+zks3GR9ZEtWOyqTRkCoY9Ph/zqnX
0AQlbS8CWKqEA8S1/QBC+qa9Y4/jpkAfTyvyoV7h6G3tD2ohuAHjewhLMrBM
mrcF9UftbfsrnQPi05jgWCm81qiDResDxOdBZqjT9fk1xYHNDDydN9JmFq2q
4uJhQxzCzrVtz77Qsw4iRj2B5SvUirzXlhZXHN1P6NfctLIWPIqwgvhdRj76
+yCX99L5mzZxAcFt/skR7rl82tQ/owC54Any/m580kdAJS/78dIJwHBlBwXU
tyYEs9Lz9bsJL7IHOWcf04y1D5DjJkip2iLF+MSKgqBctYuTk2Vfn+vePYpR
E19IZz7DeU7PWWVvLO2piGhEuvjyVgpMRw2Atjvm2jKltigiLI4nZD90OFXf
dGn79zWpEE5XG7g4Vk6AxYl3v2Pf657RZzvS1jh9YjbBG98uUNdoPzfjsfg+
Twtos2zhQxFZdsPLBroz7UbCpqXzjqL+Qx844l70zYrZaE6aKpd4NvhSuESh
S614ReOljm1sXLlrUIU+SLLea5kz9l7sdO5rdPE9cqjrMmJw4bctzSKHLPJY
GpEZQc80frnpRlZMe4/HcirHWNexhYEycAc3HCdhYWt0z2CXFzc7matOqV7h
BzF1SxAwh8VMp4bOnt5MFQAZ+U2Fvu6pZTFYLJ7XAuTlStR/SuAvHi0AOhKk
bBxXQYcJiFzJK1KkbTkxbFg5svqbCiWhFLTVqoPn8DUeaEJ5fGNiyB7hqjiD
zq2VnJ8xVgdrLYw2bATo9ylPIKViKBEw2Ao3TFtbRjpZihm0V5jrKEWzYNZC
a8CmASonpUt5nc59kyhZE8x4qUiu1TmDdd4A+5mXrn24A/6mBB2pU9NjfFwl
Albw74N+JmQy0HugZP7WtdwT3poJRjNCfDez0X7D8RM4ob07a5gLKj0piQ7t
T9mD1xG4MPmd773AraP0UZhVp2OrZ4y0QRQhNNQjNKpYWKHfx0mUaeM1piZI
/hGN70aazUAzLvCBRZIPjtr5FbT0zORj1K4WaOFe0qm7ikPzmzQp8Gq4Up3J
DifHMXMYhem+aBjJ2UjZnVqsWedyFVoDTt2d/g9hXW0cDoJxGBVKjUmR1qrx
2E5yWfDIUd6aSvmH3alzTzpaGRopzvQdnf6o1JWdQFJP/IfXSbmm4rCAIDfT
a/q6JYHBhjXhILnQqkNw9OxPnsBmRzyl3Dpx3VqifRksbDb/yPxA5aXISaTg
c5oOj2ryU/aXnqF/qbskLghlOyvitD7XXYqNS4CvFuAPvYav+mmvvTLxj6Sn
qadmkOvHlvEoBaPisNRoMjyS00R34bN02miLVvFxZY3gbzwCutu0NIJD97my
lOLCKlc+0fmc9hzWesVtZKyYS3pAg0K/DGxF7YUpHDnjnFko2T+aXxPouPLR
lwRSwM5Vv7Mh4O1tIyl3Qs9wr33EAuuNgxRE/gdG99umchlr3boCFlMIdQnq
KI1F7SjzNm5POmYxPjzf+vCEqOMpJKTEYDiiZjtA9g/Nt6RcgnswkGsVrc2f
MWHqiXGqzCmkoJ85A2cBdphVTVdBPdhDuIil8jr5XO5wt2mCa2GTdgwFxl+4
ppvxUcwTkxx6iwQFkQdW4Avnvj48dbpbZZGitI0SWxI4uGa3EPWXVZlFVmfy
PfFCnllAFJX2ZgtDfnrviA+bDe+TO8+QG7ymb5lGT6jhaEWlf7Uz1AbFmcFy
O3LEf/Irc9iSpM3tFVutgGvGM3QdJOqwZfYeG3X7da5m1YPLUIZlgxvy1aBH
aym006CL5xg5m0OivlCENTR01cqCqcHShkhVSKZz7qv26MjRex+ibClGolj/
lkMeGP3qGVi0XjV5qV5w9dAHd7Rejw59Tzx/phTpQ0G/zi9zthNi/gjMR3P2
sLSgqxNiSNc4BttSGP2NNWueGzNZuonxhibg3pn1Z1BRU576/aNGEqzVJ90Z
L0PMAh/2llQowh0wPcYYBEzWfGd2xNz0jqwLMxtaHnva+GENEz31Q+YqeJIz
/ZrVfAwmIwrmQHpE7mMgsNtL4XkS9h8/rxGVYz4wzl98gIL6c5YFo1gdmp9z
deVhrC4rmBg5dtjMP0nHWDQtkivFTBJ2+A5V9ZBQ1b4XtoPg+XjoUY17HJdV
6u/UT1n03GFb4nq36Ny91NunZsnvy1FLeWJrKnu4qIZY2anlVYD+oIEOdzmq
KW4VOoXbt4H7EHFS/bBcV9Nug9QyiT6yw3mkCVBiT9gKlhf4lVe8I280SMlD
lUS7ACNYHZUNmPZ3wQEIuLqNhlb/C1LonZ2QJY4L05Lk67CaMLQ5E6LW+e1t
qqRM4aLlQwEsDspIUO8OQIjC59wZmyD3WtoaFIS7fxBdswphPxKcNJdcmphR
fzraZd8KhC9bFlhzszg+Vno+rBdSEj6YnX6Xscq1cxYbYy4Xg4C93ryw8J+q
E0C0mLksgHDUG5Y83I3/bPo2GENWMuqvcfIBSwmdsk1erWvVZXOV1OtHTdeB
hRZwOZA3/pnghac82OnYux4dVJmxj61XG1fYR+po/irDNFJ+eI0y28/FXPUY
w9kqnveHS6SRKrjbZkZr5Bh12BW8JwCMR2l8u1wAlU0o0qE0piEcecpYtK2Z
koQ56B6m23jpvnMYQna3/lRsvq9FIewctRTGz2kgta7uLyK+IuPg4UURYQEz
ARNN9aGAv6fwC7rTjn2zOPGTVchWMj3+I5vE7pyYwbpGeQMnE5AnWX50xEgF
XICArRg+qGFjG3S4deTV7Z/n9vCpvOxoL9ytoXcFJp/zgRBBwsDFnqvCa/8Z
XQ06cmCyEtZM/U/TruN2Gp+0lxaFL+h63AUbTKKJQlYQSevYWSF0xoFOqms0
mTbnIjEpfTHO1nWyCzpSSzcAL/2hRaipTmQIv2DDPsYFu4vzs0MtZLx8mQFI
gaEF2PCgzKxTkTv1H47kYayv5ecTt29fh9scAH5Z2j3pdc9yMidd5m0FBo/c
Q4AkWQ5Kb/Kdr9oRLw8zntF/Bg8S2WJUOlHwtla+ae5yG2HVJwp3xo6qDSKa
794wUavik7zqQJVm75lI7z2KVI21fS1ZZALUS5EsIC0bxrTw5dTsFh6AvESJ
KJ0eDVz5M6Et58BxzIm12zHvbahcUnF46oLfbEqsjykP2bXZaE6S+/w3ZMV5
JnRNihbMM2c31i/h3QRLm9KPrCY+bMrlOFBx3HGkMXA6DLYvXiArJmAi3JQG
CvKTy+ysYfhdsmyU8nnX6P5ZTqb50xtPoXjeZWiozf/IaCrGeNVmSdCOH88E
gMzla3RibNC5Fr0sp6gtVPRsUnugYSv3vOiAkV1sNKxR5+mQgiWM0Wr3WVtk
IbdDlHwZQ9wb1WJV/+HL4wUs40iJ9/6SiT85moGSZGuj1BFXLrg9HNvOdazd
zYvCsqMAa2fh/xbolQXp6FGjD9zsIs2rnRrNboz9pnTgzQsz/hxxAKD4qgbc
LctLW0SYht5vwsqBj9DQqchuXuF212lC7RpPkGdLedoq4xIIO22Vw5Hjv2oB
ajGHLNvw6svDc7o93aJXBdTqoiu+sYgCIgRxCKx/Ivb4mSli9wzBNTp7pqPR
eZqDDeppACrbUdrI3tiej0bAhwbB3Vuqcb+bxKmhgb6A5JuV7PcMOGLsGGK5
ZHSagNMLvkMKJ+ZILB9sk1BkJUnyvADfJr2xxu2lUNjDWeI4jlfRuqVb2m9g
MgrYCCQUPKA3SaGGTryqh34CTGjrQptC2rTjZHXKM//V2j2epaIcjxdnE+Sa
OMUNcSgtXF8DHJHCCr+YeZw58a0Umyq+hJdxUpZ2vMNclIB08sLSIebYWbOt
jBgRP4WV11ec04GC2300uyfk3Vl6Jl56eUBDgvsIjHtc+LW9P/ygdQD7U78U
ZF1fq04ioN5jg6MxY03MRTiLzNt51DKH/kE1GBX8gF1CTqDLHHQTtLIgnI4I
VmT3bZPLc5OhaJjP0+6WpEmxdCr8/wBraCnw+Awhu6nNuqhmr+INJ+wkfxvj
VlTHBJElVWGIYHsnF8V3HbdMmmbZN3lQnjNFf+dsN9w7x7q/SV+eTW0HGbPh
45ZA7evX12roXScBob2X2wb6K0wdkbpm2n3Apj0JzQ0s2mxkMX1O9HRF+TZ8
gWHJyOwPIxTyOxpJhsPNRY5zkKTLHAxw9r6z6WtNZ9xXHaFrjoGcQcpuuLys
nQZWjVKcZnUQITQMSZNbsd1MAhSTId8VvYLoLFNlimBDWGfUr3RNsvIE/v4j
BrqQBUnFQIax0FOyOToCvRGF77kT7R5qcHXPCb9aZNDkPgCoGCharf+RcMqy
3qNH5bExKQvE65fK0gb295ekFbVP/WbDWdiAdjjMW3CFDuZ7axyWxIGB9hM0
gTuVvWUWhYVSSKHCQw379jJSYXzx/6kPq+GhTDwSTd/MEnIwc5lW7QBxjqqM
nUduPgHXK10MMY4gPDmFbYSoC/tpA39ICarsTWuQhViyNZ0CM+LEHs392CmO
0gqk4y6PVUm1Rd3xIF7k2S7Km9uC0ivh7cj6r3Fthc+UuBtmSHfvu2y0YwZs
AKXBHhX1yFWUFGdftP2lr6MBmWcWYdeOIxCzNeVQaSv1Ifq8hEFlZfsbni4L
5bL6TzInOC91P3Yy6Z/rt3dXBiDkSkXc3vgrOzaOeNW/6r3V58XKb8DYNfJW
Jk6+hyvTU9wlbfPMrPGxPu3ym9Mb4Dt50E+OnxwM91U/00M777PI1JJjxPPI
LkZagHdziJCfePZB3hOjXMPl4hImwI71ruJEuwER6QUKSCNjV6xyAVnn8YMv
YiBdlUFpGcjJOW2cuA7fPFMEMXrmxt9vj1evrgsGViGcafTnZGa9ZGjUiktE
1wdK70t3Yug/XBtlqPV6K4oiTlSAinwQboTfd2r3cfRpkjDa/dSizeR9+WEX
ISkeFQxW95sKfEG2l++lPwJbYvR6WjRUeuK1V+mmbe5Du0No6XLiDlRDsrCz
04lBM2qkWAJA1a0wGki6qlDFfYj7CoWS46uZ62dLQyIedSBPwEQDs/cJbqHu
OObM6LqkcWbiQh/kOsEwzXQIWY41FUtfEBTLQcHSIlMGJSouix3QHQaTAaV4
a+gBzn+L7PCclqH27+nq1ySpJuwK9ryuzU08sTJawY/Tx4ONwdIghIH23NKj
u58JpyyuKEWU3xf4PFmVwxqRkOOSMgmxm3n+Y/QV72CzajxxXDICPwno1mW8
sjXiEj72G5svVd0GRec/bbxHug3JMV4ZUo+MUPVJzoDCAYgFl4qjJvpq80AP
CtNRXXhaEjr/xJ9RUGUFKWIZAn92ceGfdFlu//qmTPPIdoLuGokz2uL14iQk
bogCNsT40+yF/NMxz7Tq0DaQaNuU8ZvsM+UMQMOpubP7428wb3EjWDwEPT4i
u+YjrMnoPzxUbimCMhjJY0J/nxg2nwtDvCYEeabLNKlwb05e+0o8ZeIztEfp
qC18K9z1Acxul2x9EJv0EWyLICZm3oe/u0Yx7oqTX6HwjFSmMWzxBzPMfIf0
keOqTBmJ6qkQEB7Jk670s/cyOne0MjlFnizXYElmWeNRty63VN8dmDLg4h4s
Y1buROTehcTUJg/XAs/oBy3rDk1HmEZuvPZ/xYIggeXCq3EkHmS054HZIliW
mOqh94UmwqYTPDMfxhLSUIOkmT4cmQPu2V33bL7S73c0ctNCik4lJ1VHikWz
mfDM+AHK9gIGEuwlPfxZGtpLNbehK9w8DRxrq22/VshEKrC+SJP1duX3lWI3
AIVZgZUPRHic2InOlm0iYwgL8GNhDKYk8l6O7wOWHgiHa6/imKrby3rO4E3z
YSmps8Esgcaw8c2DZ+NqIf91isSfFxOcePY3cAUUxEMuMiZh6+H/yJLkEEQ4
ZPs/nRYTFC9iKmMPC98qlY9+14yMZvd0P1W60IN4PXd+WUl2wJZYcLI8NoyM
frz5xaGuMudCsfrWmpS8fWdqWDg3vY/JWVUhmN7sgEfm5ZucRHcZ0hyyxWvU
iPOaS+E/rWD+07JlISiHR5SCGL//Map0vJDPTXB6oOfLXwMK+QSiKRQexkCl
cAugIJi4Ona31o+l04xyNZtG6AE4G9sXRQZl+X1y5l2/qzWn3erO9s7Km5pt
SPnpUlIlb5mOEvoBOdqn/IQWhREsCFD6itYJZLbct4TcocDzAp5d6bf6kljW
FNkyOjSTvrK8F0YUfq8iDgc39myFK6CIbYpWwBPIoUJovr1Or/BfjMCb2uhX
ggSKO+pZDY0rJQPJF/TS2OcemnUSiT0UCDVNjUb1IdQpFNTNqbNuFbLacINu
MRqbi+TQ3kCfHUJe+2GqwCYuEt/8cqDRMCSvALCp1npwqChZUgr4CbHzTye3
HBF5x2z1DsWraQhSMVj3ISU392lFA+ig3lpC8RSGCAxpCK9y8GpHywzOEE4U
MgcDMO6OSWUmNONvLhDWbNbtgKrCVqMvBi4ZRi8eIdDYYh+/9zI0fOwpGY+u
WQRIX7tQR4bJ5A2DpgcbIZAuU8lTBj+0i4U+ne6N8/Hfx2YaTdtylSNlaBbH
Y+lIGHcgl65jYKWg8hHcOrP1x17zz/U4wmtlolwd9/i2s0IeKwRPOjwOD28o
ryPS1zFuaEQc6uSMxhu5CDmVWbnc/JeLcQWshrhgFCdSbSXkq6nD3ez2nXSz
EUFh41pl/7Pl9TpMNz3W5EQx/ot0qZEi7lH+P/aO3E4rrAzmA+kCc78tdcZ1
fV5lP7ORzwoQXe61hc391erYF4KF7KgHbsF7cFA+A7OlFNvxFywymqOF8RKi
e+y2CRlog7RF9Fua1tkMumcGINgESDtRyQGOEQr5lExisIwk0LyVIzSvKSOc
SXknSA17rQ1yh4ah/Bc09VtI3f3lxOYPxD8Ded6eweDHBY3yfo1N5hOy0pyw
979LeRaZA6co1cb/axE3dtioubLwniVQ0t4190kl20sRC5WOpnv/q80ylCJo
qqdlo/ayEHJ/FxhTMtqQyC8ojPYf0LWtMsJk69jltkd6WhHJwubVJ04Yo+q4
9dAWs+1pfScqSaVAkJ/fecNYVf3NdMnTOK2Gnwup6TeynN2Tv5drK3+Obihc
qTb2WvjvHV6mUPvs5A6pg8w4czozvx1uzm9Y6P/sM+3m/Y1OVd+Nhy3wTZK+
GlHxG/V29A9ETIO9yEBaqgKggvVvE6ISZlLTt7JKj+P1RT9yAl0Z4XnZB/SU
U16f6oHs8Tv7bpN61LsbCFBLEMGIem1ev6d8U3nvEXA6ojksjaiIF1J2cuKu
dWP46pxdJSLws4x2H3hLUgk34kYbeZPj8eli/c2EGoezciIYYaz7CxkHk8oI
P46wed91Cg82BNdGQL637CqfHbSatAJIOWfR4StgLX2JBnrjBxjmQYY55PCR
cxUsPx/2dbtFSIjBDDg6ujAGJDeKR5u5CdjuMmpQHlflPi9m3eDpUNDzvfXR
4XFfFXpyWxkYaXBTtcfAJ+S2ARh5QBtW1kg44Psmeb9SrkIKaAIdXXmpClyb
VrdLxWlsW+JWz3w7/UsdoCvQajZMkcNzTVAnDpwlzpBu28ZxKDOhVi1aoSIp
HxlDyH2anSJfsTafBo1WBCu7x8QGKkAn5ZIRZYs06wYS2SJvFnmYYvA8MsWv
Zd9DjpYPHzgWYpNvxYMhDnNEVTfsCvGkCK4FCxgbC8YBrfBprM0FV4GYoY9z
Sb9zmiJ0yVSK7+2nDIHc6njtfY9RirGFH0B9xkiZkGw2G7yJfp2M/c1ECkJl
3b7EscJduv91/i/BLfZZ2kUS7lcvXH3EOA9I/U2/bnqUsnm3ckBlOhiuqWoY
7DGm4r+Tyi+I0s+pwoeehE0emGb6U83b7XdZHm4AdrMIT/S1Z95bWCfGp54U
lCbfansyluG2PCmnvSH7BukoHG7nJ74uTK2xDGgYUmjKPJjlPxCRwfq93yrA
EOrWGo4CtQ/ZYyVVYnOTM71GNQlSWw0RsfvEZzYdbzw8jTfwiZh/DMq1f2Am
aMyD5Zcuht/jj0/PIDZebpTizp0mpyu90gM7E3dHBuvAraDPa4vPjd68uAqv
8FMxAOYQxQmG0FRmpK/zAMLPYkIBpJ8zX9AUUT48jqaLi1IJG4e15Giu8oHq
REKaFIyEJ0/2irFXSpCDKz+CmFL2WNGloqGVtzGTfQwLfDNVBXsiUhwJVgr3
eFb9CRmYnCRXcy8dDbhW/vEWLaz8XVk9HjxVkJ4NBkKSRTBDl2LDCW7zdvqA
bO3VNSqy9ilbKad+ce97tank3Qfqd3hdlKdaqZ+m1HOQIqtPdGbkl/Uo2VZv
lL9wdEJo7DGE/Fb9y12xXogjm2XUN3nqk8gqxWeHZQ1sEX3eqJfhO0LmKob/
7KP9O6UZw5beHiYPwokrtcGM4Y0Phk9F+NPkf8z/3tbzqSTARc9VUbp4rOi2
tE+m0EJDW9xZbVz3YuzMjwZHDM+LpJPjXYB1vogAmmwOx3x4ULTK+5+gj/XT
j9hMttTFRVQIzoNM//gOkIZ00bpVz0LBomlDJnde7CNBdgD+A9sbehDsfzVk
WI4wFuY79JMFchn0LkPDZDYcCWNlAvjarXQEgTt9VUrTKhjM026dHN5Ulpog
tyrZSB5JO0xcaB4WtROHK0qWrur4BA2hXDq7G1zBwoUK2T58CUq1PDgQRuIC
jLqqn5TUFaTMYum1WOH2jFE74SCqwjCLCKf+i0j2oXOgjuGnMdtQWv8VCFTq
FAX0RTZroOmgQazdGFC7kfYzzkqjo/BvvJkVmbME9Kbkq8xu47yumYvyxLFQ
aQwqNO0ykmSULrWxpbX5fKKEkBMKgmhH7iFxb4hA7xFHiZTeEqPKpyVtX49r
b2cDOnQ/yfXtd64luxYXq/ppYWhTCxqeMDi1jEtstiuWfBjLN9vgaCEkxMcd
ymfjwX+4BFohg5fhaLF7mJrFw75b1GKxHeaJoxxEUaOOdXCYye0SyihU7S55
OLr4gNHZg1Q6a8E+QkwM3JJmOh03efhRsR22sc7QPVUXulCVxH007M5bGSu1
4e38tylHwaTlBCEK3Fb4C5ARCtKkaVzR27hjX2gsR2waNUKIVFl4j0hzku1U
t/4j0C0DROneddw0HoDUHzUsJ8xFTkshklEPakFO0tjd02bSEc89SVvzvxnw
ViY3WxfpmkcsUV1foBgHlSe9K3ay+grVrN8JA6di6Qzijk8FVGSt6Str/jSY
0HQBNon5QikyBmjZZRLfYMaTSnxfshzU3I8SoRg9P35sBYo5QVKrGPQJr02W
1mS13FElInV1TiSE8H+BKqpcOnuztCCnzGz/wPn+KWLRxq33jPn9sar21oDH
EYFnvTwAs3VUysi0fCCO/pz6LyrawFsjZBe6P1icczEMnVzDkm6oWldJN/OX
tSKIFir2x3/ga+tkDd9jRUPAU2FreoPDHEwdqydwj0zGNweiagvMje3u5j6h
6QNDwWITfrccw+Qo/YTomwwfhpU7P/Es/DDliUdi5nXYRgf64w9WJnhACy++
vHVyJrsvPZ+Xx0o5L4AJzi8vgcnkPkdTl6bqwe9gkPcX008QqzOhbJXqep0Z
YyhAnSXCbUIsXsE99NXG3pHoxNCfPGTbVfhZvSDoVmcn8zW0asF95aFz894K
+bTRLePGKmzchnnHTRPC8r/v2jqF1blHcgiR82E4wl/nOI4XO21NO9vjDpQc
jtVhR97OzM6EQ9jaCVMLopc1Nx3KWmpH6Ixd+qxwSG6rPZ65+xf8TWvEOj1M
//1pZgNZ7ml0U0b+JySpBO7fuveaaM/W1p41vcPP9tdsOk/Tl8fAmm2aYwAR
0LS4Aoock3fH4P5+6pn/VPbaE6iOdaDbddzgh/hL6crl05WR1RcbyPCtTIGb
7IyN8T8BBH5EHmz2TITPlnw7wNC1oh8hBs8JT0o1pd2BweWvyEQAqgsOBqPy
l5PLGpBMTZR4wCpgRMx6xZQ0nUIq62JYS+m0ndJQ1kofh5BIDl3bEXjt8Xzf
1kc5IShefgrZhaVN/j1CP3Qu5IfhXNAdcdhlJrw0oK7EXifzMgWOV1s2itAH
hlo4JM3XPuJDk++qBCLImws/UIRTBNXE25tvJkEQbrHMNUY9hkRMgmsW1YDB
XMihwIzHRbm2kp0QeKeK5mwVyQKmuh7Fd+p0fhqPx+sI0fiJW6UXMxMnbro0
/pCBcEq5zDRW1L/Z+0nFodIa32uJBLMxn4yllRF6QYNOWGmAqiJP8COrWnWo
DIlCASwag4l1tyA7UDCmoW+nyj6V2Jho8Upx704AdxFpr+Art3myjx61xu2Q
7+c6RExRvZIMyhxQg1OXBmQA+6SpVCwSLYneH7QwpobuZMzSdT0J/CUzmA1r
7PjA5zjjwVSMucgAm11wvwjLqclK+4U61S04aiDIqrbsNidk0tNzNTswzrfE
oZ2wevmlgPY5qmU28VOzosR2iCkfVM6cGbLlESkvg3ZnH6KM8/mHzJkVPoUs
KkwZyi1ZadPoeE+rpgFaCwd3IMpVw3li9jf9pORTs1/bdgiJ2BTPiUqALP3z
3lysOKqfAXNVrQxBCbGfPbSRJLp5SpzPrQGZEj8UQgcvlFpIPTLW5/MFwIQW
JsAHcJREAtcaeSs6bjbDOTEbe3yOQj/qqckdiPU8p9LtevR4ybbrn/fDCSlp
m6IcvQ62T0Rq45TPJO95vHxholn98ifCcg6zD8nj8qLu4YePpaTQerD0Arna
gj7Y2k8ICpetaGqhgOAVdEQ8V8i6WrRKw8wdfoNaqUXexWliaKc5dSujzWmR
js+LGoep+mAVJR44/IUQWGEYd1P4fcmBSkqKDLsHG/LxKO6FMpHQwhS1WOhY
EtWikeEfosmEDfoPYl2IYrnl9o7ZUqaihdOHmi//xYbyA4PpLa0kYpmjXi5I
HYpgUrPExpuuGDQfcXEPc0F4tB5UWIOF+QBH7cvkM249C44XUm+Iedq66vKA
k3KBK3ICHWHAgueUgY+kM5AgIBrORxwTjlvC1lJ2A5CbF4RqpHLhjLMx0kmJ
Ynr6ZqflLSMql7LJ4FrtSnABzDYXFEAw7MALOw+i1e3i5M5GDQsEBG2Qnegc
rZqG0G38zUC+N4pOVamuiWBLKZ/6KXq/ZG0vR+X9+RGVpgRbGUSv06EUObNk
fm6lGvMG9MD3s3KhXKylyZ78NYhqjBWIx8WSqRzaLwjswChNTPLEsUAOK6nX
T7f3Q5stSF025iHqoBTOQj4pqO1ZSL6pzBLe2FauY3w2TI90McKAs6F+NZRC
BmEeD/CjIsn0jsJ7rcK/Hw0cdw9N+fT3yrI8bOhd6WpOOWlPSNRqJTa2qieJ
0Pa1HBc0hCAYrhsOZgHVKdcT1fIR3A0okydG/yZbtILRVS7oZp2Qs4AEidvP
NbmVA9xOk4CpX3Dn+DF+RkAuB/2taZiGIIc4/PBwB+24IH8U61LBuxZqSbi1
8ujBLoumqGK9+G5Gq+n/6vCDOpdOndWx2h+gBkyq9Bo1wG3YunYpQP/+dbnS
tPa5G04ADCB6qScYm43SGTdlO/cGA1RDblpvIkt0/TSt0z+5rVOzhucP+33G
KJxYG7KiY9h0O1WDdJtAjkVGAaiSkIRVAKDmp706/5+ZW5sx3IgGmqPm7eof
k540xO0C6ie/KVBJKVRuEeyQ9Kwo93bAAck+DpeGreviDkuSbepD7v5+4UPj
8F6yDnCHOljef0oISr6VLfMNCfuQjXALm+Fhc9w6mbVPtdeTEkHZ4dYkz+bl
lzklanMQwAWj/UJ24paLiblcp1/n9cj5/1ImSVVxM3sjPQJ3UlLH74P5L/I3
ct17X9JXhqLO5fIAxMoJb2289ncd/YJwZvTfJ14fAEYOl3zuSo+Q8T0gB7dH
q15xiMbPxXoI5WQq08i+kr0GJ69BkQ2+PBIg5PVRz+C/hDkTrNBWka48yB/I
zs2vhy2ntyZG/T1sPfTIpfQvDAfKCWuHJ+dmALKutwYjp0GUh68gVI+fntoC
AjSstO1gnYRvnINgnyTjMeQ8FCrh088dXlrYYBTlYSWo+1wF4WD5Z4VHC96F
PAoSpAVQBDak4fER92rC1MSxKH/zaNvGKeIBVK0jHTo3y8YjKOt+vCi1cbyo
8+TyaVbwHM4ksVI8CD63WtMipy75lYwySf88NfeV9M1VPyJ548ezTOyFu1qz
bePwUtjhyhpIf56ncLRoWHfcD/7Ul2l3GZCLPIfUHd2UMlyDjkceVs/nbbFZ
WZ5+sNUgnOp40PO6pSPcRfsiLmMNkKSkGoZw4eSZZJvD7jAEsP8EgbSbfLtQ
spoavRfs0RiWAOi1DIFOr61gYxzSsAqpICSSXp1SQCs4YrP0WAkA89clj+nh
VvLnNZEXsge83cyFV2zR5aZy9QUoaSeV2C1RIuq5rbieGWe5f98tH14MttdA
8BA7uNPwMbmiF10DBVfDgZZwJ+yH8nN0PyUde683bY4PZNDR/QU3FZ4T9nXU
i6bF85BBwKy79mlsq0OYoxpTx86tLdBOc1cBya/W3yBnl7n4XflITEvEx300
aY2jMKsYPjw72jFIJC5uUXritLTKhdf/ar6ynkXX2zNd2Pzyl5p6wFgAL7uN
eCYuuvBAIz4Lzp/xP6zYMWYgrOnHAw6s2aeCYS3A1OhX7rttVfZ8UYNZQYkc
hUE+5XPdkupFIeI3gmstXbpHQQ98mfazEZUEWMUGuvCC5zYyX7rZkVZ/kerB
TBIq2Z7a2JhvyF6O3nTrEsdf7/wp67Ge1dlDqiP5TmlzHxBR15EOP7oksEQj
YIg/7MQunZKIIbgK2KD3zHjfcbtRtOhRF0EZOatuukJDbuoA24pzfwTjjYDN
ypR3jJb41BIc02TCWcPe8bzaghfGI9I5YmwM8jkjwDWFaWDljLsnLuyyUMkM
zYxIIkZs6F4wfF1An7zq5GSoUFz99aKNtNysSbVOb5gltG9SV5oMpdjL6lRM
luQrFmBFD2SW6gLS4uUl7BGHdPX6HMieV6lGqLRBlFO8ka7T+kzpMf1yxWwM
jDJHOFH9WAyBzkwIuzrhNqdSy25qDjum3Pk/mfoWspJ2Y89dFZIS/oMy70Fw
RXr46glhAY9i+Y4cxUCyimn7upC112lzzpawDWKGAX17MWdh/NJnjLHHVTbq
CYX8Beh5LFSPimC4DcPdXctysoD0jUNyQ++4QQh/fYx7JuEg2VVlGOW8mghy
R9LAabHu2ZXOKL2eGsJLnt6I3P4sM0p2i2LJvASvTKd6DXojT4zKcYAHHlR0
H5fRti1wn160XOWhGldGZcmllG/vHm01HZ6+v/BIzKlXGv0WlucqXcyVbaLg
le5ccQWBN6dsaOpTHmRqDMdki8mmP+RHe/iBeUddOQ3a1xzIif9wJChbQdbu
P+PCMYd6oQFfbSrsgQG9MrvyoWcoHT06vTCfAOJ6+OBGHmZvdOrPN0g8wrGS
b8yB+5J/PZDQZeadQGrRfEXFySFPu/yC+YDpzZn1Q+Ty2u7ypbYG2q5AMsiU
6YzcSC1EaopwFbr/8Qo0bhuPK7En5zPQvY06kZc0bwk2Fp7pCkD1EN1zsaAg
QqehcS0rpCedRYj4knWGlTuApjYbaWRqYVcy7uRjfsoJdeNEWBDJlOk+7zrW
4loHSzNo97eCmhH2aoMRI4tJjSieWKtwf7SEG8i6IVn0bRQucOCacrdOqdBr
uuNtN+bQCK8Ke5CfsEpTyBQ60IwdlNaWk3VMsrPKhFjRA5INCHpMHm0/bSf6
6IsYxQrGkzWpyoyRnWR4y9G3qDnzgWHOES8sMPf5h1mwW67zAzM8dh2D0jo3
rzXMPDBlCDtTfEcyaOzL3WtfaCFukeJ9Pkza8glHzdISOV90z03moc/yfLyj
E2nFpvVZXpHZMwLeh6RmFcgeImZz+YEGR2w+2uZfj+SzdoP4F366yVEdA2mH
UceKwg7yr9jgMY8CyetAWcExHap3MVMdbQZY7BLiigXm6a89VXHNdwBtzzb4
rakKQN8jQFkPaRIos4Ft8Uo6N+dM6obFIdLHFoc873MPURGNV5hXboSaZqsC
DUyKnm/ChdjcXjpPDG/SW8D5EBBMy043zhBMgckz68OA08ECO8JY2s8YknKN
z8THyRES0j0vXKj8gUAsRjYG5gsu+UQzJmwKHMcvXbfGXINVP9IZ/cuHRrTJ
RHDy2b6rtuobcRqeWwjxHFuz76i8Gj64jF7KMasfOVqEi6jf6cw2bO6f70hY
Acg1038ETjBJKXWO85s4o0+G/9qr6WNot28wIdp/01CtY3d/mZIUNytQT/HL
NGPfoAN8KX3m5gvkUqu1ZyeoYZCEh3s6Tma0G1yxvMom+XtZt/Ttgk7e0XV0
Fei26A4f4dBQOynPNo7rf6ULSJ82eZznxtwRtFGBnqgLIzLFYQtV8i/h1bjF
SYx674PxuWpW3g1tHGtnWzEkkrgZKd3ZSp2nLKNOqMpkrj8WABPF1gDH2WYW
184DaLKnQAaUcOGXpBighQRBG7kdjHh3/oDu8XVm0YXc/g8zGzuwvAUQ5o4i
s13fAXDFT8o+LFKCdwDD9rLhUNzTM4+Y+0yRK1IfONHUgxfZOB0JN33XasNz
HjcRrWVCdHxxUxNHnMVWcv6vQ1JxYQ0atwFvzfO8DVhrfwt38RFecW/5v97U
dsRPOkoBs2XVYxb9y2+CX/3goXotHrTukCXfa4QEwqEDR4UOiXk0Xl1m12g8
Aid82W/3zAMSE11xG2SyhmgAqjJW2VgD9RjLYtPxQqx3wd5Qghy2Lvdh9U+r
3JWTxsu/HpPXQsyAUs9NFdaCpxC7zhiCz4HDIVm9r8rpymjBNia2LJO4mgG/
QHZGyEDkkDwVUMEIElbLyv5LPUux7XgFYhIEYYISK8vusEqHCa6uOS6vOPe3
kk6DGc0EkbZieBfvMPKHmdBti+WS45qBRFfgBwtmKLC2lLGmb9yVB0NjMxKe
GCfpbe7KFek+O2xOfMIcFEcLkcodL3Ehtx2S4gQbEwHNEcjBQa5+fWLbXyff
mVcIsWcSukT6Rnj6YJzSjGUHzASl0i/fEm97ecEgenWrcrBnENhOZ8X0JvMv
akRr23p5XpDne2HDTji0uawhftW3AUcyRmEetTetJVFkKh1zTrWQ+HB9BnT8
9fJ/XMYLG8vz5tmXTjnUSDBR4iqag7jQRIZSeWqAo2u7xYhOXoqCsXXpzUQA
LUCQ/gvhpAp02dAzirXW5uAJOWten/HSmo1F+5ZdwOnTmhXSA8ruISakwASt
G/xBxcO7DcB/dq72NtUx9TGJLEDPi1AmMpi2/OsdlYLsRvEv+rL/J3VgCnV0
hEvbFa5FXV+x4UJW3XFVPmU5poS8AhdAd+FI7myU1cQs27aBci3irQJe0Uzl
UPTpZC4ny4eBUVbA8EXahQgPBLlw20Bt8nOgpKAdEvkyizDPF/e2yxhq2oLb
L4vvqJ/Fqtx3T8jqBnVRWCjWcxnZh6xtN8HV9u2SSp4R/6DKwWv6CWbbCN4G
PvCH8YCsIwocyjA0/xijyv6csvpctRYOruzvdQU13MqS/aNMMGh4DYrR784h
ubtlSQhoq8RsJP63AYmWz4N5SmICcpOEGXoxiqn5579C6u6ykBawcGJD6dyz
WIYClZEpLcJ2r6ZhZJNKaTN26GcW7yGRgAnCOdh1XBMRaOpp13QEVW2B1oVz
WKXiE9oT9PeAUXI7luQ1RqZGGRebnv9ZxR0wE7pVNEIcH/Wr5ap2sWqVjevo
18N4H4zOPbCXK1NvsLBtrIyS3EUGOxLY3x99kI6mJ8NpFn3s17Gp4eTcM5mS
i+MG4q2OxWI/cGPxrd7UTMyjJCP2lnGMskMz6XqCBkn4a2EAb0TVWhwfIeyN
g7maoH6dRdHeXs9pZ0NCH+uDavqcFMdJRTsdRIGY9S6u+ugM+hCUoJ+JEx6D
R+5Oouc56esM5CMpqGxAZRq4D3Jhu0dFizSO5kljNjiO5zHKkLMj01n2m/5p
P6WhmcIf4ORg1mnu1kSwf6nqC6tdx3YY74w3KvnPAHM0Jh2jjy+xGyFvrebX
T9DYkzyh7/scTgYTRFAhvorlkS3MYb1s57pTZLGO0n0OBrbPBDJkkonTX2vT
aVCKAIsSjVvAxPg+dCUU+eaS4/wJo8A8Ly36s8dRR4qax/lI4pVQH4jT22AQ
oJq8vJJrOKek3mpNQVT/iO/InKHr1nalNSzJnCTKGu1XShjhbKGOyA9mGdHf
2fzQAYVAadjsq9jrAUhoE+DSLM/L447WWYeakpFefGN3m9MV77ppWgsm0GPj
8j4F87YEiMehzTMgFEoHUUvKOMuFGrmoQvaWc0znW5rEjv9Sb2kx89ExbWlM
qzex3MiA2T/ZIVmlrSf0mZJfqvq1BUZMIRWF8CIZRGK2w875gJsYyomfcc+5
LIXuzkBOMcI5RIS3Blo/LtHFSfSfN5nl8Znba972uGoPCiPgucBcW2VQN6kf
1RrP0zMtq1pt7utXnhDEFTRydTI/cKa4YviJKuWpoOIxYZ4+XUCYjy19MS6R
AFJmcU1Ygj4rpGx3ruXIo0TGLgm859q2VAPInUqkgbfI3A4F3bdKKToBIJgL
2bHC65958x1LhEnTjphiJoKI6W4Wcx5JUnV7PMViShAGb5IeR/n0yAQSlIPM
M4HTGqzmisAtxc32w3Rm/vdwukYNYyoBNL1ZSv/pUUrQ/E+GfWZG+eIRWQE2
MBPpTyrEuNC9kX7AFgnVB6tLLDTyxJI7b8iwUpFBvXlXdfJv3aWuHsnm1sQC
f2IA5Imh0C2DQGP4G/N0Vfroc/nV0hYQELqutcrvH2DKzPgntiKGEG7CLZMt
NQe1DTvLm7mJLHadAvSZ83NLCM4QDSlElD69uBWcuMGvF9vL9lCE1J/t9aCq
KOXW1kQECZ/cS57/23q6M+ElPoQpeb4F/BdHE6p7RQI3VTyzBEvkWKvRF6r4
bbe8nJrOFGDtcnaA3aHt3HSyZBrAG238uCR5xvEbpXYU5HnraIi9cjnoGE9r
C+8HAXvV1qeVBQ3CWGFLnR1lRPziNWL1ViNLpIBo/bqM9MopsiuF1jkH0mlA
bbZI3Pwwsm4yzi94b4hAPCC6Rs3mE2PM5UYnqJhUBE11+JLE025Afoo3N2+s
98GFiTSSBwf459yIspLOqAqR3f8UoQodUpAHN7DEjswVU3HgO0LEaT7uUbV1
lYF/PWP+PRO35wYwWU+PcnM13nd5HKMA3LIf52L+MDO66W1ZpRGL57HDLUvY
1eEvlgEUfprnuo6c882Sx5IQgeR3p5dHgE4oylnDBXIPomVycPHRbYRXUJV2
49wWxl0jnzQoZ+hQbipwQT/zN/ExPRa94vQSAVXPGq6R+AeDk0F6zb7iH3l2
4/K52kfTY3CeLnFDz32rQsNhBU4pFLpzIWbjECAKyJYRVnn5HtVCgqnRagA1
GLE013XFnk6gePXzU4dvbw32FqBOS/mV6b56bDN00vJos0mPe8HSH5C9bgnQ
FcHBl3WjGWSx87NeGo6M0M+IfYRUL/64FB5t79WiZJxbl3oJuQN4vPq6kGPu
n+UuMLEB7IuAm0Kih4r8FYs56cIl0FC+ObqJ79wpnaw5aY+fD1ntvZS74ML9
GnPENJCdd4a64ot+ePJ0CtqTvU5unVTCv/ATd6NkhKFcKSPhNBxcjbQu61Br
+z9BeIOCTonBtiTl8dn893dznRAl8ZJlAzkQOZjbMSLrnOusQPED8E/Zgm3Q
w2gWXO30t1OotK7HiuBokCMo0NWpSN5yp6rB11v0wlZQPQkqHgCLHn1upl7R
6zUeT55kuPY73dT7Gr5ol6qwwOywx3v1D6LS5SeUuQRqak+Y2lN+gDahJ+SB
WK06FBuT9XvEGFifhm9RGwILbpMyBLI27wIBzZ9N+IcWqPUga+F7ZXbDTuwc
hlozJP/7XO3Wj/FRU8oRt55RDy3hoP9JNlV7sqnaPu4RNhbeHpxm6veI+txQ
OB7J3PPEJ3oGOQnj9/faKM3B0hHYY1xsl2RNqi5dU2GNbgBvwLjeUU5JjDLh
BeuSwEdLgJGYLxkTYylz6CA4BtwMQHMtAnJq8vn4hsGH8wjMgO8SyZC6/fYF
2u+kSyzEViSaM4hlpFqbxCeDqMTIuEX+gN3IPdQag1zuVrhLAqg0/hxqTskO
newHbDTwPhVyxa17gEyhlQT++8QO87eKfCn4mjqxsMmhdQSzwh1QOn2nwwXb
0Kp5roREXSy1e1M6isgAZRnXn0Q3ICR3TSmfm8oAkrnWBM5CV6tNQAx8ONvL
6n81lASHNjTpE9rSsEfe6vqQY/BJ2Jgg3jfZ+9FCklZVDz8nUtgUzSl+jtU8
3DM6GrNGDOM26nT0+N84l6C7t19GmyXj9ii8qeSIb1sMI+v/12extjYtTlDh
GkCaMruZKA3ATMrgO+hdByL37e2bKHBlq3GwVFbVp8V1hDu5C+H7JprNgCDV
2U8SmL/trhd2jwUY+zTBtEwJqisX5kBGjDVy4sXvBO+zT2UrB5jxBAul5uv2
rcdqJ6setMkbn2Msw34GkR9K2KBPrl1/7dtePM8AUf4PwPQmTqsEyHExI3Wr
Z7ilr4zOI7muA4PUxHQYzMyQh/vVdYfRp1Hk7+oAzu3oFn02aQmFgfbK0olH
7L5UiRn2aXa75iSzjG/hPdPxVrk516JHkZAeL1J74pA2/18NiB1HdZv3JroN
RVsjIUhnvIXA+7cist1/y22gLibJ5i9MIlKlFz2cZrl02XHQgG0ymB8hjagj
GM1r9hdi++GoSo+P641pf1vsZs0D6yuQ05B7ei3tfQvKLHcX15LZnkY+Zfl+
v4BiShW/42Zna+6vI0UeiaTjZnfN5UjHI2hRmFSbiVQd7/iQ+vpj49sw88QX
8tB7IQIEBUkOlbdcp/AQ/pTjjSx0z2T60029OPEhCidRKFQR6SsS+nlkaE1J
OV5sndCxZbo4YFQlyAGInw5I56SyleiCjH5cHvtkE874EcTFYj8dHT++Nrqe
3NIN4KKdCaQYoxqdUD3rQUeqx8u05xQ5RtJiG/q85JyUDc2QRkgQ2bTsswzh
w9CRKeI5BOwWrcT/x+fDPrGsXVx7hFhDA45Ch4wgjPHC9gzlyIEN57tABKGi
HQg8s2bLkFETR8Yq1dlHD9A7QntPlXo5vLSdx2RnaFkNiewX24RbTn1D1kSo
8hazlsufOdLsiboG0hcUjOKuLtzQjQfhkuAZWkRF5rqERIipemze0JPm+LMP
w2BBO2N5EudupW5AyYU3TYNvZn7MT2Dl0f1Z9ojjJoo8HOzFt/vZRp4XxoJL
4+jrGrpAH6CU9X6APu7jAIQnZWWwP7gx4KYVX/5jvTXgUoqy8IDOJi6it6WM
d0elD2P6uQGFX+ewaX+KOXBNBarO1QegkFTJ2XU3aYC1nP+Ybo+bcIEKVWq6
piSjgK5H/Btdl7T1nJOU+SjeB+J30CYUujlsEXa/jeIxLH0b4+8ilkvtxo59
/uwEOE+NRcNmzvMwIbXrauzPI3PhQIH3D22/XegWiEDdpk33QFRlKdVKvqcG
zvf89XV1PSxQnro+IxLDKEzPuk7Lobgiw1SWJkDy+1wY4MV/vTl4XIjS6lTq
dvw194yCnK3nSKGxoGCHYjtz+eLkM7flDZh1Yt+Bnv6yRL/lUnuNmMtZu0/e
yd9o3ozTKd7ylwRiCQrnjSPqkSL6RiN0fJNie4vyleGrytrM/4IWzQvRs+vW
ESCEEDEq92oOMSuUE5ka7TQ3+Xkn3E1+Ly7xn/HS2dS0KSANND1q0pyv4Ick
apUyV21yEnOsFOcvJGu0Ex4Z0S7SWXRZWGt8OZIk5vXE75HWW4P8x0XvsiBX
09F2ljuI5Q/F86+mY4CxgORNGgVyWNDpeNYevg3hJRmyMzi1/P3Edv4+0iGp
+R44s3w0YN2T9lfmUplVC2j5j+L3MT67vUvlFz2Cf1r9/IFNy0FBP//bVDaZ
kd7d7nITEsOkNyNNIMxpjGAmtMusQccmgEgP9xwRZrtIfHJNVETq0QB6Vwdi
quPRRt0kySCEj5TvViORO0UXb7IA5dcmsNvbgLD4h75tJjNg1fAEUUYbu/o3
CtHHYWfjmO8WbIW9t2WAw83clwjNRxyQS5xvg8OIwvxWe6Gz7zxsa8bpmyzv
AFTXpHsTgjIve1OCfzz5L/Rnb1Z2ewxTtMCO7G4zB48FF6p48H3gx2XL4n71
wqFd9Y3HJX7MsQKIEJaTUmVDECKKh2cknxJDIXEXG7zYIf1KZiA6AasgmfL0
3GfCwh+NIEw9O464x6K7e0cxjewED9NiiBMTn1gkVlPXBOb/Ka//9MkXmsFY
D4nD4LdSkDlr/Eva7O3ljtiIRcHxBnc3cgWXeKiSV8ZjQJuskTOFpsi2exsJ
+7lxT7TgbAfIldVBaQD/niHaiJJXpGdD/4P8TIebSGoMDA23ChXW7syvEo78
MoFDQfqiV0Bz4F6AVLua0k0tt2PSn1WH3Yq6tWikt5qd268e29yLRK3QcJEO
T9DSrkQ5GW382eBvGcBNdhvtZiZ+UtNKUpw0ChWXVdKogjLwTzgLr+UL+55n
1Os+2YABKDkU9eFPACe5N5uLe74alzMiy7m9/aYvHNAIpFT8r0MwUD3BkxTC
dZBe9+BJPTnVT4wb0szq6Yt1c5vg5FjhZ7oxHatrd7QcIIGHS8A0jGe5ecyZ
A5uh/TfnPEePiN+YReLKVzq+s9FzbzsoDEtLDpIew0OPzzbnxkvJWlKyXblm
55jLbzs2BIJYLXShYuXJf0u2ky0ln9Gh/UOoxJjrUMR6qghFF2i5XK3KznYC
UedPCKHLXRLonpdqUcZjF/ZnCaI1Q0p4T0HBVGIZawzXwtam1Ml3Twj+94FD
1RuVYwM+4jnbPCQB4E4jk03uLGEWrDXzDDMKC6lKBwP/dkMn9OaEMkl84qzu
hrfGh5SQzss8hVbu4v//fIlV5b0TxuKMJJ5zoJNLR7w5XKfjFMFCLY1w+Wxr
gBQTSHZDI3KQ+Oa7c5I7zHdl7PR6JngaRFva1+eELzvphzsOQjIfArh15XGs
L2JiOu7Lfo/ZWc0pnE7k5pgxgOl3kQpg6lc69FjamSX/xmVGEBisLQUtrC5D
smXFrnywwjdUDNyJxHPcanCmZ45/IH7pdlsMCJ8dNjanBFSzMHiclFX3Ov/z
ViLgHobfG9Kv+NuV44di1DiH8XdEbG29l+3jAFHYl0JdiV6MIluOo1TdX6yx
5rTBAJpggl3MbJQUw5KJ8sSkn69CVqvKN/mVD2yTU7/XqCofCuwRZjp9USO0
WtPEq3Ei+G2ImXUV6yMI0BuO3B8dvPVXIM6CQfGdFQiGZMXPCpNPki+fkyTr
JFpzBfDCFT6G1xi26TOaZJhN0gu2rUoNUaAeCkXNWA022GIlCiMIZpKwBB5k
rooRmD7yADGggoEWkDaG/9nSo4Ve4iKEQlkjEb4bSdvkouoD6TNs+MmOakmo
aXUp5tv2TUvm7tftIukP493lWCZ9sZrxI3EzrfsnyWThsaWKNfirU1Q9QGA7
3XguEkMwLbqQgC8ZSWuy1BpNHjBYjhWe0/EgyMXpK2VNiFDDC6hkx3dN+1kw
6/ECfWyIsSV2jlljwXm9BxYo8cTZwEMubyREyDOXG3V4kn4yhDn0aUESyhgv
9lLPywdD6MtPMPTAotqPdruAzkwPXhVj/3wUS52QEQzgDxrwgS3o4/xaLy91
x0QFrOrJCzjfNv3rqXiZb7u7lEZ8QMlCyFKK3JQAttOHvIAdg6KmdP29FmKk
sKZZblz5mBx9WDdFSnzlb0VyyggNuBWDVi5zCP8AUp/5ouJa0/SEXW6uv5Ml
rq0P8nO9jt8zyRn+kLW5mFCFq1V6ncrX1dfv6HQNGuQ7SE4wCmXSjumcWllH
qDKo3BZTFpYVv9Qa2S44y1C4FUbM3e+y6sbKISF95Llr/WtKowuVuOt/EISB
32c8Jk510ehHYyNqRyyIQeE/kCZwhPz08anUI4He3iM6PccdmlvWRzDG7tV0
u0iDW+8UHTwH0lBNm0eiBLgAVF/S2yW2l2GFe0r8uooqsMjJIBeBiS/2CfRC
00ed13xIWenxSUQNET/W1z6vy/n/5Pzjgeva1SqKvUHcHHRdwmyOSASluE+3
Zxt3fmiXFz3U7kzBsq6g3w6AEE4OOA57fARJHzo6KZIcE3e9uIe9w/tN8KDc
jLzA9YLL6Mhr6gfBlGWlD1yAz8vTMOpaxNEE4IkaEd6VdyVVj/26ClJnCrOn
5QD435mh7GOVmlIo9iNXtOPCJU2oRQcu6s5n4H41B+7Pj9M4QfqQAI1bSe5q
InWEJ+0EocFNaF3SXa/+QZta4EkYzexznnd9t2wTMl0Pr4gRHIL75fY9dj71
uGckZsUeLmB1hd2AZHF+v0eN0EmZECwjH1NgPOqWh8bFtzv5Lm1GZ+/MzZHQ
3mZ+Rku8RYk2tD3jtu0rBZXOgeL9xmNmZemmoOmZO5H2EctSt/iUUo8ZF8ab
HkDv23Oq1DePLdDppYCQTeQWWdHwBL4vVhadjKOHwSNppdYHBUt7ZZLCyRDJ
IG6h5/QGrqIPSaVUbGrcnrMl24hDvhTB/QsPrOHQBjG+aJyQD9ArKQqbceiD
NTYYk/9nD9b71L06klr6bvK8i2NYiIY7R1EIX9QLj6gJT97o/uH95H8xq95Q
V1FJFAkBGNmlBCP2Cu0rFOVBLPIk5lY11shnHF/Ml458VsTDG++wgJFegPo9
eDLMULyF8ProfHHGBskETiOYph/ToHfzSZy73D9nIfpIFfgFCGkT4kgntMnf
KeJSelvNWMgnikTxD+/fWQ9cD6tlCbFGusQjaAotGOAeH3I3i0yHqmcovVxz
cojUkMvf2ZgLRNSs0qidKgK3oKIPQRxCzL6XPP2I3vJsPog2jTOOccGebBv8
rXwd33xq1r7YkoSQWkRA8Hqyrxu23mEhTr+hX5EXQs/9aqffVmSq+LjYpY0Z
YRw2auF8aF6DZHxyk2BT5v5kKJCWQXznZRTYm8xApwFctlg9dQzC3zXfrm24
qwej+8q+AbbwxCFcHGUX8Ep8xiNtARXuK9Tq2PewhkO/X21CYGYi0xj3apHd
RIGgQhnz1BjidqIyhkFS8V4KAmzDEDJaVtIu6COulL/4oXu6mnKorGu3h7sd
sXD0NSI3HTrPX25RIxYt1E1M0tNjG7h9EW8cPzuD4J29WYxSlQHyTZjG4cwt
r1E8jZgHt6zI9TI8gJijgH40JgJufrVcMcr2l4RU1QraTGwj4oRg1odLzHhi
A/UUEHmbFscB6XruH5O4JXwPtH1rShCoJF42xubC7mu9LaMl0aFFRQbjNhHP
uFl9Nv//m3krpF2zuQP3F0LHu+ltSfkQJ0fVqLwBY0taaDN7cmC9ZcfrgrqO
GFtXx472xczRoGPYJ2rdb8+ovS1g6j+GjxUpFovoDSWITxQUmih4xEaewhNx
HH88GOoUSH+wGXkHgErIn1QhY0pGbiwH2umgXSFlkJlB1Tj8HBIyhkpnD5jZ
s0myQxeqpab55e5lmvRhXd6Fr7bnDIsH3J7RCZxLQMzaj4gQvExHwkYmLbM5
0xDHmN493kBXoLFed6FK98g+OD8D/fbviD1hQDr0q9dj0B1bj1W0zg3PFhv+
YKYE1Og7kXd+RknOg+fFwfZCiKndtnNbg9CG7BI+vsTRmazirtpTXhAQfBQN
8mQO6UJvSSW5QtgsTTG+fMP8pFBosJnwm9IDr5TBvqcF0vx6b8ie+dkIRlEq
cVW++FbXH7+AtFuwAWRRl5EpsmQKcHYkr0EMjaDQqPfIQJBTAiDO2t2nlJl1
RwZIJdVskJtfNuVHQgIU2eu4kHxw2FNS95quRbE/q0Ct8tJ1GPN++Tvz/mUi
3+JciZI2NSJZ2XCFbSN/ZdrGykaxRwlP0lgQOejYcGOGSs0nItbf+CaWEx+l
VhNXOVX5N/TBzo3ZeBqRBLjq0F+t7q9vGa2+BzFQUGjfvRvR8tmLtcp3sRgA
7dhsdOf6Ac0IUAlPRmrd+afD5BBZksRlMxNbfMlKkBm/+BfbuX7smjInagmm
BGYdCr5awgENL7PySqKB5lMjVeOFtCw7f09W8JOHqJukhqaH806+pg4V2nL2
3+TjwKWp8cFeFBSl9oMY5KTa4F90RY/eCpK5D9VtB4uD5/Qo449fzZJWkS2f
ype1bAUh4jtkI4/b/4vTb3pe/ewf3eqa22uFzOsQq5vg2CtAA1QF7naydOsA
RBS1cQ/q8zL+QqdFKuZU2g55axt4JwoviD0wTMP9zH6tFyRZ0B7F1loCjzsb
zHfgMPqP2DhOOE13Ln2YGJobJ6RYz/QFlylNh2ufDWHLpLpEEu5VggxceJZ2
EQvO1ztmxu//46U74Y9ZRhk+HQUw/AP9mr8YgBiTReNfyl7SK4FP6WB7yCgR
jyq+n31WaC6fcTX1PFdiXBtolwZzdbKrrhv1XlXo3PvsMYoqBQgB1T7msOcd
Ooc7t7fvgqIfqt0wy8Gdtpw1h+rakSXOhB4Kcz+0OC68jsPgqc/0HhLdPuYh
fvyKbvA6eYGkZMxbXdPbMN5eZ6ZVZ5hcLx7kl9Q/mYbWs382o2FfEqGGIS85
hnGqnd8SZ204micrROYTcTIav2vvhcMkqSfBh2fWeKiwlaj1yPwMCHWCAeDS
3mbgXJ6HOhuzr5nL567gMJhaM4j7y2qieBmTgBa6lB/N5Aj8LNr3Tyhp0GIm
l2IHnHvvUs/dfCcOF9uznVdFz+4BhUmKUYh2EN2IYkNTfhkk1lh7+56S/Oof
J9ZsYaq1ZOwArpZBFy4hB8OQAzns/kPRVbOZ3CtdV2OM22YISql6J8XTJlcy
coriYiU0mO1dC71rOnNIhzPw1itiU+ZAbTewKDTuXAb+1D0auLpIlH2LfUHp
hNxzhIxvWP2qD9kAfw2DrC6psGuW00JVyp/4GFUYAvCgtNKg2ujzZBk2ePlw
M6DsYvCUj9Y7PTrVMvS5W6Mo+Ed9LVvv46DCFwROxv92xBbJmD3NC1kctSMD
lo3z1SmqR4cUz1CgBAunRSHCxctEvpVpU/63V2PG7kHYdDstkupJq/xQ7UQx
hiE/4DuSOL7NUVADhwgURdkqq6CaRmZspS/ZNnaMh1pLvW5PThk71TqJNenx
ovh95UctXHK10x+LdjE20DqfbSFazk6Yaa8oZ5BE9EwS8OOLxk2yiOvE1wK2
ziRduGFQo8bRhsI4yxsHL5qh+76hgU53Y5XwD+0v5DA3T2F4l1RKM5l/50ws
aFK3PlsijQ0ANs8833l4AsvJDfyfZg0LMw7bSeuvgOrSgMiAdLuvmkWoMri+
DsSYhtDyWCsyS2bJeupo/qF1BW3Xl1wZJQeg19M0hhr+BR5S/C/mBTy6EXe1
1yzDtt3zNGufhGu8LVl5SPLtyTADYdVn3vfmdc9vUtg8P3FYokcDl36W6Yea
bVFGw9dMeYiciz3Hi6TKI5UIKqDcsh3EAMj6vmxIqsG+0fGAofGGKQw9QNSR
laWpH9ZKhEOHl1vgs4VDlGrsQ2P6Rws5DDWvWvw3PqK/Sqz4u6qq6WGlFpMi
ncFY5msDZjl/6tmNfrhvF4DwPQ89sT11qMFJ1IFZd7XBBUh4+yFn9UbHCnib
helIBftjF1V0CCucAcM5w6ldB3WoTaFW051UqCwVDWRLJKSm15MhWdrhyxJF
WPath/umt5V+sFb17hcCvWmXin/b3BcIruD2Ah8LUlciNRvzeW1U1NVfE6sh
PxxFIlB2eQDcaNu6xGENVeBn3DJxlX9hhtubVpoidDFcKQzKgCkSbrGysNUy
NBia3Zk+jttfkaI33pU1ILwyqPrhi7NxhIIEUzmRG31cQVL2JKaox6/jfoF4
VibjxPDJyTjVOBYIe1mE+HQZZWkWEQS4cW9u8O6rWn+0qfP5h2z/radYEF3y
JEbBMbMWy5EdDrchxdlvd1rQCDG5ES2tiu2KwoAkkoue0mJ/wgg49+SKknNd
iL8Q7SGGa4p2clEeBUGuaHoCMOFtzjF246k++6Zeu6i4FkMjv8UxeurFqbWB
9Ko/RvYWPb+utLE0d5vTStbMcbLxng8ZPTE/ly4nT7XXIDHOoeAJMPsUz6lj
HqG5O8uDEMdWnV9DuI5IFMNSjIMj37IBsM4/Rj2sDdruf8D3nDwzwpU2ZYdN
+ItlkDHHAxEblbmN+9cHc7olurfSJ8SrVtVL/CzaZ5a/T+Q6YDeKlY1Wxx0+
ajijo76s43hIOYkkpFFht0u6ddkaZauUBzwWFIy92FLurc9lXBLeYN2GBWsn
i//X7UsRHKW7fOExnpxrUw7LHBjsfZ/KDhm5w12VRldcpcR4NDDkjdOqPzP1
C5plRpYR9mAXuqD3xh7eGOiNZrLfuRDkg3nZpRaRKcLUwxnzsdXuoiyCRotd
X3DA0CdSqLBzE6fMuRYrxEAZJ218xDaDdRaGxmE9JlesK/PrMLhDT5Q2E4A3
pRiigWLbj8+5cA/Te3+tXUzszok33IdjyXl80Gjh332ExkhAtm4BJ2PrUxvK
v7K5d1be/6KAyvLQL4KQR5vYNUddkpsGJ/YCvDetVhboiVzo/Dp6UDk5zchh
Wc4Z6dsOMOsS1Z5hgwVvmwutsbob37aqXZ0S3FJxIWL6JXJkibgAXzkLyDoU
cJ7jtjHLkauv9rlGYceBi44jnRZhYrHluh0M5D3HArQtnYpYYsTXVQSQAx/W
6rOSXS1GU3FeYJ4CVvCN2oRq40tTnjANWBKYoyK2Q+s8XZNgregTEglY/PDg
MiKj9h5YwRUIL18rTs+oy3MLOyYjA52Btc5dYRx5D/TJNa5YFqfjEHfzNh7b
VkTmGeRYU5fzrhpA0j3qIILnRh7OrkARrZd48oiVa+FxFmedLUrecgkwlLh1
jdo9b0lbNqhsMGOXJt4IuGvZt5TcuN0F/qTq50dIHaZ9UiFQliG3EiYB1Yp6
vZrdz1UovEaT71xkA1FjDHrSXys/G4cbY2q/WuOvX3DNZ962P7v6mdotauJH
3hBV7HQE60CCXrIsm5evrgZdEXJEspuTmr45C4q75RyJHnidvGbNVNNCRjJE
0BZ4M20bmKaD3nJzh8/y5BQU8aRBUnmw14nsQ4ouJ5tZm5PGExW3gh3dl8sn
r7ZQVKzlcBKDWDsojlkCkWne2fkn4X5jBp7uKY/sr4ZCfE9zlMqocA3PwLf1
3DkNfrXyROq5B/gGfxtEVa/AQdGqdFdJgsd94z4O0C954DIXEVE4pXhv8aTr
Dy7CQPQbN7fT4bPTTKZ80jhRP8AtZwgEI83jnhxpX4d+EvLbfVvMVYk2rcMM
QwTdYH1P4wJz55jrV1/DWemt5oH+yGtpTJwgfEeXasiPywkgAbNt267/Nn3E
YCaQDBD2XOhlXqTSgRNY2RIicGXl//BVsUHn5ptVZmHrIsQ451vdyJAfj/3c
r+RV1UEL1i8gVF8FDD26EThdJGFlOXB34cwbHhKqvcj1poFSUNgLEMe/1/oR
e1XCUzz6f5ck/E7bAyImY1slpCAV6BP0xXwi5wtpZ/iWzEyMfdHVeahF5vcA
dbWzlZze0YFx1KxerS6rFNVaZPeauzCMZpz+kEDUghaUOu2hJxb4RRQRS63p
pPws4k7iok8i8ytlRiFjCvpIYHLBxzpqR0aZ4GAjyCIevlOGBRqzW8QQyS7u
roI90RO32aNqIgH8x/uqj8PxtdFseMdpRG3RBU/C44k79wZ53pZ+5PcxQb77
8eU/lftFYERwyvGG/SFMCFatgs60KrhkyClVAgdvtdusffABzwp+oCyJGuUm
RgInx78X/ns2ZMdAXatRDMfZnRkz72GFEjYiH/MW2GUQ+OiEriH56WhpqObP
xNJFbowrCJYo9QBHeZ29xlQ+zrzb4cuHL4Imjl/bfKK/RZ9TDCOZUiS+TJms
aiHuUtvGOQZpvOl5MAxf/aI0HpoT61kOx4buHgy/ZbYCYE6OTNNfByHmeJq9
ab95C48gz1k7bOSUJGwghTfl0hpJdAmIfHb7MYDf3rqz/EB+IBZ/BuAYYQBl
ZdQ2sI61vIbm0M0sul7RpZbscbJ7AqFjcDCaPfXSsVqq7YVLc9Tta+MF7/+/
7OekpBYXTz6te6tv9rjfoK1XD1xvSAYWZooDuPCHnOWmTYVKHHn8D0xDzh3n
IJuFB4gRmHbtC5FffUzbbMs3xlHLlt/CxDge8m9aiCSSH628l9LK5OlxRLbj
34bBNhfmWWJiv9umBk2z+7ueG4jAhyYNmirsX7oRNdCOXeSw7PABKUSl2M92
WvqMwjd710gRTLkMb9NQUN7xVFS2LykwGZ2Qkn6RS2DScPVDtjFXy7dU+7s1
U5uRy8AKyJ+/nARoY48vdAnYT71ZphZ+ksL3g+jm9eYWPNrwIQw8YuXAYru6
1lxRr/47sw8uZlrei7lVQODuamPTTpkyZqBD6rQfbIODHnGFXiEP0SnUuTUC
hOC2uWOobqLON99cLo8mSZaeFjfy2WvTOAXhc5NbTROGVGGbbj1yP93628Uw
mBk7QzPxVZ3Aqe+OzOj5fQHpsIbrDSVPjpdWa1Ijq2WeGNmlOwm1OL/PIbQD
q+J2cxYun9juXYYJYlAkJJ3ewcDQh075Tsanc16GsbVcL3KmTAOABpS6/mkX
jP+SjHW1OxPX/iSs3OWOjvW98AhOV+cs9s9MtWcEPb1XSXkR8cRJqhYHe+SE
uw26d4AjqYeLJGAE1ZDmcJCTZoqf2TAx5d3RdMjY0SncW8nfuvhjU1Yqmhcp
IvilhORDdbUwaeO1MgZTHM/pBPVf7a1/Dkf/DE0vOtZR5t84m552LEtVpmrS
Q1Lyb7Q49am60DBCzvrodBPDj9xJ7iCB4evzDGsaYvfWLQZ38BiDpKDsdRJ0
VRdV7DGXEKnyMeMWw75cJ733T7h3tz3/BCNjQkcY+JiXReNhYSp2kEkMgvLY
upwB3/d1SweXNjnXo6sGHTYXWl+pkhsE05yx8jGEihYiz4zL017xZjfduFRT
dGe8FkKjLXSykRz+stQ8sL3UGUE9DbUki2T0rnnECK8kiRVZY6ZVOURIU4/e
grqZJtNnBVxY1l1/ExVI5sTzGD0e0HDwvYNXswOy/LafhFkjuZt4IzW1lrY5
PZKQKOb81lfp8QijvrfPOmetBSPiY5pUgC2UFdR0UC4JaCZPLCp7qiI9mpab
ffGkfZosBzNFY4njApEWb6/eWRDZL0VWmwrcDTtxgxWPigs+tu+0cLe6Agnm
JD/SqtuFh6sfBH5OTvVRBGJTOjLiV2K/2iDuypwm8f8v9jQj+rW2aQ1fMB1v
d0715ZIV7NmWxKmvIDMaG5NmEEH88r3s2JQYXewrLxnGOSFZKKLHOTpMezgo
a0Oo+y9tmIQ9FP3ltQdZiy+S70BCEsZq0wOMfTNyXG8LSDNYg+IAyUiF4SDY
7NUkbJOM5eq0X9/4YOV3M9JDQwSC1ZOihuHT8Cv2EJ7yESYSuG/TIAL61OXR
Mm0BVbeKWH9Qkvy9lCz+VslEbUCLxb2AN9NjaQzSfxlhKjob5mOPsOyYDTTC
yIWCV0WB3OdBHD1X1NSdK5G9FgA4zNoSN0p/wF6950XEl/SME4adbRos4APB
HFOQ0c/BtRCvucviwgSM6a3iQLOfuh20np4rQOMtZwEhEgKkPanFspKoy0bX
XxoF/OI17PCGiUHdHK9UnS2rpyzk+8xGVfuRyN98s/hrSDWgXEVdEkN2aIu+
LddA8fHwxUS5jBkvxrmSLcxDoyLbXeqqF8FVKdvH30Y2IpLhoyB+SChvhANn
GxWpTCuMaupHppETTRtpx9xzXBVLsyYOrWAb6EpECHTCdJwbeq8ZaDcsPm6c
OBrX/ejuf46kzymJF3H9dUpfSEIEy2MLKZsIn0MwOnhoIoZubfzaReYw441I
wEHxVHF8LApM/80USH7e1Y0S1i8rvoAMhhYTG/fM7uMPcmFkv7ENM1exFnRZ
PADDye5tTQqxQy8syRCWScWzXw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+kz2GIoi4FeYBn9iUGoLkGo2uSwX73awuMIr6uszkItYAEwTZBY1TM75cjcA5WEszwh28z5Z3k3434dg8CczhNEfAPuZ+L8VpicFsFW8TOPvBZk0qWc8/8xb2QciHQMLKVi0xWGUSm0QERBhRqD62do9gOKMisdkPQXrtCf8b0hmEliVFPQBswIwiHprvijsrsqWiexpHI3UTBWaLmymcO95V8XNtX3045bV1qKWneh8lLBlDE1jcIgKJv35UbdDdyozFD/wNj4gCh/V6CAZABc9LA57Q7cf/bxQNrnDw9id4VHIK44r+b3sdVoF27I4pOGVtZUeLRHBdvc/qz6SXGqHVK5afuNf4Q9ut6Um9Rrrt3dh31//5qLXC4FkqQ4ug9/C+kUkOdQRs/V9vuWXRmhsRCgXb2T1FbDgG/4m0ju+HDOFWggLHtOo9EYDrYHcb+PhNNXkcnw7xYRsdPHO8pj1EUq9yX8NBDIJhzo57M18a+GYA42xiyUM322wLfCyOgw4RYBhTZJLATcToL+5nlro8YmGG7FZH/C79NhoCDvnyCwa51PkTE2q3gdhtwogTjnraViy8At2DLR7+PWSC7H/48Z9rG4vsrRl1sf59/RYuBXbg+fE1LjFMCiTZypFd5l8ig4bJnIPUvXDKc9hO39fWTkWTff/5xFRpZBDZ0hd3EtghoHbyYwC67bK+dgMx6MrTNDeuQg3Er9OAe7Lbgqdow79V2PIMG/SavygcIk5dK77zlfozgbllXJfKIAXJcacMtH1N3OMWCpZnp/kTGZ"
`endif