// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
0OQqPHDY0J8sNk7p6VXay6ee5GxekSuJSgta2LsA6VZuuxVbc9G6wHqyyE6y
wiN9wUYDCdKaB86+6CYcQTHDPovFbUfkZAqwVqKLdC/t9SXvk72/7QYYYxtp
WtODnXAG/WSQSxrcAEAmjDYSoFut3EJ0kgcZ8n80uOgqkrc+JVzMNXTDNoCR
Y4Y8jACP7r8Flg6+KQRtl08Fs4Pc70aMYPFnOf5ItBwEECP7SnH7BJldiy9R
IgV9naA4c31aErywLg00i52g17zazLKXsIt7QcuClyCth/2c34OHnp6o3pOp
bDwr1jEgIUaGmvnbm8NCYO7DrppAARG9Ojql5+CSyA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
m9Tga83h8DtOgRkZdtpDf/GY+AZXz2j8oo06ZMDeInbrWhENlRsF8vTI5eME
xOu2/f7HHEFX+kYvkg1K7UyL+Ul5R55IuidtjyzZA5zdkYI+ViHpi2X+iRi7
plS85U98gfhHR80aRwqC9e8bjr/hQcZvLYr0ONLxxsCSsT9bZTQW/Aieq8Wk
tcCkGrSTeAeih47Y32OTppzYpcLLuZMp/8nNuXK4WIQKQyD+R3hkhpjraAzP
5cnCSYS13yobbgq4mEifcz9a8gipl1yuftb/NligeGx4G7i5RnvkZTHELdXZ
74/LYwItRHyBbbBPxUotXA/2YvPg9TUOLm78y5lj7A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NW6QCl3fHs6MtcKLzkW0EcaNmRPCjjD+/h80vlYCqOpL/eMhE0N3hvygo/WZ
6cKAmoCuDGqOy7X7fp1sCyE5NRWi8Zq0SLyNMoL3ozM4n/g4NwFnva4YZwvp
vzlRtEyCo/hYJAvSsOdXYMAKeCVfx9ycfqetdgIO5Z+lEHMA88k2lpahYnVG
S9N1g8Nt2MbXDd5nM1B0VYboL3p+RHEguRRfyV9EZ4oGj68An1F1djooz31U
SMWXPorSmAVZNmuSgxh7igyo9qksM4ZUrjOEcYAID3BwAXhsdqMPNhgCPGUW
bY3Xwd48oJksijV/3FVhp5nvLSMpUGHcqnlTpfPxiw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gZ1SWh1Snl2nYprZjkqQUxAGxiFGnTdLGCFYiYd3xJXiwOaOkYsTnDU+Kg91
mw2gu94SYj7Hj1nyAXPW6RQgPBlMbKHQtjlnC9LT/bnEqmNMO8WRmLSPXSB4
T6GwUf+MK7nET4Gmna3uXUl69U3ZHkQbanWHPxk8Qz49u1+vtqU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LXzuoxd8rmZXFe7V14w4symtKz+sffovAln2zp3ZFHU0VGlb+VfrLW51x5uj
0YIYBu5MKjz5PwQD9gMdkFnaiFFUia2Q/T7wcWlpL2v9MSQD2MpWOn8O0u6f
Caz/m9eMkOicl/nAv0cukeBQ1ATqW0pi2XQhlHI3e92JH09kz3UDoE87fPsY
KpBoOCNr9s8zBUNe1BRy121eFAfJSdGr1Qmb9K8E8lr6/dOwFjlh8nO4Fo3y
XTt1gNt5XgFdMemojtHls8SAHGjhfxZvUxa1PUI7UYrj1dGcib1AwBcONp3d
iLVmAjFHvruDwrHop/xk2pgCCC2llbKpYmlpzmYbE5TtTysd24U/sT3brizl
CQ+iu1t3f/pqfq7s57IK/I66jb0209BqTbByCQV7X1Se6Z3V8ygUhJ52eDsW
KVZnRBGelaUyMvV+FKxDn0BVtTkz15WxeEbgbfwbJnLcfqtfyOG5JQs72b3E
XjScfKAWQ8ALWNttSlDHTLyM8dObnJVY


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YFYaR+/Bm3/K+dQ2sezmTWmXMeFlBYl5/GMQzFiRDtdjdJ87VvHuwV0E5N/Q
RZ3oEPAyVJj34fwe5vqG94vROcpTh9EDYiuJMRg+PKVIRWSo9T/9K4vSM2D+
FTWXG2ZcgtW9Hh1/95EmS6uMzEtyTN4XSeRXezAhprVEIp072DE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oh68EVutJulGzwTAQ3E8zF+Os+vXLZt/IqdpbM+I/FA7hfei9xCLygqQ+Q3E
yJbHkDOYtllkacjrzDcLZ02EAjKCdi/iobVAZvX86Of4Rp9RaheIuPgimLup
HMPrPEygqTWGirzSP7M35J4rYgmL4BrrN/fGsYnJ+msVnZT9znE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 22720)
`pragma protect data_block
mSHMxmy4Y1Q2h8NUDEKrUBjnT/9YWCCxeLkZkZMMSVSh5pgj8xHiXwH1Ms8/
Go1LLLosOjRGaWn1KAH2hd4JqSJcIpStVEtC36TZ50rGFLin0Uh1SH60lbhv
Ma4ivLBPcep4KM1euvFTW+q56cinWYiqr3edpaaHjKOtUj1OKdkbhNRpSp/D
feWRYC/XuA2TTrKqKX0eusCc7hJhxFNz+pPKsO+86/epZi6HxljO2y/yBmt8
ZR6wq1YCeBYa6t0DJISgpS3r6VpGwlOynGZk90ubCGC1mzp5rqlSRJKhdx05
6wVtkdLq0/x8U52Cb4H1nutGByuBI+HFGWQ9gZ0BriVU8UCYTUh1l+SeBPLG
WFaumsSgZLn/mudPJDLj4BeoB9HPDDUNp4eEgj+hD9vgEoU/oAzXS3aHsUZr
4avNpDiVXv5ythuLVUq6nbgyOoa6xx0nJXAQcKovOfzTDym9NIbdTFMh7X7n
0SQi8WHDrIQTAOxxw+FoYxHDSRWhST2v61Nn7rFM1t1hBzjYXk2+q3LMeZnm
po45cbe4UOCYw4jOyJRk1pXMiS15J8xrtjJ6BLQUGbeHJApxkaNlhzjLpUbL
VBmfoDt/ZFkdyDEoLlVxLGw+pmy42qgFezBOo9QASP5dd9kCZ9jgpGaIcSX7
X0+Cwb5sbeXIV1sbCLILYFe86/RSUyraMpKsTMk2KAx00ozqDqyhKiFQeCx2
Bz22azinJEiQnwFX6B50ELaZq/fAmnoOp1c3tusH0SaDp/jnJA4pxlG0NUH9
63jDnbCYiAlZasFyG2NmobJTFaCwD1niJ3AAQt9YdZTvS6e7xzEww26tA/ZF
IvFkOrAXPjwiSJ/IECEtjdtyXsTLVekhRct+a3Mn7Lq91s5m4rPbk0o93JZT
lREa7CoYKcxG4tQKCuRHpPgsMKCLqFxvBpPu5lVQT1pVlIwKbqX2uCrrOo8w
Bb8EavuSiOENphhYsUAJq8Id/kU853+Bl9F5ltu7W6i42+o8npnnJ349Bruo
+w8wQBtrW9RhWuEmGNXTaqCigzwRJjUmKp1DJWuYqjlIihfmKk2YiXsTImT8
YYQYyUzvAypjpp0xtdJ/ORDI43tV8nfH74zirbG4+p0xZJWGCe0R3xW/czjs
3PNbKOc8Y9yBWljtp/K1M/S3J1RAWLSlyKHuT3hU+K4ieEQ+3IX9nAmpE5Ch
5CYSo+60n/VutMNnUtWahCtTA8AoRGldvJKqyMtIgCxXFdxgAsT30P3IkC5P
WR65hV0Z7asvlyv8LQwvSky0rG6IlXvJx/zej5Hh/Cih8u6VNEizqPbic9xO
lGzJq+Nv5m9+MTT+OqxSRRa4XhyIW1lXMu5NB7jduPtVdTnXs2LRiNl6uRXj
oWgEvZAefKHGp5Sy5KlvvDPuu4e1s86pfQHPYGoWMcLVdaNuXa14oQsUIvO4
Qs7X9Yb4+KBd/HSAMAq+22H4N2ng5gz+SUQs08dDtMnu+lqJQdHmY4t8UCgg
t1p57Y8Yh5NqPePGcyXUMzlFk547DzSIKIJDI+MsYqKwBwG547mewIbKICbM
ur5MpO2SKTk5FtRo5VYP+b17QMhG3u5GC20Uh/2C/0XrXfhji83H2yHe1uA6
BLhTJZiSw3k5Rli4DIf5hCb19MbfRG6t2OOnhhBBd3F0NT27LhcVjAiNOTq9
dML96MtLGnMqDkiYQCVKPKK2aRT5/GDlf4CdaBjB5V59RB1sZpyq+LxdAmPP
+2XQkP6HBlPcnDc6prm5FUk5g+o5WHATD4H7Z9hdlk0AtCG8R2GeFgTo6i85
PkniidSLOZFexQ/ucr5GwerhjPAz8b9H+bAMbG7puBdrQJznh7XKJuuWsRfi
+vRlSErhtmaLXrViBVq4X/9myf2u5RQ5PulqIBopqGt86AxR/GwpMZuSGNTQ
5IEZ8Pg1wBDXuwx3sIl/bN5hz/bjTiIbjR4O5ua3u+FfMbLpXR/BU70AmQOo
CjAZeqK+G/iM265AKb7XeZFt30meICi9cxbBDa90YrQtPeI3WIHjDsTx6AGs
SuU/+J9cAe7lCH7TwVPko7uRjSBMh+IsDobaRALr0aJzKDAAqLuXH96rd/kG
riUh9vPL/wHsv5T3IOYC8RZKM/Sn8FvpNXLCXKAbLDnSupsqknp5G4/S3fWi
qJSxFkav6jVJaH8Kq3XZn0etazG4xB36pImrdN1tMUOnWIlYc2OsVVyCuH2R
V6xL9O2S08nsAORxZuaBnVcabooslsXSBLdhRmc7PnJDBmyFpeFz/BXZ+CtT
uG6N824PSHfyAFEHz0BMRe0V6aRvIxrvnR0GJMl9yvEJFYQiA2CmBwUmgSlb
KqZscqmOSEDk9UwGogK9O4X6+Eyvux+UfjhFzIHsvuMZ2pvHOQJ8aFBxdhJM
Q7QonuhplOtj4J50qdmYkpN9LFb14QqcJCWrfIHNK8cPVsu7dv7NXDkVNJfE
lc39BG1rz8F8RDr+YhfKiuwVmDxR76uTD+SmE4GCiMS8c+AaLXRMPpDtR/+h
VH2VREoF2zk8LUHyShM/qQR9ruFPZDKLRs5t8geLAB0NR26XeNMnPJz/ZAmd
TcJZnIUFAGV0xjCrGgnIFFbvZ6TYFnoCPHVM3FXarmXuk/JgrmGB67DmJuIC
BEDd0/rGD9n6PmlD5WsuanlNEmBT/y64D7VisEGLcYs2qSzN65TafST6RXuu
CJ6KZFADV7vpJhSQh3TL3QEO26UtOTi+Ok4VwtZJOO1bJnMLsJxy7CDHsLhW
GmbkGsYjgiW3h6s19P0PGpBWphTTTlF+JRWLE+lyk9+YDH+349uF57SyB2bi
Ufx2yqOmRyeDXYqCZnncKnuidFbPn4FOQ1V3oIoqGLWKHBPNBwXMC85CZ9ZA
l1cjcR9G7W91yOBCGL3w7GFfev+ipr4+Cx6kDJlfjM+C7G9to4NzNTJaBkuW
PbzZ7IqnFTyzY3PTq2jYkJ9pMkqxDLegi+zng0OzyvRhNcN42rSPYOi33NUE
egpl5y4X8Y2VfYTmtvJvIY8NuouaYjn3hFO0ggWz7RWW8VgcadagsX9JsyWP
Ij63+pMuV/abv0N4j6VwoFQ3iiikZl56NFkevFL2XVMcHTMPALf1/ZpPnhQ/
bweUMzlicBCjiAxUtdgPpzS75zsZyptQ/dOVJTTHuXLeo9gq0uIuwHvgzp5R
1c0pA+r3qXkHBGiiVBoQdzMtG38LBIHEeKPFnvJuGK10S4QhsxH/3/o01zhg
JDPNUONtQPkSYK/wm1EyBVyftlC0yX/6pKJQfsdg8wnVluYBf2nuPu4z655D
oKSPb5nxZv4pp72FRD3VR4Zv254vrVb6sIjQjBtIFGqkHBcm33vHKIwzz2BZ
d91VduAWOdYSx+gumBN1WPXX7Ob+UGHD6rHAY/4oiupxwa39nPQK8Kn73i9N
yPooiyeVFasoIMKfhUaXMZWYwKjJacx72HjtKGGdTOG2t8PRcabPr5KtBVJG
ZqnZuTsR0pyhiQ5CgGGaexQY5IFKv2FA3+qXRT45f9MWR+K/vipPUeOmxP8m
oFfpn2QKTL/fdEOdVAAPf/imSDSYi5n6KfBdj/wm0uJzgZWoN2zgmIN9pWtU
YFFbDx6sSi5lVgfMsT1XGHnjlaIOljKwegDyWqO1d7mWg5FGyXY0YLdvMkig
FADNqR+M2vAUozZyOM9lW+Gt7brKMY/mTKco1YMkWIIf914i8mGLnaxweJ0Z
mLCoHhMOpBbszn23BUvZyqgajzoSaqEVaBzWk9uI2kb+GRpjaUhxCvuHmhmq
XhD0U9y/vlB/fUai+u1vx6HrZcMV3SHzisI33vxuXC8cs9auaafxmZottaJp
0aE2UlbmVcW1zdn7F8zi1LV+vuw1Zfa9hU0wkiosP5j6EVeAU+UvwA5TWtqp
TnywQYXfJYDVNg/n2thRlj+qPaePC4s4A+/9N0jjfnObytqcBotLfJOQ2Ye0
4RqO5k+mkUx3j2oAL47VlxXAaU2/uyzUn0izOoiDiOS2GVvuspDhwWylnh4L
O8/VxfH2z1mCdx6TJ1gJc5FsldSP6DJrDWDrqy4YHghVyAMtDpVga7OwqEAv
NIqkGSPNJrctEWLCivCvTwwAIa866v1dyMvMRVqFEF4XY8sgIYvxs6uhdD1+
OjyxTBtEbKndhUYz0xJ9Vc/AyUBr/bfgvid/xUhP06L6Z5/vf13tnRtrHawo
f402yCEFVZpzJ5oYDqQPNIVXO027J8z0bDOjLHqn/lbDjHVjG/YOZ2E1cCrS
8WzIIqXrxEqY//n0JbRPYzO7rINGr8M33venanbf8sC4Y0sCPkoFQS64STk7
icAASiLo6fXLZckOxPSH5wstqjWH25jhBmy1RzJBZYRkAnB7Mp0A92Gg7ilv
euU+NhCxDyg/ENMrCe9LZndvJVDvlxlhxKeKC6X/BDeRdueDdjs8VqQxehGL
D76Wf9Q5bim8Jmks+pnUdmihE0vEO5K2suBjxrr+PduPaP+aAWjXxI1Ii/qT
RCbudFcLYgSHX5vIwBEpHQ8a/rYpqOPS440D+laXm7cGOl45YsLAem3rObAm
WDJGa5QcDCj4Y3K65x0KqvBPeOnJRpdflwB8AXJIemxHJwf58isq101UJDvb
1NOOCw/MbZzAHKTo/wEL6JC732qDIiwOcHKP9Uveqt3O4gfuDEZ9duKmRyBF
7MWUMFTfG5AG1Q97OMKvU91Nxv+nVQ9uLLqa3/dZZ7Q82bDku1Lddf4OQ+oj
CI7Sp+cs46gcKKQVnr4zFMezB3crV/s7TuQG/ymh1bFqxK0CkurF2yk/B1oA
bNijBOBlTnmeS6fGPBpbhHjpN4Nek3EjijnPIjNM4v65S7vL1LyKI2ToSCvV
WKvYC6d3AdL8gsL/n67eDVFa5Zsz7Kb8rDK/sLMIdsojDE1K4+J56JaXhZPC
uVN8/5uJ4YV2ZAYLL/xRhIqU9ZGWvfuvvDzXzfFhjv7DybaMdYHYRTlz4qrU
ClSw3YI76VynnF01IZYpmENXBky1W/O47tEQpbFkZuiyJS5sBB9VZvThWEQa
XkHVBb5qlU6Y49rtikhI4ponBxtfSOrWcpLJ17Zl9gGaelK3YK+elB6P0JB/
fxJFqzqTBcXR0tl9rQjfNE6xerRuwkcvwUeMBuLTaJmxG5w+OO7J6T7jkS/E
IikOteuQY/J9B8VV3gEAObWfdADbYjEaedI+BOkEk9gHXpXTawqNrpVIPIKJ
hUydJ8388Nn6vWZhSIOOijvJXloS9TbPDNez9jlSA+ltUTPoDda/bxr0sm0c
v6LH/Or4hZKIN3hIl4AtVOlvE8/sdZPUiYxYF4OSvNt2uIqqFWRUqBuI6KuF
h8Rc+uLqAGO/ldfLbo0VZHISNoioAD0NK9v2+8165tU/26ghU9jFrZQzuxLn
gSrnaGtoBNx8yA0mhQ8ieNSA8I0mEFsOkQ+LvlcHtuj9tTw4q5s1pOYeljTF
iNTR9iMDW4QKJ5vBvVUOFucDizsiaMZnCeplGUGUGeR0WQ21wPtO0HrtP8as
XUn6F0rhNH0HxIGKK2pkJqs3EEXZMGMw92lvoaM4dM5AplsRaWwk0Zx7UNDK
DRS7SDpEsBB597zoh83cJP2wSW27670srCpH1UWJmS+I9YBEqxCMpIJl+PwC
8VTr0XxN/5ObEurz5IFbp5wpDugbFBoALkinHvhswYfSdyVYjIfCslOGLo11
SloiGeGimj4GpeRYvbS6rPl70V3WiPGsXm9RcWrus+vJ7Fys91/UZiEF+3gR
yokYsWPEeGE+j4ZYJhSjibVzo9KQ9Tz6lv8utCF6oRXfGgnEsrOKZ+MiACIp
YXj12YfUoyRwX6X49J/Asenr7WJM2+6Pe+Fi8reskDYYqaCoUqMzT4nGh+EX
cQfFGxH17wcyX+AZ6DHhK7R7bfoip24laRKCrgDe//xcb8lupsaqHbw6LZOP
N/pTn4kP0CiqhzqrT7IaCncCt1dsvJZ4qxzgJ0B7ZItAalYhkFBOdA1WrubI
qy73QTo0AL/mEjqCuUZaVusv3SGkhLSoyXwauNKC9mziDCpC5tJ3im8jgSK0
vd99Q9MKyHzqOJRWf0PTxlV6y+OgQDADt2Y9EVlhRJ7TYkDMroQNOn9tvFrF
FeM8gSKUWY5P7snsuB0sA0WcI/t+IHGuLdLbZ/hdTKA5aIS3DOMgXjYUhYdq
hn1lz3xblfvGWz5fRvCP3U75BFVgDk8bckpCzmGDxrAu2dbZ8py8OxL9Dhl+
s+bfCJyHQu7zKPiWGxtruXiX74rZuYo+uvRFJ4shuI/60OML+JQPzSgPCxv6
oOscHyLdrwJuwop4QAEUbVLDeo4HFkR3KBUwJen2bZBe5ueS0AVTUKVEO2HH
r+vWsxjBIrjf7p03XMo3eGygFo+QM+DVgLHlUB1e1QXHDJsx6WVIkB376HH6
jMTFRTzFRFWaR4aKsrc0tJ9pcGRBIB5DToMh05s+LVb5MySB0b4LUvHGOx8a
20R6saWYj1q6FV11z16icHWLszHDkqmqBONppBy7tzjHL3qJpqT6GXBZOdNp
hJTU1K5R0MKuxh+ORFALJjJaNaGSh892cFyVbpje7We0VicyddlQo+VFAv4N
ntioyB/RwgVaUrd2cFYgsTYRHuY/EjNiEOPciKZ+VoU0fPnOnmLzKIBUYNOc
bcudaQFqjfPzmI6ijyAMHcccyuxB+w0ZwcXeBm6i05ea1a82QKY0hABriJrF
9/G7lYNPcmKFOTVyXnCrOpoXV1knEOO5oNJpCU/WsJUC8t6K7cEhNUBKzwuL
vYDDKD3Wa98lGAND9qkXrt6SH1c8fv0hcJI5BkKai33MJjP4Ykj1qVTrWrXG
IJdNy8w0eCMo2EBJ1CHHTJW1/MQjh3Se3dHz8+PUCme1gcK1KFMJ1Kskiej5
Bdw0YjxxFdC6e14RAd2t/CavDyuCu1TLQKpzaa+ozpT+kDrogw4SeTWXYJ2Q
+rnU4mk1YzcWUhpWT08Qje5+mp5Snnc3koUJM/FH3gqH9IZnk/TU6Df2UDIR
MapobqZOZECj/9tm6w2CoV2aNZbsig8aMZCah0fieIaUVvSeR0aSFZfaJA75
1lAfTRyIkSTb+HfwW46ll3aafLS0HOR4z1O7L4i+ZRrCUyGO3HvLSM0da/+R
SNqe3ZDLvy2/eO0dutd4TrY0YbfAlqDVu0/tU8PSK0TFJOSUDoQoaDuDrtqk
nkQ2IAQ4wHukVPgH6a95C6dFAFX8lvtfHhnYnWHaRn9b1F4azZ7QJgVVhFLt
jzN04K2FlsYfRUAvOsa0B3KYgwFjXUPtZIAr6VHVrZcu7J/4VwkKcPmZI9jF
IDwJUXJM3BF/9FGWTFEA5LQpc+QmVzWzhTg/oczszaEEE4t9ml2gGOuYJXko
DUUOjXA95Ao0SZo+nZ20RShxcNAfcQ+Z07FsfyXEbTL5EYsyzW/8HTu6Xatt
cVgzT0YNgmn2elpY7c1CluAEnMmGgapC7djwicss9ktkfOTDiE5A2A27O35u
IRpLRO05RGCTdUb4HYKClkVPmABIzayLJ4LAGwUiw61HAiqyRLRkhCuFE5gl
jeBeQ5C3sfJ/MgMG/wQ3FoSgvhkO+oOVvPAZJHwwac+xFKuGPhY/C1AmPdvJ
H0vpCOX+zWMlwGFt/wc9Ej7px/VV4f6BEtBaM2UnCc+BbgMAzpQaoaelM6XA
uVN8O/6lPucp1z+T1Sr28NCDD65jz/6A4T28e68YumMPYIBErZ4vUKR0Coj+
wGs/qy9bOSWhnblTNJX7g8rCmZhnWrn6bY9WabQHReEO17DLi2DszAJeWOii
j6YRj+pj/9aiav6+dNrjuGw4Y8nc/hgoF3O5zxsIjiSANZs7QdVYEdEuVhsC
l9Z/D7Ohu1j3fiOrxzald7qr+jf3xMctth+xvG8lBA4msMpgGax1aT5tZN8K
LGkSNntMGZstDB9OTraHR6FugS/viPmS7GtTs9AH8ygRZM67mdMBmX+bgu1j
X6AQJViu0SQthyViU9rDrsWFwvIdIJr4Na4aqSmycFijXD7UU7bsua7GDD1/
QentjUWMfMrEP+8LBXr22+KXAmF//bu8QItNNb8JtBH8z5oGCuzpzfed9S5R
Zh06iSQ70rrnKxkgVNkXB204KEQDcJZtUAhyuBiyO5HYAkvsuREKSOSCyc/Z
4mT8y5hP0+U5mKB6PTwgVskWLrCpj+VVZvU/DVREwMboZk1qIZpfyucSeTYD
q+iMX6cHywWEOwaiqVGYKH0v2V3WZRyFhDvaIi29yhMVH25ID1xm9t815b/+
7FrmRKsPnNKrBXGditc0XwbjgIKSOcCYJ4YI18VPxH1+TmL2d7ECbpX0AhkJ
AIbfM9qWEu2Y9Yjl+yqpA2j+R7wopXXG9T3GswcJGgoc4Re9mlDDRguAnPq0
xuorR5hScQj+dkY+Ew8E4FGHkPMoT4/G03SG/9zgc9hQNeP2yjaZWrYo0xg9
hahmsiPU4jeizX0kqj8GIllhP0K1hlnIbQjB6nMTfnFC02QG9U2OSjiun8tF
t3CG1irSXTgNQQJc6WiNjDhOG9cQAGd1Z5HwseDGte0wW3sMwsrD3lRpVTS2
DLKpuawtEv7gocwMQ+DMkm77Sd0H3JbfNun5RiA7PKpFFxhiNWa5DDWUsQu+
V0xBT8scXQO4EaIgzs9miliJth+3axedXws2+becKtbuxH51cPrHNYJH42Nf
34xL9O1PN+c0QWA7mYe5yjYooP25DT8uA5YgPssrFWHAiHMIyt6A9zDvhXPI
l3HsfkII63ZBGFZNksCPqyRI/LKUsaVXVM87T2Ht/GasUNYEbJK1Lo7xQWXT
dY68NPdX4/cAJqp904MZbJcahpkzm7sj0dq1ezChjVoJOpiX0RB7emTTUnc4
TGHIGwlRmwBeahFJTmFkaXU3ZL2Oc3i87gfDA4SeF/ScdOzZ8PABLDWKsEXD
gOCQQ8ZdzJiTpeTE6xqCB6xnazFR1R4khXdwpsymm2Xl2HalYe7O9mlRdELx
xm/q/v7HSMsxsqVEJ5mclvgDNfzV2lu0BrpjkmU5Hopncs43q0Qgd+SCmzey
FV5FnbRu+NuDLbRWKKp9FpTG5D/GGDO6wa+010v9bnYdDC/8J6/1GDbSqks+
TTQnd0Rj8aJ+PzA7kPds9QKMzDm+9S7VL3DHNTaR7HwPRODjIGgOrVAFXk1u
5gMarzo/Fs1MZik1qgC3vUBUXDdCqsQjcXX9xqxUDs9zt9OqMWVv8pDERY47
FF2Q8H3lZ4uDe+itzgYxUyNW0pove5RsI+LL+K1x4YcSaQedHu5FinL5yrmZ
tT7WYWsYaUuHMC1j8MisPA/1G1bvUGir7fysl4lUHiuG/SiwBOn8YJHWQMMi
5qkC6e4hN1rCnkSqVBhDk4b/SlGpN5dnckEJXxbwWS4fxzrMUgvQ3OKVgPgT
srdSRiUKk+lIWqQXrhmO123CEImBnOX0xZtoz4IcJutX5UwRADtmw25p5m51
pFBjf+HYSOI4bJtMXlOhxGMAleHXZ7ZZMImo2p7g7ZX3C19RbhsCHiPq4Ij6
78E/i94rBFcoFFrj1oA3HZfrOpiG3gOAW3jYYeiwjL3+Eqyo+jgrs1mFn55D
JnQqQp7YbNgJLNAAMsaOaPc0/VZeP6u8EOLC/Ez5qA1WnNKBDI2UnRCky0N/
g+IRR/s9dFgD4fiDem91+ftvfTu9DySThpAnjlVrIkNEIg8wcBGA9GsUrCLu
BRYJughimiz49wr/UROjLc8AQKslTo2ZGvHfawLdai2o9ou+e5Sim1ruQHns
TQNTiZnQmkseUBf4iswVz8L4mrQ6SnQOb7GvpvTEA82KQcs+yLLkyJshk9n6
ZVpFbnBforhz7iPTZPgLjQwhqUzjGWA/H59o+hpmDS+mV9CmUNyObMTajguB
cE1mOs+NSJq+Ll+LbbQHFWzzVy5F5aaTJ1nt796NEKjwghwGhCVaNBrmKWOM
NL6ttNzbLHUZekQKTgFKXe5yZbs4MdcYWfG0SJuY5+CaE60jcyhJecOw6jlI
HA/UDSP0iIER1KVnjtMlaHs0jsOZ6QaAGIXrQKwOVB8p/DbQUEbCZiDAfAfs
9OrVDAci1L+88dQxlDjCZRDqmoryoKak+wbEJQrUhuUFU9ivgnxxmHhH7TSQ
566JUP3j0W1yd+7ZtoEJi1GUiXQpUkTuCAQuJxxjUhJLHYlPwj/1xlmt/J4K
7nEnjOfmZFGm+1nJD1RA9R3iHeQA4WYze7KVKr/OZlWzLG8r5inuLVy8AfSe
/QIYcPO0eLfLndkjjCoz9dp+OhWvGHzfspxqTJ/mCyF9HfuWv3V3WksMlQoq
EGbsM9mLLbHvyqTvtHoRWFd4h61eSU/PKRNQKmkxN7XcJbUAhwS6j4rHc2Ew
oOQLB81IH55ClOXXfIlpoYVuVRFP57CtD3PexbtkZcYQdi07nUyfwZvc+B+A
UpXbOdY/R0LLHiz5IJRsjkBsHoQXBtff2Ro8obzKHKQcQZyqJzCnRITMFbZk
Fnls9sXFEw5Ysirw4xrFIYK2wrn7yeAKKpQ5r8KXRc4Tps3a1ViKua48NHHv
xJoJUcxf4lnvtgv8STpMZReRY0quuQGpSnEJaAy8KiIudEJyy9N4VwyDJIyP
/F369tKPVjWtssOyo0RnJ7dZ6qzUio/9aWSyTsDMxgbbk6j79Cj5Qv4QxXon
eiAzUNO+Glku6Ho/1mY/oP/lWWyZxCr3KwFQcuWUO2dptAPNw+z7RCyvsclQ
Zfc2wZlUkCY1ZY2+3cyaUTY8SznYMT6CRzWVo2LvCVyDjj6mJFoMPhMYyAKy
wI6B+Jz60D0PaPxcOxFYdSYrIR/Q8YsRkpceHy2qLf9lTD+GYvCfbpsftcoF
8hlYs9AFYhMahKYMP+E+rvly4rPtSTyeoyBK+fuJJyAaY/wm9leWAVG9uDvF
p+wrW0JTIdGklPMqnwNLn8lxMff72PKa8M86jiriRFm4AuC7gdE+FSux+tbr
Dt2SJGciVtlssgbJRR/D27lN5CLP4RUttv/WcbZKhuen+iant8meDHL08KbP
ycbhyXVZwnKDy8g+ZCu+LkVhdwXUCSHN8IqF0RWgPnBA+uWBVyflx+EYOSII
7dgpqPK9ZwL4ybQSs3FZZDOrpbnfOHpVw8uuE8TXJow0WX+IkGY8Jb20Mszp
e4QlDqJ2B0EjkrOmXPDZQ42KJ2rGANK2ECe65K5e9fxHSct9R7nJ3neGdSWx
XvV6JMhvvzppxCqqd40pCXS0G1RnVyBK49k6/2YDxztkJAeml4I+ieL+2nWL
3Chat9FaILwwp09Nrb3ZLXR3BUC/ldnR2SBwpPUGp7CPIaW9Pn5ka5CLvYDg
Hf6jhtKbSEb3NX++71dp9k2zIuDcrNYEtGib0lSh/nYSEdarFvG9gGdT/gY2
2wjRA0pTbiEUZszsQpoSQdiecJV29gDNP1vjQLFY6PBq6D+GNQp1wWwnb5T9
yAJaI2R9t+3KDubblyplGjfzmcxTTkVTvHFHQvjEHLrsfqfu1Xg1aVIfJ6yT
ExQDYurYtmAsTNEvWTKnn3ZA1hGxUYTAo7nbMVaaaD6bJl2LQtOjgiZJhDDT
GnkaPoKkqQZiEFQMk3tYYJ1nylfTJMvejfA3DrX0aqxfbqBrX3qPv0v1Uz+A
q4dTAfN3BhHF/Edz/7sjVSnZjyL9nMNh6zi8x0Le0a7UbdOjp8xSitHo2t4U
dbF09MA3I8sZfMCFbOe6PstIIQAR7HohUvvQedJblzJ8HZlHldPxBGNx4BKU
4j3cwFKL1plIdTMXmSsMbGN/Hukrc7vzGjhsNpnYl15SvwXMt/RWY7k+8qqP
GakFPGvLV7SlX5omEZpNpW3FgSFJ/07T9u99hCW3xJT6ZbD6PxHjYvmr+ZfT
7ApL3fZMBAFATE5u0s97ZbXKzGIvv929+yXFO8ThMzk+sGySbBFRUnhlzm59
1HkCBdojQvZR/FfBZMa8rvSCM9OjDy4xgzqFhUYGoi6z1u9DQ/VdEkNZGPCN
VYdX8RN8Y0VwmxxO3Ewa45zVdI89FJpKpJBg1Q0NhB3TDdHoUohzDUnY7n/l
aRIllRZEj+h1nsK+UifFNFJl7SAjkaQx3DMwb/85ka/yeLwtMBbdD3rD8B9g
JgVC1KNx4Pdmb+uzFm6nFz+nXpQoiMCnahezhPoNByMqmVo+8ZoQQzW0ej8f
9XwSZn+kB8A2AUnpblPBfWI6BzM6gvFEggQyAC1z49/m+a/hb8Dd5Iqj+pPt
EFcMu478aAwWMdcAODgIm8ggXN0uyuwSXsswmZJX9MIHpNcSt5uoA4oF1Zoj
Y9s0XQDzLfjw7RS05U3eQSei82+ElIg/6CHUuR5zAX69GD7g546Sz06ZXtkE
j13GgtZ7g6w4vzBUvkOS5WZYTqZSjUhkflNAb57MM/lz09IaPx1L1oiNMdpq
HZpded0CW5ahk1H7SUmt8TXC3M65fCuoxXlkIM5vxPJismpdAZ5ZJCYj9b8p
gqmK+OALgFAp2+yEeAidLCkRYjymfumWLqf4yiiOi/b8aRsUYAndsldkk3ds
KstKO6enhpoU/QwaNZL4uoq7nwlpBXk/kXEjr+9MdQ720W8BsQBxCQJxYy9s
yGF4XioRTRwPSGo6juc/dqC/h6MCruS3RGb5M1UhNZzz+6wce2tCAdtrdbj6
+5TTIIOfDWeWZ1mdB1dksqDO71v3YWYMeWBfWmD5Xw+LTLgGy4IaeNDOcPxL
J+K44C/mfSGyvp4cLOHBS0NFf/0fRFuEOiPjL2cNjCw4LP32dop3bMSoYB3v
HrJVpGpYADqx3+3twcX71d4dQimWyw9mXzvoUwsDDrDPxkjXle4pEJ5Xpjbg
o09JUaau6+MJiWd5xSTzQ/3n2gWkVnabrh770fho9boi3npeejbsx5Zgg5Hw
2cThJ57BKLkD0UYGKTbimDGbHqmdRR6QUOIvvknYsCjzVg6IBRoQU40tCHaP
9FF/3hJqhWXe0BT9DGuVrkmXCPdGwEW8MjQqR8mJdOn39Jqw4AfCjdr241c5
uguol2Ep4FAJXJ/jd4Yw8//hgS0rYGqUAuP258xiKGwtEsLCNpRxmKJwwuyQ
4jKDdxg8JgzLRu0tghJUAiRj6Bh2C8WCDz+r/zmupoR24b9DVmX6/oy2W5H7
HYwpaM71l7h0Cyes7F5dN9kgSaldTy8TdutXHClxahTqQbOwJ9qUZn8SmGEC
8S04e3292+T/B6jzfVmyELlV2qsQ5iFnlG3BYK4MPSOGh//SRpAvyKl8qp8Y
cEKorYMQjCSga8nH3wu4aMQKy+eEzgKbgJBlQR6Cu9wxs9G+vew6riz/R/7H
ycYC2sibecxQnvwBo8MlRyeNeGgismi4ggyx9qMZ6AvI1I568kPOtdKYPBw0
A+9qHBRwUZuODSTsJWP7xuFRQNdsTVKt4srgzQ0DvCrDfJNdUjuuOKwfBah1
AW5pck5JvABimiRurJEZ8snVZhp59evNjpGB1fglfQ74vGJ+SNNxyplZCp98
lcu+jUdReuA0wsxuiJ9DGmcx6q77qbROvhxGfc7Lcc+jpxK27zljIMtoRmH8
K9aRtGJHdDNOL/C23TZ5TarcBiKrAEQtjr+FBRiihBR8ln+ouikvmR/ZfaTO
y6/F6lbaDO9k7zRAXsP/r65YT6CmQpyyuF24h/RFuIOckYLTze5YBxfREH3C
g9km62fXdQ5YYKXg8+TYp/jw5b8oq0lFv3Q9s0LfPbBTYfFjShc7zd2B7CEL
4HcFUT1rG0O1WCGtaifpImsOlU541kWy66NNqxuF0T9RpKFPouIdPNqEbO0w
UdERcdZwNyZYduMc9bo7/YQfwSefISdv3MnYg0NI0egXEMPrDeGU229k0d5z
KQ/IHYaUrsO+l/0oJBQT7f5k8RjrFa9+9I31RdCqPcAGmUa6SVlN/joAZb2U
jfL5/j2Y9wqsCWJLeuKJOnqFHoWpTB8SnHBt/DsWH9hxnKWMp1b+TfbAg/NH
/LSjf8MbuwzzCDku7Hu4GY1tLuVh3+ijWvu9lQiZRumFE8XAFxs3AuZq9Qgs
IKBs6VFkH/nsgIbajEnfn4gC0Yw0MamMqicir7OrFSdIJmMEfccpE+mqWVIi
C+gYrSS9qA6OQFBkdTISVJi3efS5QydMCQoq6gyLrbxv3KYXlJ2NDX6pPiiW
LtftugPwsxiDubqQ64KR0z4WksTfcPXmkfgU26V/GM/vqyu1kgFlmLjGCD0b
UFq9pSQcwRuMv9G4qMzVLec2Ow4zU1au8WQ016LJUB0X76+BP6F70CN7gSH7
Qq7IHV8zq9TAj3igNTlLTD9w7wlcRGsSOrvOzVNIsZN6g20rV3xLgqHqHQ0n
AfE/88wn3Xakw9tlwgeKyWWqnhXYEkARz1qUI2pAAjvVXMKM8AooXOEs2Hc0
bn4KBhl/zwTuIp6SHsVK+Jb1nZBjedRvwBCCOpi1EezED+wFGnHlBWyVR6xd
ppnpe3rp5QEorB9RUCfFbOEnB+ClJFWCLf9ddY8GX4TqjdjgRpik6AI3JwUK
BjXv1oFMVdhp8uSxpukH1KlH6M/q+i9kc0Orehtx4iuTkuZwGV2k2j3Kl9dt
NLY30TBatwdeFdrnXotqNYv154ZEvhPQnxQ5BxTeWEysZ3dS2HGljCUT6gvx
K9tWSdNdYrBET7gbk2nYI56byacSbGNWyMIVrTx0f+6qliwRAFC5aEKepmXm
OjWG7vWQphtO7q9I6APCkW795g1urRJGUzRWFFCcFkcunBps2VLg9ZzAVack
gE9USvs4FDPdEAuvdCTuVWSkhA5ui91YT2Dyl+5Lcqzo4cUb3MbYnl8jtvMz
7EpGz+Utmt28A30gyIsc+jkcWp4hDFWByjaFBQBMoP3HOY0+NvdNKn7UPYrt
8TQOh4vlMNSyU4Yt0vA6fqC2l0JJnkeGLb8OuCOn8/ixYlkdL1aDFSiuBe8m
TKhiDhy44UPcUwqa/DxqL8ayIZeSgIqylWf0g6Jw1w1YQQqWyCwzytVV0j4q
z3Bd8h1moYBN+B8GoOUrpVCgYwZ86YAQIL/pMpi+ZQN5baHrEVSICO9LkdpJ
t2w7+3lJunj/B4co2Mnk3Z9KT8kY6cNHZNuzP1TipOYpGguMT5bAxSwj4gFJ
0NnlNGgbbXr1jMoUH/nq/L4ajRFQlCggZEWeQ6Fee4x3uoAE7WoxCnV83LCo
LY7D5WYiLlnPLewsTyz+ZoErCykVD3S2jjhW9cikY0krr9ww6d41q6084wfu
kcdsHDmp3lohpqu1dZui9TGldiU4f1i4YZfMEvZVkU3V+5UGAkbYEuAvsfGW
cYkiiYjz0ljP/IQPnsp/lALj+/B2ehSxdILd0kZrAfw1mzuJb1SaE5YOXvnR
il/VJHt1VS7FWW+OVmapIITwB8oDd3mTfWQWwwl0b0//GGMezTedfIODRf6F
0fA7drpR10IjBy6yxa/UCgWLr1dp9PulJskyAvz57tjc2D0ulvEYcLCGgCx3
JQGAGWlWcOZObVZYeIcDe6t7qt7LWFOwWF5rlhB6V/6JAdfU7ZaUxoPzC4sn
S8Lu2G51E8i0ogetphgSdfQV/kwdSvdl62wHPsGWAjEHPz+qqdSCF/TPOLqZ
WN05YOJZ5UPe/ymvbGWbhmFgN7jnxWGow0PNxQ1kev0KlfoqliXcF4C6wsgG
OCYevYeCCyrYbWuTIdazftTCGT77KfnLpvgCaxGBtKdIhcK1l0k13JnODewV
bnPaNESK54nDbXpQFLMZh+f+uHDdarV9RfAWI4lTIEPP7AC6apVrq7KtcpKx
l2cvvs7UF0L47ldumfcHJdSxQqybgt5ylVqSV+eoozbnm88nvZe3xXc5tDqv
4QFBRWWDJNOoJSUYBtJIpnZ1pv/JiNk0+Rtxk+gQSrxjIX0MSK7G4GSynI4O
q/glyNn3nUrInXEdUKviPlMzSTGXxHoH7qxIdhMAkwD/xWtJ/kXE0p5TsHb7
6vEf+g91I0ces8raUHVXsaPGqHWbzYjEknR6LEZaj9kSM7cJC38Whqd56pO4
wT9BwK84Pc66rvHkfgOqwx/c4y/r3ca/WS7IuNXd9RrOT957hNlP1Ytn4X/B
7lCv9jnb4jyJnfkjIkx4G48Es2BrJaGWd2ISwtmwr6Y4vHZOxRbLDQMer7fm
UkqRa7oilyYNBG5r6f5ukqQHrAUrA3xImBS9wXavTpqmF+2nZ2MeajdVkXfX
aJOvdzByLv7TkI16uMokTEzZcUYdG6vJO3y6Yg7qXPNP0FV2r4u8yvpLLtzc
d2qFM/yat9A72488lnevhrTn2u0la23AcEaN7HO6kViPv9xzzNgPd952FenA
H02hS9+Zyev9rfaO529mIKioH1bblNVeLuqnKIQ5ynpRLX8lCbqmmrB3VR8k
sO3aLhna22KqpPqvWYYmKB4sgwOY03SY4Oa4WCpM58bhj4oULDTIOHvbzVEH
wZUu/3Rb16PzTBKbcXOTiIAITN42zq7BmFFWhJ/JJYxw3Q3Ykfs6Rfhy5FDu
VAcGmSITIoaFcRPr5uaDPyAGYWYBN/Hc5Cp+kGEylSvKnl44Pr0H6/NlJ1AM
BrHdZdOIQelyxkiwA+W8eM8eC/ELtD3hQ/sA6QogQSDSVTwZyYEJwtYOMu7+
YsTZ9JQKufLdsBoDHsCVtauMVdCICNoabAYB1yYiKcXbNMIMjj0N6C2F9aun
sDoiQB/dMVcAYVNB0zABc4OV1OglmKCW+JxShCmjXNxWstrGNRGEYhPX+DzX
L/f5XY4IQXph2fXTOINMmo0bFNqPP+U2Oz6PcsJ4MMgAyFPrytQe84B8jzyt
Ol72uCwFxdYvytm8ytrmqQpAiF30+vdf6VogykTsrNfHs3bAaCttKS95qh3k
WQl+HZilBSk7TtC3V8gMwmtb0TkMOlFFpeXS1BLUtXfDUQdiSzYlgI+7Ct3w
5MWOHnOkTmv487qCKhLVCh6hleRbhLERUV8ytFLc/oLiYmwTA1nvNDG4TQuF
GcZq0SaKmeMAwdaoVWATd33Af4Q41MkmXj5iamOqWjsAu1hqhLI/Cm5qmIFW
qSV5qhS2EV9w/fWbw+KWjSoZohiC3pYWTBHjQI2q4htKrjixoSCocJYWQhtw
9sFFDRVSuw5gPbKx97EnserbI5KV6OgltVTFP0mEuZjFnvbAQhMQWadsWamc
hYQz1VCVM9fL3IMHH3QX3aD4ltYwY/u+C8xia2Y00HvNFz/c/jP3YxVPAfz+
cab468E5h2MFvJLwVIDh/nu3UokI9SikmlhXMMQmUzt8go+AjM2W5Ssq2dF1
qniGJgAuwnuYC8Ct5bJug9W59UbBtaCZFKr9KTyurh2VMj69bwnPAhX92Wf/
EXETI7eeKdw6BojBOzgpIZu5WG8+Po6KYY4wH51HQd1w/CqBK32ba/RS+tIQ
+G5QpmaLw69LDjUqLsdo8gfWDMaWIQgfgdGnxiWoPH3TYKFCpQYWyMsF7Mru
OgCKpVEj4PZO/xbr26c5Z/0eXKb0Y9CROdqdm7tEFnC/+rRFTmSaLxacFQK3
ZP8EeUg3I8BiAJ1l7iWlv4/MWFC239crNU+gAP9TNzaS4xoMNvfBqyhhroGp
e7t6QZ9+QbaJCRS/QS7mwa6h6aOBz82jjfHdxybaLyBnMoXxG5Lxz5Ok0GQL
Sudog3rIwBeB0zq56bFqlqEZ2IgDkI/uJydg3I1dRbCQOw+GetlHGGQej9fF
Myj1sFehYB2dchpH08DJNQhLHzgMOJ4fZwdbKxmzUraeTrrkD+8m3eYQ91rq
UHFe/d/xjHbcacoR6+yHo2M8qzmK0p6wy09FH4gXpeJhO0TrqdowBm5F+Ev/
y5gE/Hqm6Re2WpeXcckmlbZzwxotM2Dphig7QLFRqx4d568vkF4B2+iDUtwz
nOwq3YL/aQlFZ7z0O+nP57Xsp7UOfMwxnVYZJU12NK5Ki52Ydy+RQcd6RxKY
vUy94C6slYC2wlQoIUziitfVK0o2UDz5MJr8REAwmXVbCHLG/AeWGZqHTVd3
d+FNrKIjebkwP808K+bUcgOxG7MEK4ixp6Z0NfhqBSJx2MADCmG2yFlvViNp
cVZVpD43YXKq6GURE36PzK1tSaxMhjhNkrtKcGv9AfaAL/D57OhBpdv2rgDp
Ck3lXrCzudQ1sK53kmNGtg9oe9GvgMnImJWIF2yGLgHtFfxD1S8JveJlnlE+
8co8Iuhp6R9mJxcvWlKHKvarq52rjomWoeX6fNGz3xJklFW7ecAGc1SbLsz9
niOMDvpu2P3q2Kuoeu7qqNYDTtLGnP1cYJ2Ty+UyY+CoKeJnaHxTbjKn3gFJ
QHijsDUmB8Hb7UFrLB1WfSkXIiEhYeUfaFZiKxqjyqpyULa8jD+Y+hIBvZvX
cfIr/Gylh3TrDSj692NXltvFtorh1qtmuL7ve5QqBqSz82Wny95iCeV9vQVL
nY0n1cMabXc3k6XNaOLC8YiALl7nU4NDh8aqcME4Z8vZpR/cLuoXZNzL0bik
Ugtc8seM0Y45ujbGVT42F1nhx6RvGFs4cZXsgofU0maqkDfx4Y0tCkPEUhmV
i22zvlZyHi6AE3Mj7SohWMhb9FRYtGECBTDHPwvjWeEoKtKUvDslh4FiDD1A
8+Myq8y0jp7A2q7SE9EE/lYwi+mZTi+lRdLutLd4AWKdR0/a7ZDhxuMdfvH2
u2Purzj3uYSDS2SwI0X8Yf2aa6I1ve2a5focWi9to6FceunqjxklJ6VynjRG
PjdNM832AJcAfgqPOd75uK/NYwinspmWpz5bursYwpMvfDBPhLQlKmdF5gv1
gsSx6FftaXriQ99D1M8mArRqHrcsGen83aiP+xIRR05R1IJnphJjMIyqvxN6
okOGAMDvV7DsiDCFOZ65WnZ+khXCNgVQz8M1v5QrUSynMpWnd0wi5dAwkAK9
aHNQueJS5vTaw6Sr6RDrIoWH6EWia+GtS8dMPOpSz1JHOpsTikqi4IQ5oAEx
bWtwa1MHCpTcG7/U+M8Bm96coZrf7nlV6AmfqNwOgTd6NwfZ1E642WjVRPQI
udrZ2+gP7dv19tN7t74/1CgzBs5dFyIFB+OU1aqYL3nIVtU+EkpksG3ARo6G
GRQn7QU2YRgwMlkt4uk9mM3A+CDbBHq4mdke5efh9fnAMse7zN6d/ErbH95E
e/F1gFNLKz9cTvS1qwcQYJUk16Kna+wpouR6lyhCdH4G6oe4enC7WbHyfTu0
BrEP59ATUwUKa8n0ZFneY9ZxvclBzUA/lfDb87oqYlTlV90ZvdBI7+sgTxG/
aCNFM2iR48OR0vNrmpmK6pEfo+E4WzVRAUCQdHYxXkqPmk2flCM9P9Ke6MQL
1Xu2h81pY4ETNoEI0+Dzl5fz7zBx+pDiTm2qBzJ9YBzcB8HpFkMNGt//ZgjL
44WNC7fnH03Kl9iaRyl5XrXtqXGPH7DCtOe5uKXBmge7MR4HfPcqvrJMqWLx
BHEEoXB12xhefccDEftOZPCLSFp9v2juJtkmdFFzTnJVESoFQbYqI3AnPGEt
wiwoxOE5iseM4phZk5mzouRx8GTItwY9r1rDq0za7e9znuZRKDJtAyMvzrA8
oW70ytm7iFYq2lx1DZp4LK/JCEsQOyawMkuSm7udEofdACenS8leerYbtR1k
yJE61eHOXS6mNDedDyG/65lnYp0W+RR8qE/MUjLtViVnMdPnuX5CaGC6v0ms
k9H3m4ekahPVbkQs+xba9/cuFdT0XgeuRNtShGs6wSKJaAJCW5ZjYSjAcN6Y
ozv1y/eph7qaQD72vnzXvTHLXZ5l1qtsfv/TxkkB4mrVYSYJ+4X13/aOH3ug
FqPZGjvz1WvejQIqugHqf8lwlq1NfTMOToqlRVBzSwvbO8WAUPNlWboJRDSe
yUoGpwgTirnLOPTR/b6L+fMluaRjA/vNbcvP7iNzlGP6xK5Qi0QBxqzfCQh5
0j/ZQrz58AlUGpfPIKygMVk7y6MsCLICByhziL9TqJEmLhIbrxyr4hGZlhQc
+LdsBUWTi4s2jRBAFHx7j2/zIvjDLcSwHyBEb6yHiLEZq1zLvNq3vF9Nsu5r
V5yoVch2H7GvCAWuKH0PzbLOc67Pj5CU5RxWkfHKECKG1bcyJRUElMXR6lYJ
5ji0wOAHGWgB5I3fNlblJ53aHwG2Cgi1rUiSu7qVxuCTZUPdfD8PxESM6xQF
HwAczCeB/J9dUkNrcsim8zLdIITsslExBtEMmYnLbz2WnTyB81eXhWNpuOM4
HWBiOU0x43o0e3Sq6nDNKQi4Vxdw/GgE3y53NjPROC5xjKg3vcapTm6nj2YS
z+dJn18Qa+gh8aZ2Chm4p7+oFgsGLFI9yuhGPcB9oftO4FBO/TMJYN9zZYzC
qTom4DM3ZZpSFa9JP8WI6jnHVMU7HLIV1hj6lCR0Ls4teeh56gm/44p0MM7H
RsrFrapZUM5z93bwHMl82wDlx6fsGrN4P09tI9bnqdUl2mTS+g9CxhnkxMQZ
DxpMScV0HTJS7GcWVLRThAA1vjFx70/WC0LEArfRQSp+8DSE55uCfyhtd8k2
KCYVZRdJZS+cEXHNodQYsO/MC8yctj4yH8Bn0BSeBTnDCDbwoel4O187OL6f
0xRzsKmwngTLZcOO8p9C8KoKMUxLAnPV6gr1cpTr/9oxGBTyTGMLf/r1TQDJ
aykwxH1EqUdcMJU18ISKDzGTNLaIB3EdLE4spF99Kxhw3Jfiz5A5IPJp2cSa
V+e+VfXC70e5yuqyoo8W/v64TAYTXheUSZdTCmcUEQxmr6ZI+zQqVrm3QO8w
gvKIgHvbUmhVmFBb1JeDsV0/IZSZRjRYBFrDhrBzo5se+ANXCXeFvPZW+x/f
OxaZnA/iNpUYFa3IJvIrfF+7QdLbe4VvBPLx8IssoJzj3v3jnrg85Uj3gj35
FG8IiwsdxGVxTPpqc3qJDQyV/qRSgWcpNDO/Sbx9lesQqHpLyRvIrKwfukRK
yedEGh8G3Qwlon1OTVfDjQQMhUaYmLHSCxr8V/gyztlVyMtIPOkqoD16sICG
Y0LZp2oI0s5uDnU5YoiT5MU0W2Mhs+rfhNA9lZhAJVn90R+zykMZATPomx3l
UnmtPMC9nr0jI1u3Yu51jFSKVmeEVdakAlNu/knNF0xFqzSQorkITLJ5Huda
p48bVWtm97gSR9Vfb7CKF3K9YoS2wgZ6r827az9Kxj6cgf9KJkY/ZLPOMhlL
oEnHR1LukMjcLzFxYGvK+rWxuPLsucPi8Wj8Yr2+LYMOOFyMQtkZ1WPZzDbF
PGh1B+jHxdMWIdN6m8KE5Z9TEz+S9b68XPdABRrIuaQ3OitLZkmDmg6N7V8r
IAvpMot41eZegeHYm1QEUcvUPtKDREJ2Zc3+Xqt8dpXY3pV9cgFInah3xmi6
Qv+3fnhNfzIyP9wiMdozvqh7RI+DpJ+I0p+OiKwSCaZqguy+CWAcikYwRTIf
erKFGhWUkI8OBQLbYVNTMoKeIFkrJP+e54o3QlYhLdM+XvkXmvAS8Eh+9RA8
d1JEa23nx2tPBA68jLR7qzTki7Cp7QrlnsQnAI9SIfgAACfcnX9pYYB2pf4G
z5tZa5HKotwrsX3+/JDdN6v2QGL+guLjWVNEDtp4jGCWjwlHaxF9KOooq6HI
9dYR69o3jwpN67mgUTQKZwhedyYF5v7QY9OhfBAZfHA5ZzoxysH88XhRBsme
rjS6SoJ7HVSv6Tjw0hkbw9gZ1zkjEP9PcXbyeFv5T4htAHZmmCP4jodxGImV
iniASXiLEYIIpzvp0Q2kjWHbgNhL468Sk11ww6kt3Y9MId3Ar0XLOGcul0Rd
8czZPFe5jzr4v6Irec4pR1VoaP2o42/jX+V8d6R1jOTqSveMif3EHt8/b6tm
P+B/jrZ/O+t9ffMmI8rly/Bb56WidB54Vriedc/sapjNq6wL9WAQjVMKmwmf
uzsz6lxaX1yqEeeeTSWYN2wNUJmFRHSc92oJf3CjWeOG+03+KJguRxkNVDOT
lpYNrOWzmnh7IC3Ft2Rgg/jb8zOWjvP0M8mMIlLLLmOnqW7JMt4MtpN909gE
9SEpYfspvGVNKsH4inB2aAGzVeO19rqZwBojEKtiI+LhSXJFPk2GaN1SYYEM
Pd6QSuFBRnCEkf4yuJIPZnJFKBFWtQzJsyCx7hDE//HxFM1QzUIIDpjgLCbk
n5uYN0b2olZE1QFWFq5vjlPjCSyRc2reQbcVR/Tzek3Ia811PVuOYMjq3R+5
qQvM9abqf3E8Y2vpJlXw2OopIm46cQ/ed2w8tx3EUqnCTbNTORmtVv/KfXOq
Hu5HDV9Zp7f8gR4uyi3s+tCwc9CbLSqPXgyPsadg6v8ARBk6SRwrPnzlxibV
zgwIJaEXL4jbq05Mi55ENTmBIZOnwlSCz8ai3aligjwW5dkq+zEaB8t63oeZ
TuFIEd4U8t3UykFiDgL+CQBxGHisL/AoUN8wCXaPXc92avctuJoxWxHbc+Si
hYOIje0iOiO2X1an+V4URcsPFbS6sUa7Ar1eqv0rna2IheYxSG3iTDJ2HAIF
2mumBA178S400h4zl96Xin2rOvPW/5wO3kx/uob+uaty11hgt2r39rllCcz6
2RSZym7M/ZfQdc46KxhegPiXG4D3JGmmPR1Wi9XCT/raAu6FaFsfppGmzDuk
bd/MBSknG1wy8/VyQBQNLaKJS4a3xnU/cwROdZgDgBKn3lvQ0kPwPGqV8S2i
9atVGuinKBVXA/KycSwPTOCciJ3p/+TRaml06ULcfe2wGpLd6wv81FuJZ3CG
6Hj2xmcQMGkJLDyhqIt8cGLpv6d8IrNDmizJrl3lC8acyn/Mg/wS8M3WE+Zr
rlXcj+K/uT43g9QDKgZreAnJLUBZZelKk7749GsxDtPUton+vidGFto+q+0d
DUSNrKBVTxyI99nyZIY1yInEGXR38rNJvdQQG3n7vokyNO+hmLoC9M0g7NN7
ZC9tm7pUWMiO6q13ugIxxcyrlKMyJS5p5Zafda0Trcg/KrkHiEih2XXhbMU8
7pLTnwsUDz7PpmRm3/AIrzFjzq6SYie15xl3cIMEEMrV3/h7mF4+Jb6uuMoX
F4yz4PYzOVfZsotQbBt5W2wyAfkgzex7xWeIcyPewpfetTWe/kbrDX97S1Io
bvpdE8lKi9X53eziV4xoylIR+zIFWUfy4osO/8qaKSEbtuxxeaovgOP/b+Oi
gb/V4bcTa/KHjIPCJSQKHHzvJUgoQzzdwo/LXAWRlwYNzRfhC5XHKpBLRKFQ
Wj3hCEmVLzBPbtSR6uBD793T+ZaEwLzhf9vudn6dYeyYj98YqkPOL7RYaPc/
MehAnfJh8uhN/FEMTfohSAIMzU1vsm+7vPJRrnQMtAhgTPCSCTzx+EjhNWJU
GiJOwdZkugrGnqVp/TfUDg9kYQuVCc3eXVgIMZGOTBSS/aOL90ejDrIKWVIy
b1LkjL3uJ+ntMDlp8KhRl52Utwg/u0D1akKHXKirDPdQ9MC85lokq7gfYtpf
5/ihgm2SA4Uz/Z6lXZSGO71O9gB44uS3C1Iz9IfO/aM2CGIzNtuO2apNK5Uv
jgTAQQHc894HWVSxBkih30FyJfumUJlheMIly06UVgMrTrW6XiD+mYCa6K+/
qaSfERZ7ftVyb5RzPPy6xFrb5otUO73ATX4ITznertK0fBLAqB2ESWDx9qf6
4iNzyh7/fc5kPoON90y9ntmH/QyHvwOVwKtDxx95EGd+oSKM8NVP+93YWLrk
O7oRUevXXszkxykMG6X6sMY37yGW3XFmaEUxw//MsBo0QdMs5mz7aEhNBbqP
LK6/F6B6+hIRCKkbrnDbGezcEp4A8CJfrQQvkrXOJ3kNynYvGoSguFdQgRza
40quEoiAenElSo6pWFXbkzd8a41QEYaVt7Laqflu5JmFUnL56zU+faXMcgPn
pup+rMa4FbGVgv7HM3X3Iq2DXr+QGiSvJssLO4OXuaEnw3yLvb+mmcM7gj0Z
8iNUXz4AQ6GfYHAHFgb/8EH4z+xtCi8pU0CySv/2fGbAiwlkKL5rn95e4oKF
/+SSHcMGq3yJBDxQJEUJDMJuGv1HIYoQizoHZQdq9HQBCVhN9WUP7rsDo/90
R+xfHxV4afVj+h4kv4zILXm3HnjJmXMYETpIhQfh4/yhYJ6rpmDFJmOFF6y3
OsS3lzMghLVKMcdnGtJez1CbORHDX2/bDzUH/K9wS+LMeif5iV4IkJKgllFH
4aXH4ylJdFsQI1aWxkjMdUR7CZhR/ytg1kgOy2hSkKv5YeeqhRg+xJuVzb7a
NVrToJFN2UyUb9gmrRV+0W7+/KWEdWwvrZrQNdEmxAtA465hvE8OQfpFGOKt
Jf6wz96/z5uXtNDkal596AUl3tOKGDoCocUzfMCfvSR7IFPqQDs6siC43zI7
2YqlLdFQEm2JflwRo9u+b6Go5L7S4n9BxD16jSYBS2QAHsTfIF6kwcWaxwh9
kRaDLlEjh7rx8r2FCp8mxCZPkOd2Y+x9TdPi2D4t+UBqGTDB0XE0Fgmwc8XL
hqpeDj9bUlbrUXIsxaI020nSHykfgd6XOQ58aTnbc5/Xb7gngGZ2iFL+hRyN
XFqfhZDMJOBPkNpefZyMIkYvjvTI7pJgMpV+KUxu3hWBsAi2WgqZ9vH47BNO
nQn62i6e1bm3MrNwZ7MLi1uAubRBVhxWGqVSUR10Zh+kDU81UF19X5/9uoht
najsJ0NZxbjKXE7D0KW91lQoJPVoIMKTrHrqjnfryiZWo3oWaxeqMyvUNGhZ
VhlYekLEVpFZ3EXbs0/NLS3b2vY2SIb9p6w/pxkJxeiiVYejy+Ky1MPNe2mf
HJsf8h2Q7lv5IszUJYuJmCmtr499NLW+BKWyz4krCyTWyTnZjjJfnIS2N92B
KZun6F11fyFtiZeDU7Guv1Nv57kFPB8BZnpqqHmmnoSA9WtGhxLXPenqgKHP
j0/GaROjbTyuvrE070sOcmLb+r8QY8y6y/ywHX8sMKdPXvKt3pCIOLrWTMNc
sTd2Wznk+C/bKfjkdOvSjmKsT5t9mTkAfPo5YixhBHSeZXACRa71dSQr/GiG
/XR/lwTxxb24SWKl1i+RkqSpych7f7LKvRhQtDB8mLTbBPUeJODn8ByzSX9o
7VJ0VidhePnYQJMAWRJ6w0aBdFQhctaJgn02pOdD11XWA/WQiixj1QKfhQ8z
JDwtJU1UtQa8YQD5BYXVCjAi40aZsD8/rAIqN8ruWUIjl3BRmXOyqnhCXNgb
nh0Q5VF48mFMuSHbxNg12RJ8X6/MgCLO4+zc8Q8BEk6PjIFInxnEKx5Lqkpf
E39GhRKkvtTvLDWP+xP5EXMKzs95rqV287YptKvAtXZIXFFBSXCdJjiyFPKF
tt2WmmhCCwFZD7VNm9O1ykldB47wS1CjB8/VQVYzc8a96633Ncbks/KOlla6
iLMaZk/XJT8FCPKKg+cIPwBUtMbopfHQ4di0WxUhhObYDud8FJmFW/DZe9L+
usk/7sAgCzFsLuYVi7wJBcApLDQBBmwBGhi6CBgRDkCEvmOkxHKCTrzAgBnP
OSVt5kyPEBFd3teICLDEsXuSSSLY07PS+Telc0gEbnIZ0k8se9sx+u+Io7RP
74BbdcNG52Fd0SKn6LQxh8dOqp7vc0rUE/o9xSkbadoGnsK1RjNVehGSGdAS
ENKjfyVVusB02ltO3soA9L5HBzw69v2TJepAHcTRPDzJPoauus1Wzr2fh9hP
SG7a7Mf3mK7FqxC4oSUVVdpgVvIzuPnANixVdvRb0egBDAZW2dduT/TYCKmu
RcgR10S7Qn3aopdmCUCdrc4+whWSnIM8rjl8DA9gunAsEGVUq53lZFmqJnhN
tJ+6sMw4BIrzw16+00+zE/y0mUCEdENmZ5X4vhmbR/fNA7dh6ZJU7p8JPDS0
HlKyB9b8AnOyX+Q5CO+glDuYY2cAeKMNDwXPsPhr25g5Fhht3C81jvF+HClP
msuIkA5g4wrE+1IS99Qm3AbSZDdKj9EYZX6twRADk9VelJVWah7wj9iXr2cb
gzmy1VYoPp4Cbh6oEGg5jtb2ykt7Mq7RA6mZX9rVFIjRMQtTdvpu0JZXTTVB
SEJ+bF5cXinM3tqGt/gdKaXoiDTrv2VJl1mSBk8zkVA6T2MPBUr+ZJM2MO00
ei7Iie5ps5jhkrHyJqhfDyojDCfvoPKrjyFa0CBlWDcP5faAsPz/7zZr7xep
4vNJmXlzmf6bGBJp3csRM7a4Trus0Ui8ZroptMbCCBb4J31uCoZFDJZFbiFo
cyJ+YB0fVQViKi86aUqpICQvhXLBju6ZJuR7dLcUbcoUoJiHm5g/ZB3TGv/5
7u+hanKH1Q1hIG6GR4Zm17bTHaroh/EnfOhzwp/k2TQ0ht8Yv4+Yq8s5HaRW
d+v3xQTYSoKoMEYYaE5HNt5HgU7NKU05Onj7ligDymN/gUkC70+HiwNzvw8X
NlvXbrFwof/RZHslLpnrF2n+uZFOfnO7xZ1lNNtq2KchA6Kwta/zIFtDyC4k
2G0WhRROOFttr+asiWhdcRp8s40hf3Cic/qeKj+DhdYlG2KouJnHjHMZR6m7
p0CGFQBvvulTjl+KkjAbpbESRuO6T/WPZy05zv1I6lmo1T9oxPc6SHef7zaH
LWl8XyuO2+1BhnXn/wLRRY2IGoJdHPWCldDmkwJZwwbc145fuEVfInPME2Lr
uulSYgj0P9VyVjQHXIXGWF61vqF1IaDoD+6PmC9QmYPuFuu8UVsPHQJWjVuV
0PqErUoqfYTDk+1NiGtOwMw14XjUwDZ97Hrbx0kI6+JxL2nsnT11E7geHlR/
Z+XivOvJkSmHSy49sSyn3+A59ylhsWvdODoovlZNu0qaqaJPAIX+uokz8iSq
BRg8dZZ+XYYLAZxSS1adFaDLgObl83NJ3bZPwY2yab3AWN+Awp9R3JBglOrM
wrAyAWqdQOKL0BjsJNteoV04DNoWnxJEVK4XiapBp0xvH3rt8FRw7NqMEate
vq9+pG0BDP1fF/8NfhDivd4RtC/Ih8fNG+u18yFYLwZVTOxynpnO7WGCVM6d
w8TTmpS2mc2Ennaw3+GO+XffPfTit0TmUtytF9cY/jBvMUmgS32SfGiNkGif
g7JyhZs4KRJLoZUJIlR3Mb9EUSBEcydilssQCuxGONo8bU4f0Rn+cZ+i1beB
DMv0uZHXLMtwWmP2JZXE5NDA4g8tvxUtrF8nEUGenqbNKjpw0omkBUZXyL5g
u6g2rAJg0fErWvAG1SrmiEsn6DqNv6ghPGHxyn/hJw9S1ue6dJQfVYkAp1qb
TtAmXbWGxoRVvr0sC3GknzCT8teQL1h3ztXvcQHbZWJioiEYbwjKervNKdL1
0h2HmTckQnw/ORYaSI/LveWeGARUh5YaU0EF8vAiBpiMFgBQdPd/KXZBqbYC
X2aFodQnsrezFVHIjKli0R4PG+lXInMuX1VkiCM6j6/v3J0A5Wl9AqpAAsd8
6uKxrwn96PDaHbkOfVPHG7PpZd32Um+MuM4ELrY/Lu8jVAffipoNiusjgwtO
+6zfKGaXzw9qjx2U4QTfpaw84R0eUlloXdkqhNijAt5STYlJ/F8QwowDYluF
WKsjXmPM5MEq7MTT4Z0vUO3hu7fksT1421N5h6FknVSoKq3Cp912wtF/pFc1
0FPP26SzRXb+AATxgoAiIVPO9Q9pkKhVBNkM2ksgjGzLXVH6bLs9C0PFRbf4
rtyBf1jLJEQ7O9EjthaXw4ImzN/rk8aHoy5wE1ZbYBiOfjyvuEj+KT3kKffP
dF4CvGbuAeAaZVaPDEwHIIOXTHZi8bKyJL4LzPLalZdsjbP7vQOrZCeKjK5X
TYCIAIyMb/DtENvxeSdoIO45Vcnst87wf8wWBJ++3npV5Ewdt+l2kxmV7bF9
OcyzPsSVxDwQoJ0oxGe1pXMi29SgnF2KUIIpdicRCN/qnKzhcEJKzfS6vZ9G
S/cGb9CHf4i6ItN4kxBIBCLff3ONM9mcr/0cPEIrJVgyJWoGNiGegfh4VI5Q
JzB06VB8txn6m4RZPFH0ilzl5ruAjtPDMaAOZy8tA8g7V0oz1zEoDdZxhHy4
kpDfKXJ0AYwTYX4zdxb9SHihiciW4Ozc5E1UVGqUvtCqP2Akx3t92aiD1Bz/
MBSNNaXE8wO/k8apFeDKl2gkaQI7EYCEP0tOFalR6a6CwqrkIn1QzbmI0jX0
gL8qnbqU3I5QFZGkUOJ40TQlBakgVsRSc8eZbtrzgn2daHPflceUM3gVPR84
ixqOgWEfMtKmIrKj7KFCnSxoMiySu0YiKeK7IRjCb6IsRmId06WPJc9Pkb/O
aVPPhB699sqWhFsfVX8XDEpq0V+jXzYUaWvMRSPB4PE9Ou3HUb833UhuvZC2
gEs7k6CsClLwYn1jL7ZW+3z2XZO5I8jYOwgvHMur9y4y0WBAtQMmBbXyRX1p
a4xwo5Af698noXTNybsBOj1ukdiyUc+oBqZTKzf0GEplOopKmUCgp8vtDUjp
TtfyC7jGqScZRlxtVHkf7jnr4gM0F3lRm9GEzZZu0xKUvF8dSSbKavhZffLH
K3IvzlgmGKnOcov9V8cE4/DG/DAyvhpCQObynFfmlfoO9C+UOtQC4bq34djC
Lkltu3DN+SuLwxAynbhxKWzW7XdDjN0C0eXqoIIivP21dhWmg5NTfsehJTht
TEbs4o3HhsmtV/RJxalREV6T46TQfeZR5ZYZ1vBCi/1GWSbISNiEmQXjYofr
D6NHJf6uvUbro+JADfktph1axo2NoIR4GCEGl05M/Mh6ECzyKPmB8FShk8nR
iQRz0RrzwNVtJ7eoLUQnhUFRup2FCnngXJ4VdFzjLLdWdMPvpPokfRory4Dw
kgumUSttb6+nkhvNB30+gMBsGNVIGf2uIam1zvMl87boViRn+EctB1nFq8NQ
fZEartzs2/uZZ27VobOLmM2ad3OIK2b4+uHa5ENnmTVmE/uun+PKX9KHqUuU
D2UszfPUO+5y0hD3Hf0bPJH5m5c9yvBd2FNeuJO77D0swdFkPOct3e2/X7uX
EJMy7nloUSxK7ZcpXPrliP4k/XYv8YAoPpnlzLHYdPZGdyD6DJg/yyd60m56
0DhRmcssHoxYu60/mSy3u+gVEuZCChV1ivj3r69qwtMMBW8hj003zkWcLAU5
anXNz2XHWfoKejqzQuidxPL2jYJA16C1L0lO3OO/zYBd3duWhbiEgPAhloa2
0gxfpUnqe6Kg+n23GMwApbflrwyC+ymNYTCZwEtbfrzhqjnOjErdsuSotXx2
9S1IvkWbmG5riw5x7mrJLkbo2tMEH/h68PZMT3uPrpUK+lxnOYuhPybWrFjG
34nGnXteAiJy3RiQxanwi63hifQIXSUhLn4tgD64qFPG7IhbMWI6MrfFhP1d
ym7O3q6H4X6oKp9CAEtaT1P1bNVePkAgIBwgOIDDZrOkTAorohsMUndBKtBY
hRpogeaTn4if1zJ9P4SYoNoTYDRqk3Q4NvXwXYbfBSJZhHP3HfjDO/AZxQBz
f2c9KYefVsjFEV5YAYU0AHsgGIIrhkX3HMhTA17IBn/1JLzkT8Jua9J6Bb6+
g32i8j+LH8pOUm9pBqgOlSJCVpo2+XTvbYeuyqxzbhBoYeHaUHehsa++IzCq
YU5kNUQbm1xicoNROcEAJ1GGRhQvCJ/BVbFLLqJMd7LBowSOnz7F11GGvome
EnglO3G793E5vbPCww2g6S68mO5PMo/W/qXBLzaqVpe04A5xg/c/KURWV24O
dkKuKVHFQ334O3F6hbyTsQdvI7tRYSUzFDpD4kF114RXgkE6mdbmLbJlRjhj
TUf99UmUrc9EasaojCK0hHtjkTB9afbxMZGzKUoQfIek3lYSgHhpopKOb2vs
YbHW3qyAgV0HhqwgJfOWFQZrbkz8W/+T/0CKEuSYlB+mYyo24E39GuIkB0yi
ewctuJI6eSSMANoxFnUc3UoNz8R/H94mAfITBGZu689zEHq9z+DsuNfnWVwV
WGiYfFUkZyhfq1RiV0+vzelnuCS55bfok0QVxuXfDel26eoe78gGuvEYqm3B
gdqXNKLG1WQGLaD9spkIvAXBvfJwGCs60w0IbISFnxrxklSdlT0QbTEoVYNu
kRDMxlC0cejvSQeacTQwwlUUcuR5Sm4Dbud+rto/I4tZ3OZ1MS+niSWoglnu
al8wkRW6ooybI6O3H2dTXd3GfcZ5UyzbMEj3vR7bZTHjT3FToXSKI2UsYFjT
lLpF9cksRxpycY3OzXY0HhfCyMx0fCbgZ49J2Tq537nFgOtcd3Fxfa3d6Mem
SSnf6QTXewq+Gfq7MLbBSpvkBzux4wYoVD0I6lJk4abc8dGTq564qw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfQNwzbpvdSikAOGk0hORAwlo6c0zSF7+qx4ZdoCk6NrlfxCIS0HlJUC8Q3pup4V9wscjHoSxnxGpJAV/+oQFrcSDu7RWZOJuhkW8aA0bwhgYLrIdFPBNCobXp60ndNgJlw/cPP/+6SBLcUkBpJBS6hN3Wrd7z3vEWh8NR2G6Nfu6m3nL9XaxtBCCOMFMi3mKC/7LzMhZZI5K0RP7oIYc2x1xVHegV/0U2YBGMgrxhav9QlAsQt0Ysr/vi70NrPx8DZC+jjV1WDq9gJdi9Xeg9hrOpbXKsrPxHIf0pWbjiB1c3N+hb0ts8hWafRTWugS0UaLi3LPwbIxK65yz480pm7dE0V2FyGczMpoYlEqWNhZDri/892i5iZcheMBzLOJ3a01cFvEMp8aKIolWzojRlWDIdLuQDksCP/22/lHeqv1gCCnX8MY4b3lpaK1fA0IngSaKaNXXPsYOQIs2p5NTRXtaYxmULcPkTOgzpN/Ve7B7zZfpwYqheU2vq+EhQChdYY7w+E4ynuXBAKxsQ/jr0mYxDUnnyagiw9kCXSvfos7JDcd0SlVAXkpN66IQcszT8oENq1ScXEzTqsUQFSYWhlG95OUNysUZtpd7aD+/sWRXKO00js26Mi7UDUfnPIWWeYmvD48hmH75t2iduu/bxmhF6/fXPMLxaVsVWSL7HQZeHQELsSFz6SyDdAp3OGeBCw7yJ/jaWd2Wa4PmKkdQ/ceRdRpH1M1HEbvJUD3TSZY11IMK7Kj5XbesA5HK0ygpTisQ0GxyurF3eobIvjtNl5D"
`endif