//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Wq8hOpCvnZFu/BThw69u2W4WuFi98gDkIZtJb+WkwwZDJ8x18+3wW49WhxW8
KY8R79p6lpTtDgYczXyx3WI+u3l2Rm+5xNXA4C+Y1rBy7I47Y75epFwBtjT9
37+hXkrR4j6suacGC6XJOBpVjtV1kxn+F20d0uWfs/nLSHr9NzFGzHtI3+Ae
UMrOJZ/M6Wp6Brm8wb2fOfwF1cC4FSaWbFc/4ptt4NBGyZXpHmMalCSJYY1M
IM+zROIBPLVj+irm2f/ptxaYfzgZSlXhmA4SixWaKJoidAkWdk+J9y6ta2Ci
XtKkU7r9xsgTR/YpzLeGOg35gy5agaYHg0JihDfyvA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YAKM+coCszvWGJsU9STy5bz3mr4ZKi922Xmrx/nt/qaKG96CA6/aKW1IKfj2
xQzsACGndrm1ZAHTAwglY0g3eyoO9LsFQH6DEsxjo1Z9aVW4pgrruxehmIjW
e2E6To2hrpqRCWJoaBpinIIPMdDGae8TPGbaXbK7btuNFXlH1gqFcm46YEY1
vn+L93jVGfariiQO79GLfUTsmOni7cdnNqeDOHe/z6uX3JWRm1mLpnLh2ARm
qKFyBzIqD5l6vEN6TaZTA7GXh/7M2l8+7EShMJbh8VM4A/0/vJd5ceSvXjj1
yPr7gUcE0Zslii5lmA/g0WiAPMRAgvyeS8qhftbMTw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fdu8JNXHz+W4lwaXSUCZ831zoRMTwesG3ZWEbv1clS2XoASiEF11uOod3YhY
OF7XDH8Ap7d8Ja7JQjPXl4eKjaq53GwQNnSbtHArbR4O0kaOEcUS2qwJ89ff
LgpHiJgFnNOPFtN4XBUkKeCIZFyHT/TTUiAyCfRQ/ve1f5qfzOYl2zZ8nG5a
9R/vAGvk1XB4R8FD1aw6FahQ0gXFhBTiNIGIYpxVsncQKOi3u95nJ8e4UCua
8onNDpGdXjQV8iqCp2IXo2Wipk+PBlY0q8J7dmI1tfgpzUGdjcgJj6EF6AqQ
tdIqm+JdjlyDDnVnrZBDDjZd4usNdpUw9E1JAnllYw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bNtkUgEg9afw+juRuFqzX61ItmIyBwip6C5Wmnj1P8ZPdj05TKPR0K8TI+ep
Iv3L30CpSNPc428pYa/AVXEn3hpIMh/v86AMmZk0UupZaLP1I7azYO+sjYoU
nISBn4oQSP4orWS9WFRjLV2MLlmUXkIon5kqdvjw9/WvuJnRjyc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
DB1AVVvIOMFTrcgIKPXEmpG4cR08pfolFzmxfz93mWh/0vwZHwn4GMcHyNWc
C7+NYQIAQfoaPQh8sxsfbLeRsJd/fhZ/0uhHktfNaXGl7FJI41z8gL6Rl/IR
x2aePYWJLnA1HpS29iNkvv2oOXYuWSaeuCvNgrwVA3BTCwvGYyjmWh2dbUIE
zGhJa5UsHGwqLQI+fimbUiTeW4xTq9vlUaqlL6QHhFTjOsOXKONjR+rl6mE3
88qnzF0hj+RGLnP/UzcLPH4uddqJl+NQ3loRKh3m7XbKaWn3M3XpXrS0jLex
TC2HUgRJ9875tdJgQiyqlNcCkPyfPrHrm5ss+1RLt5w9/msmNHD8N4QMrFXW
NbnKKYxhRL6J/UL/wOArf3wfR4zaqoB4nByAMSEeH9pDVKeZpDZZaV891EEo
mvwtXLBFqciwxtEaWnmATjeJCNkxCR7HKwN1xqIvOCPTPR7sVWZaY8qcBPLT
vxuEKL7Bch18Ie+5el/JwrxB9oz+9Hwt


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uzj8iJy23DxYwBwplWm5t3VVj2a8OjejgT1NvJ4921vnfzDrYYBIMAzaDdwc
5RwPG3HaG5qznlelf5O5UsBcwOfYb2ATUcbi2zgn1XAfFVxWcJwfdPpZVku9
PUVNRVTjh/IIpAUCWu7G0oDEJ5wGn+nss2uD1D0JNdiKId58gEQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ohMlg/RNb0cHqr6oLIHint1ggHYcW0dFFGJD/0cj6qWPticoJKYtmZc0fbnv
51y+POPX/gxDrhW3l3xVtnyv5+5CJUzIosTh1ZPbRcNF7OlESfWOMVTPtrtm
Si3rYlgYexxBItWb9PPf5t8N2fFy+V9Q/9m7oD69JrcInPkRhus=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8560)
`pragma protect data_block
Df2FFBnITfSSrEONIY1IppsGEr3XokC0J36vkqBJx7AUqa/yEJ+zkGgSHi1q
SJRNzgSjV1RufUiNozgj+FFS4ZVgmVpZLMqWoR7ImxKMnCjMRnO9YaZ7FQo3
1u7gxQ1h/C+QNbUx6nkJbgp0/l5A6xrrK4QiMkMnXOa8zqIgNHVKrpX9yymw
UKpgPc+bJad0uSVVzFC6oh+6hP8qh+mV3PMjnmNkye6520b4lGGDPnPzlJCk
7vswnib0rZd2jnlZhWF+dZm8WXv6vfBH/kbbcudbosFgkg0xJCpnkNBbzv9E
26PuuF1cvPpwPNgHTuNfgxSGL2s4UfrOAWfGoy5UNZRQblDBbDgRyfsY2fV0
n7kKW1iOiJCr1DHTvC9RenoaQxIAbTTpx78x4XFK6TwO23xLUy8fIj4hRYGD
LSZLF+/lW36iqWq9wacFl6+NKsLdpiEL+L1dPzQNK0zsQmwJsoxJzfRmZCk+
kfvhOb7UGdeYtvvSJKf3H6M16bQtAwldPdKyFSwr60rRWX8VSvoa3z1eDxNx
Hjx8H95huxkWbhSW1eogkKK+GAO9sKCUXh/ZK6IJpa94oPqKJbYs1YdrmrYM
HgVP6S/yhPoWPh0icCj9xzVkOYXqQ1rT3ifb34BZEHo0y4nRkopzDHGz8/py
sarA6KTTyMluUScMRq9Pfeo/kPOYKLXf6ED4WCXDoi8RAb2PFNQB/ykr16Bp
PHMOppWGWs1DVnkH2uvAjU2mAb5Iz1GOPIceSOT75Eaihim2ov1FCakJtizs
dZHE6uSu8xosOCiwqLtUJcFNUgcPHB6NyT+bGhXinr3/09UEUfWFrnaJn+a+
GZtpDZdgSFnVkjH/Eu9tqwZbZHhE8iPzHS4Wr+WiYVjoOd6WTX8pCqx88CaN
R142kJ0r3uUK1z3LsJdGLtv3JStiiN7vDbuHjsokPVfV9I9uTFz7AosYURI6
fCpwyQtYPmMynLXBCKEbQCTBjrobodkYFN4HZGvf8DncD8PEp9vw8E+b+K3k
aVR3Q4JxGyRQDXWmhkxi+WFAAFDcnme1ABT/D7BQryV2D1bQzPPK9iOy7kXL
xemSxJXD+18ePapWzmHUUbdfkqJ8xFJOsNzwQKzsHJFxJGQSKMEbPLh1GSg9
V7xFRiVErBjl2s43seo3FG89T9qSJXy+Lg0fGvENMLc58KKWq62TVHpYVbMK
JJBTZoc4ytNvr7Rh17pcKwgEU068ghECQiP2Zid1kpeyA6T1NqtgFv3umWPk
JlHxHglOj6cE7WqNQ/VYbco5JYCq/c3lvHJG9dtzqcoVNjbqgPUrKMC0WErw
gNhs+QhHpihgg+xMxGyDIbGQctVMtLbJWqTpc0nkBb4T6Rp5/s5AWw9PzdL8
oQ/xNyeHfDXiVEEFgFz5Vnu0eMbfl9VXpdgNRK3gUzR2Ic4sUxc6wHSuDgJ1
bA+hMHNsUlX9Utk84HwSnU080B1gjI35Y3fpt4cBH91sCr+NJ2/aQ3jzkXYx
tVPR72lYzOoxkMO6Xnv0mbbTV4sdDszt21a+NuHMoFe8mKWIjV5FrV2QLgOu
mIYu8MOZZd97bnkuB4Wdgz3N0NGiwKOg27bpsTUIp9Sk2JBxCTx/ti9Mz8Gr
kXAzB7gxca+lu3g1Jg5e4xh49rttACUnPDYyVCoxvV21xK2UBUnSajcuEFKt
GvsMBSwF45Jtn/U5j2LJ/R2lxjj9xPkCTtVPVjk4S5gukcs3JwrHMoq0VVio
BihRuC/dn2TxKKC9uXPys5Yzickw5ZXxSRspccP5k+c6ySmwfajG5YjoFYzs
M0KbEQ8LSfj3csMC0aiIzSW/Lx01XQmLgbUaQOhebR83X+e3sO5DvM+HC0ag
V3P2tj7SlLgUAPdVUIQtLC67ZFhsx9xwNldyPcSDGxAwy26OcM0Zq5zTPsor
BI1V2VcBMwa8z3bw0am5Lu6CEAbJn5NuWURKuQ1eunEIMNUkTDVsMshr+IRm
mMf6NyIbacVdK/NBf8uSt/adi3mXcdWhNvrjGAwBFIqZsBDW3ig/Z4T8wVqv
JJoJ0/igEsTUeI+NoXavCrE2peCRhYjM2icX3ccyhLHnr+qlbD5WgQybeMP8
iDmqQXRzn+dtG5jidoKhc74lVHk33jHQZ3JklBtczNqZm7yOTTmx1RRvjc7t
y5wmBri2l3phb2ORMC9/hu8qi208nvIkzrSAX5RuTe+QntbzpKzsKTxFGDcv
xXQdvpxJ0kFIwIhFkO9vfa9BnJVYxIx6r+SPz/TKLUf0cw1JvumhzGrsjiNQ
X87Ruv38fM3Wp6mE34RqGNyYxycNbcKwk5zH6BHES6zfe1vms4hUQimwiyhS
WXhl8j35cAB7TAyjg20WqwWQpRytWVp/WAuBekuhaGsqLhaCm5CVueXAMSlq
SIgZ0qlwKPyqx+LFPbnSC9u7jJ+z0gopqFXTq0xmOEsu+97wpr+hTGLqprop
y4IQKr3lQgSTIAtQKqCm71MNSFj7eHbREC7dTQm/wKg3OKmoGoZ/wU7iPAMm
4NP0OfMaNj3nKFLEPbRzN+ePZDJV7rC9vswy5h2P3Uj3sTBEXnYpiODPBYqv
A4lQnyPn6fDde/4Z+NABrMLGRfL5wFDuFO0lQxyhYM76Dfjwk93S4yCYxUZR
kUkq77tbBrmz/co7BJ5eGp/+HL3YOryWUhtcx057J8FkZANkrhNL1n6ZCM2D
PyY4eQbml1MmPQ6Wja4q69NMtqkXGUtrIcOzQHZzG8g0w6AulFcgnPKZSeOl
HfN0sgCIojruc5R0J/sZOpPKss+OChTGk9eNXa6+VilMiPC849PCWQ1LX1Gv
C7z6ixniPfwgYPRUd/QX/1JdHi+Oykas/NYgSDFDQ4oG6t4mFV8Rgela0pW3
pV/Ok/JpISZ9tV8AYTv+kUOUI3s6GyxSmy3pH8cZ4ySSoOHgMq83KD+qXF+g
x7v05tnkzNAHNyWIhCTe1lsm8rBoQ01exZmCYYIqRkOlzVB/qPfOvjVAcT3L
9aypuudZWSAXRoAx3G21OEuJVfC/vkdQdWxq2HVZgs/1H59cD44JPgAg2ITl
LkNbBXJPTNqddHl2CCnuficlYm4SiwjLsIdSETH32WJnTLbuEJGVug9YrI2j
lGcyvcEoXev8BXTuLBonkqkImCURsi3rWsFq2QD5xTmvcFBW1Cwsef1oozvp
Mzt4b9wQgX3+zYPHUKhRfPUOiFHLEQYJAHrMCVflknu9t6Iu+B+bKN0iich/
pEBAGrbnBFuAOAhCn+G9xstePZkObXbD/c8Ta9e9hJxbkV6ge87tf8bhFnmt
YfEd0zFV/NkRYkDkjGindDshTHpHSMgcueRw/RqkBqnJ1qR//tWuOCOSHtOc
BE7/RWzyd7vH7VC3DoK6X9g44SkQOzSLxOzqnTRZv5gPwWu7yxjmFWk5wkHa
mlFIEu5cdff7p9p8I2+i99Q6R2HvEutuiWpQ7KwZJRMfp6EQ4K9z2NlNkXNL
XtyIZ32KCVuofpbuP+d7NHRunPNt7P7/1S5AgtAG1szZiiQkPa8iEPaf+YeK
UH0JAwXo4+EEirO9DAXCb7y3pcFlWrUDyyW8JgIhGrLwrhVQUMM8OHwZUpCX
e/kTTHWVrq9RSpstzuuu7bJY/gQ/xPezKavzA9E/qZ13/YZmCe+7TOBt8yPi
ljEE262b6X2tYVViuaQIrBz0HAoWfCGSzNZ1WAnzJjCLw8/9wIGvij7oebHi
s56tQDXXpIr6s8k9AUG5j0gfx+w0tYv4jReNKkeJQixkbSGVLgJheoNiZ20w
vjD2JWESWg9HwWZ2mmGVUIrMNkjm02wP+Wf9CK7BuiQQJlw/H1FXCtRyBHZO
FuGaa/X3pHolcqVGnoM8EBLLEjSMq2w9jzf1iIcVDp6GWmTwhpoicYRmKc3T
eKsPhScE+dIoNVAYRGbjvOJl/7mo6RY0BQW2AUW8fLhJTNWdOjVMh+UZ5UNG
H3s276OXOf0sVQMcMBWsol0OERG4bVqpyA5jntOe+b287sQJULcfRzcfwfhr
0e9fbduTSeJoF6gB54Mu5urD2/2+A0nyGvFXN1DZVKjNjAyA5bBA8nayHmUL
vBuJ2gRqIbKxEieqbJoSvusVRrGmTkQvjWCutHcQ1oZYl3FyrQtRFO00qwmM
hjpc5j7KJUYtNvEMJnf1fAgoGB2TyGmDAqolNdll8iI3tDE9tlZKplspKlSz
MjzgZBTkW64BhE7HgOn4X5U08L/7ZurpFTKTYJ/VN3gkzxTgybGONlDoVVub
urWdWgE/AakQAVSDQ4TGtDVL1OLVio83mrO89fOEXvzsdHwIBgktIGnPSORs
1k1bg6IzBEs13NDQJQ0Ps3+9VNN9GebVQVF3Gk8v8pm2mnUGV+GRfx15Jyk0
PbnLiq4JrsPwo3o0E/Z6WhgMpXd0A8Axcfln69CdrzIB8WACBw1SxLzwwfQ3
ioqotiOaBoPfzhfHNGRH+BnWMjqLcdc0uxgmy44jOnX4cxqnnJrKmSetCp8A
eoa9RJA+9sz8N+8j4hrkkImwR222sXeWtR09SIqzWthsjOGvafsLATk0LEMz
OmKb2PgrFJ9uAPLKbd48cu4bvyujfsUV7Vz9ZC9W6nuYRhyprrraXLyXDcEf
k61PVa+S2faPtKb1SJ9F3UpqmbJfhNyjqLEC+rYI1+FiWIb8E2kgc7iB1O40
0oEQZwJvU9/FM1FYnnj81BjH9tA4luKp2r3nSWGW2jLrDCCk1s2cPe8Je2o/
UC8Y7IdfjvsT6gmvtTrPOt1E0Wf0JzrYALfU1zMb+VrrLZuGywjNlbrUvuQT
2CEc8Vyc+YhiwsNB5LqyeJ7BV9op0+dH5IA3zIBcNeK1kW1BQ2/xm/li4vER
ac6xLS/tFN/XS52DqFOGOPcx4XYAtvgAds+/FVFilYUbFN9V0mSVhpTcM8u7
ps34lLCOZE2gGUW049SzPiZdQ5bSLtMShWcnvzpkGLaRUMCxkIApurDMpfUy
FYrMaz1f2QJLyQDUd4GxmTYnjyt3UWLLNbXoNX9Ftc0Pywb2h9W7DDvoqb7F
ypmx4ZTQZXdYW0suFjh+8Vt4+I7VYXVEWjDGF8ZS6Sle/yUaqJ6LoNQwsuGo
U10slxYUp7JSVdV/H7vo37wxJXem53ZotCtlbO/H6r7C+RIRj8ZPS3ILMVjp
VGIEqmfMLKWPSKSHjkrNiClBw7cax8FnTutNTtyX9YZhkY76h7mS3caDlht2
3VWgfsdup6G+bSx8pBs3DDn4G2hm/sd3TGv1+AqASR4SfYRDzwYKGU/zBgT4
E+Lcpdh1655QY/bpskUJJBJ5D9yOISANFbDdMsbEiVopj7u+cn0wzDSFuwCk
QwFPcXOOKL9r84cGYQep7VJgs++4oSFEH/HPBFCd9Y5IiIfAhWasFmldtqYz
cJQbZjCneqdTWvNWUBl+na4WwHKHNr1dAzhaVoj9buJOJHZIDHgvRRFBWLnt
Xs6EsuJrL33CEH8uoXQdklmSI14Gdo8KQQqg67g01cMYg9OfNEL43DlLf9l2
r4D0IvmFlMVXy9YKGVNbcDzsGo8LuuHzFuN1yhQnZb0zIFuik/Lfa76tYtzc
Zz/Uremk1vs4WApYwtn3KL0GFSHdVRcazTU2NMtq5ipNobovBV3UgDRB+fbS
pmJL7NpcqvN5fTQUwGakEi/faPRUbwygoPX5ttenKhk4S5QArnC8rWNebJ+m
9kqSgsjBwri+JW7b6f0RZQbXSKaEyTX4w8aAif+rzSR+vZd5K9ZhF1XBZbFH
Ac0HygTT1+Ojkas07NV+ELUmZp8o5H9DmQKdLSmuWhXHgIO8UBQe0Q5JRuvs
H7CWdVrpV8x0NLX9AFOq5VcX32D8lcQ/U27Jdcr7HCqau2elNWKKuyWSoOIe
CzjUhyMzPYVu2FeZnkhRWYRf2UBtu9mQpPPQqAetiEvovwtNntHQnRs+KpbW
MARRUo3WhPcHZoaMKWYPQsZHqC11+68EYmxusWGtnK0p0HUgAWsYhepes95x
40AaNiQ1SzqDDupmRYSLsNVlZEZuc4v/84lgFVawTeHOQ53OYt7oK8Fx6kak
nfP2CBQAPbi6YHdpvqopj/JJpdApPR3Z+wEonNuQM33QHAodRswit6geIK6d
c5ha9uDLlS7VKkia6gsNHBaVMW3FXoS/9wr1M2pyPLXKozoN8XdPyNoB0Vsn
6vb5qAqrJUaW21oofUIYzcHtrWwpuLhNmedmALXfJRdfCSfvkP68WAvY75Fg
sMcR8C5pXiazjxSumd1wOmdkr7/dwP0MUx9VznRPuryi84CwxD//dfGR13ay
c3Ev/HgXfFJxdsYvU7DX/cQkdEnLY9dyRsZPlRnQCvVqaD8jKlCvBx3QGTMA
54TBniJ7irOIchniB0Q7GVCnV8+weBLROLd0EnaShLLXOSz6dwuPpYp1njKI
0w50QMzcOsNHEw0oKaa3imbvKkQrS3NiUEhBPL/TH3EFZ7FRLdTq1g608kNk
YcPea7EfRN1065ESXpPK3SDflnfRTid0QQd8z67b16trU983SYk5E05GdLPb
LKEmMZ6TovXves5lExcVDTww7J3W9i6IYiX5iIWZu37i7Rf+3IPzWyzFwqdo
UoA1VDjJFWXI6GSl98X8qw475l+I8dUUP60ZIEkJ1x3yRuKywhUPbW1IKfeT
AErNWYb6LlMnqt8ki1E3/51Z9VCm8g1IWPB2yWeftBqdNB/cF8QeD01geIZd
YnkT4zC521nqN3ZTkUK/6QbLVOHgDzdOj0S47hJostbZCKTCbfO/ix3nGqeT
SUC3OxdG/AGuMbMX11r2qN4/Fz34x5rRow2oXRvaVltIIhHrNSx8CjpUw1TN
uL0MVPY3BANN14TXMSBfeZodQFUQ84FWBXll3NS48M6zxUGbfOOW1D0ZCIZd
db2d4EARpAw2IbkBhFDfahg9TksphO22rb0FdayBt115Ygg8ICJZZXNYOm99
Owne7xXylBMjBh+eb33SaTSfFGCIvdYXA4feoMk6kYCGs76wXXX8V6JbJx1v
U3/+70tDJ1oTBFFEAz5Snc2VUNyV0QYtVIL2I8sfZ8nujbbpu1fihHg3YLT3
LFxyPtQLnI8SOjT39PITjyqkYR0Jptx7QW1jsJK+cPezPWq3P++Ko6HrjV3Y
Rev7FI7Ho93iAZmL8Jw/r6kt5fbXI6JsLAzNR/fYGhLqeJsJBx5It58EWpRh
VEzYBs5EUGmXR5/f0fsdUyxTSn5oikQyM5EDwxwjAXf3misHZFPOrVc9RLc2
hC3d++76yt+eirqwoQTYVa+NqWqIkZuIo6VO/oxRkcjohWP0hdaev1wllkcQ
avC8JtKW+youmpwEvt4tjCElA13jCJEIr2slBsmELLvIzKkjPiny1u+gKX0g
4UrTzWDPSpEfmgg2l9i+NjR2UwarBmIq8BpGUzgP+JAnUczS3I6S+ODPtiLT
w4HO3BGJGGTMfgRoFHLBT/FRdFQdQeYErf1CkuHzxt+ZBkUfk8wksg7XUwXM
SWIgU6k2CXJjn7aWKrG0QVpA2FC2DHooOYXfMzcAEm9BD4Jk3Zod7tTRormh
mT5Pi5BeU3HCjB6dDMGOBZi22CIr/fj8pLdqvGLp99O1Bg2Z04dxC0wmJ6T9
akegg6eAu5ZEatgT0kOu10Xuk5PJ0XgH5dD+AdJ/mF+11JA35Xu5eZcIe9uK
ohsT7hD2GQfznth0KuX+HRyuzFscj+jOAwnG+0vZt72dAvkfOlzP8oIj7+fn
S2qD7NveLW4KlnlW0sDib8+BKaiI1P1BcxAThbM2pRANc+AcOp3JJFluAra1
dOwQx4tzEUHocfKkX0zkhsoorHVEk1jagt0VxF8ilTzfte1whLOerP4miyn7
E57C4f0YB06wuV981QPsKb6ud05a4M06kF/xyLdB5sEjv4YyxEIvgEMgKjEb
5kHmMpqRCoqUh3Jn7BYd6GLBHXwrL/nV+kRWhCoikA/nybReWubPrUfkd41D
ovwFnkqh3TkXQLarC9umutz/5cEQFwdgzbRDgFbMVX2xRI/o0FME+ScJYo2q
TKQ8zXoBZwuUZ/XLvqjb+R5DFUu2JCaCs41cLNWhAna74UDgECnQV/aKUYNL
LhyvnJiuMy+WcdP/s5DFLoDrJx2y30f3jXe4Wd8XQQWxQ4mONXgf058AdO9j
4roufNqHweNx/y6IRQr/fup0wPtgQK4pXv3trQnHtIyBFMSuuAINkjar8qvi
b/wkfey/msB1/loQACS424RdOC1KXdl33znQoR196kv5b8pZcYwgThX/4/nW
MFgfoc7pR2cIZbqFkx7WiuCqNOn9Zvx+O8SQISMzypRsfGfdhaEXwulQl72G
dlGcGX/YDzPgnEVXiAmu4Hm+h9wNfVQMhWFqAFiy5dzClKm6RXWub2q63VlQ
NcF3p1rmlCl93awh1fLOeKov8d4opC7DgJZUxqMxOj1RwF0ECw+evRj6Ql4I
qvZu6eaVM6FfB+Y1zKju2eFF7XWCsQfASul6S86JNA2bSYdcdItUh3nKjNK6
DJVDOQPWjijWacV1RI2ZsEvEZbrXEAfaVvuwSnfyUAyBqXynGyO0+65dV+N0
h+sy9i+nceFdv7EFD8C8L5di6oiv81lp3pr8KxOd9/Fj6wcYbFFfCP+VNVUD
UcjpwooyqoIZtPUnMrWx+u5EogbPSU90EUptXIlQ2Mu+1vdaiIGXM8cYuKkW
4OwW+EdCtrYQ0fsI+Iu2RBJ+jq7ZqAmfPNu7Nuo5zHKJVqM0nIglCu0Jw5sU
F33UmVbcyHqQjDaK8GNGhc/Dgvq7JcTAW8QQr3IwQNe2kolWXIQJ4yT3pjHH
11EAoHdZhHyjyphemCFSDjSo3EncW4irqsH5WNY1XviMkOPUm4/VvNtcSJ+x
BX7kd2Z5kANp0q+oNfJ7lDW7tFN2oc+YqCtUSkmLWsOT33jfC8UwC3vy+Zl9
cOXyXjQKUk/YPWjuN8E6dDsAIUnMCRNLbTPTNbhyUAN5XTZI6GIiGMJtz8Sm
seudf+jeBzjyk3I4G4BjLhZCIFgis205zelOvDDjJu1z2a3I0Qwna05r/JFF
+qbYu2LkrhezqnyO+L+E5Y0FLkYhh4jJVSFr9m4d/xY+u+aWUee6cknUX8DG
0Bdj80kre7xKeYWUmrhg6qdJ21sPN1BLofhgAsRNafl1GIbQ0WhiDkUilwkQ
nsmZM59QMEeR4OyXpSItfTw9t04v3LEDVo4gL0pcrjz7wfWvRpkuJLT9Gp1i
U6cMNR2+Uocg6BpzpgGQMPjJR9CzcfJG9/LzD9IpUoUWCjiRcXBUBoJC03Sc
XF0USYTwFjUfNxqRhuX2nF1c/TYfQcdKQ+kQdPdjB1P+ENFeZIalhMp3oZ7V
kWyeoLLJzfUpLzKTXkV7ypL6IMKnaPGPElxLpZiPpYsepgnmCFVd2lq7A+iY
2wPr0o4BzTP0JHFvEND6zv9xJjUZ2Juob8llbrezcVxL1MPmeQtvhwt9hAeQ
geeo5OH7MTXR0a9glE/F6lCTufrp6WCcSS8o64BoFLOiqhHSZ/HNRifJZoID
6f1Ds/aw08kpCaDxPqTt7P1y7i6rQBXjmTVODNxJjdTZ+kIcwe6fHdKQe3FC
czli4hMOZWsaR9VD8cWoEvqwp4424O8vWwNlnv04c6xHNx3zbjW9jXn+qJUH
JtcH3CGlRE2aTSc/JRuJdL3vr2p1d7u/7nnAPC9HK3D5z1C7tj2wqNxOXWB2
RvA/H13rSe0enBKqk0N9B1urV8RGInGn1QETnDwnMI6VjZPqgerAdEpsV6d6
2lyu6kSVaKgKNs/yOMJ0PCUn1NRJlaWCL6OVX4aFMS562To8PcB6WzBs9Irh
y+tu6JBkKMxzaGp88Exys45eXKW4U+VhFgXMUIMm3FLikj6D3ef95+69ZiG4
SOkMufeTD7lrw17ma+zIcOcqgWlavZZP1UPZJVbUDOu52G+Dn5X2XStwWVFk
GbANHc2byAlrmcBvp54F+wWn28OyaeYy26VgJHB7HKZRosOEsa+rTeAg58/Z
kpF6CVO4H3ICd1IVmX6dVQlfmAZsH8Ar2YY6+DL8wnv/LPQBNJI0RwdTmFCW
uM21G/ApE2NMwnmjGAsM0J3q6nlsuQgP8YEei5j9dvAjLSW7EszmwYSRi6b7
z9dMaUpilfTmtOIyuXiWvilfnOFPZ8gHJqyCYZmBjkqnFbtHi0o2bvo1lJA6
KcbjErHBG//DLZtlV02JebV4DQiIhuK6mhWoY+yHLQsko+YhvX0DXOGkHJ3h
NdcU2UrjK8G4GcWyXcrtUCNzq71gX0unFD5weUTbUSpbtehX9aNf4i9Yod/d
0OtsbR6ypXm1LREIp6TAlTf9I8SErZm0K7j8gMe0PbVnoguZgXHYp9kSiI1U
LjXBS9mae4jPhpizP2BDF2LzVMcMFOil4CbQilxcDdtFoELC0jxCdk7rTch5
SK583WppFx2+Bn+x5Y6SFOGsNQWkqnubdxrxgm3h/bDw21WpcXaW36X1tywS
b1euk4Av8Q2hFSyiuw4FbL33036m9yWqM4tkKIGB05wETvL3+QS+hPXoMFQ4
EE4i5pPQ0I4ZfP3ws0E33jRiorLtT18czJwrdq6NCaANr1SMJjNSOCbcXReW
spcI3NISRU14g14otTjokt6XUkD+Yx6PO3Tgu+27OnZ9GUZ55pMXACS+tgf4
CxJHTCXdzKpPInbow54VHSd3JybFAn250nvCu/IUz7hwf/Fmf4NzI4/OJejI
fjA0z4WbZdObdU8E+g6XUd3qtueYjGwVKslSxdsPtVYxzuBlw/BSTOpuz4sv
hY/3GYv+M6Maeek9m8cNNDpMYeE//n37loihGZl0t07Dric9R9MSkaU+P0PF
9MbIjlilifyxD8IrovljcaF7zwjGwafyrElAEk47AJLUZZXLkau+PO/WVhZh
+UztN0n2cGEvH9k+5WsWlYCKOgjdlrXkxB4E9vwdhbBRauofkzTl+21IokL0
WkelJTo/fhjtQ2m8jC29t6JkJOCq8mRMd0w90ZpoaMZXwmAnHkK35+9YuAYw
LffOQM2S9miA4UmJtfECTnOtifwWrwomRoiYEpsvbVWmnC5nsLmqxt0dw7Xx
txxvmqgjJ2p4NGmOH61t/Xy6ptkrOdwnkV3xtPyBB0i4QPlbR03+qtZJCqv8
ABf0ZWAZniMCmVcY+6fC6b3OG1wL/XAnfAOzEK7WkyDh70a+ufMBLzU/fpN3
Ww0frwhxj6cE+BlczAynupMkBsXPhDm00q94NEbVH/GhFlJAHC4d4I/LtS98
BSaziinqB/4umqexTqYI3bCaTcFRm9cjwDdHblsjv3sdvCYWrbxjnWzRI0ii
/HidiKSNKn9Q6A0PIURT7asDt8urJxKJkRN4ehFftVQTafU9dZcodpa0CoqW
Xlj7yYGpYoGWuw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG0fjUXmCsckbCIhX4taIDktQDgVA1We9TKwLi/HJO8h8oJB7uPFd61yW6DXXG9wjrzkLv2Q4aS5n68xcFvTqqPuAus6mJ+vE0tlx3aFX0gWz2KZd1WzRuovhjUqClyG+CmBhiMba/qtaYOMq1ZQZ7NLWVIBxBoY6P0ojnXVrkGqdoJ26VtvkyyjCwPFi7DookA/P9ZKVvK+dwlhrk6OGsTcvZYP8hPFHd5U6J3RHbaMRSsV87QyCxM/f4tVx4pMr6qQyOBLiXH0KYadQaLgEwKAz8v3RTDSUTrgHoNTUa8mk+PT7/AKagDA3Zk8wg4cQ2i/hcMSt5k73A5suuZ5sZYB0IAb1E6cdWosRHquWSmbamWfJ3z/DmoSDd9/nNvCm7ZaIFc6FBgO4VVQiHZuB+bRiBGO7hu8PYm0xtf3ZcNMO4SLsq1Ldhf122geot9LTsj8GSo7CJFmmVdwEf1siHJkxZrkjier26r5Fsm6shLdtCSjhpXwuN83HfDDxAfWR8xf9v/qgouAq5M8aZvIhXkpVoMqLwC4/TUDPnBIguSCUXfBF9ZObpjJ0XvrqO5Xl8nO2yxCTLUbc9+UMfA86j3dukt6gi5rah+3qXIbGTL7xJYORcD0iAav4LTklcDgXsDEdSDultaxk8GNpZyOCDr4ZGHhSw0yDBuQcdj/hkF+2e0rqJQ90auQhJpbHs9fF11ze3q6IJjlikjfJkLheuKsnhyiPCOgeT1UnvAqFP3qWUqAvq2yltdotokFaCByrNCI7TgUAFTxrYnmJO1qKCBW"
`endif