//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
G7tM+ffoPi4hHiKVKs3raQIUboAdsUeUqlP75xx3itTD+JPN6Z/zfBUCGTtB
Nv6tcZpVUQrV/s8f8QdUJGHYklaBcG/cZRrH2w2uJTkPE55mQcHnyIoLwZpD
2BUzWpY52/AG3U+cASuRHj9tR1mUbskvqfEpXQ72g2HMBMYjJ554Ju5c6qvr
ncafAEoMnQgFASPmdm64g26pXIUFBAPX9hlwvXQk+LjxcCSB+5DGid/WtgcO
ygXQL8uP61HCsr9Ik1l8HCDtDsJxOEUZXQgKlFqF2B5DAyVuDkibsrmFbsq+
bmKNDheMicNF2DCFtPg87rzW+4uc7tphDe136Chl7A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
eYTLy5hUQN8W0jVaKNJM5oUafF5leHLN4SETPxUrwBJuKcArzEBXp1dCvvlD
B+Eo0PwHoXFrMkJ+FREhWqRUReqsjspONFRbhxo+686oaakYW4RC8V5PRZ2d
vOVQERQZGqxv+Oh668W4VQBOBHAXNrDcNIopgAKN5GFfclGo+6j0Qthl2b9S
YetlXAeT1LxA6/TA39dlBMdumzrKoDt/RXcyHNTg55tYiD8XJMT9qWrhyM6j
M65dr1a7UEDnJdEMSCCxnVnFByyxFOec8EykDBqX+hfHiynpBzdsCYJTgP/F
R9pCHzvkjU42bxPFhmeUGXZZkMGjmqVV1V8hm6qy0g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Sx3ZwFElzbWbDNIjF1cK7uLtmR5RrPPwBvQWNUhbS319tVMJjVD6b0kpCpq1
m08xhrWzQWcIOZvhqgMKiou5yOegmbVRs6FnTYIXS8eGOasVwqt4trkFd3EW
cXrIbPJZypERC3sdxAwebP+9uncPDx7soaXPKuc+Irph+1FMFaupxk8U5W8l
qJCoM/A1gL6ER1qOHirpzyYa6aPhP4/j0p7Fw8t6lcm8q09mNQsZ6g8qk+Xy
Ruc1F5KcnNSRgM00TOBveo7k7Huf6EMh50s0ZjzdXqptygLF4UPjfJyGrePD
011s4RzJqlNiVxjMiNbc2f48mA2oZY9tPl2JETqk3Q==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Zt1Orv5pnyOxW0XueKyFsm40jFKd/IhbVOc4z9uaewAT23L0oJlVfgAhDP1O
v0DvNCISYe1KyQy+l2Xnspt08sijRO9ePVvQYCwN2DPhkHsY1dQwt8ez2zA7
jjmQBGXu0eFmGuRxlXwEf+u0Ta5CpxswX+Hsd9juMR81B0jmYgQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
XkXBn5vCxbJnNVZX1RnnuvEtvGaDz39LYImG5S19h52wqNN54Z0QbFvAxzrX
ZYiFRmsqVEp1Jsnql754GagsTcHRAPcUCFpW5W8gSK25Knky3P/BencL6re7
oUYrJYo1OM4WfUvLt5LUp6NtOQZgi2rEh9JX8KtnrIne5K7+/j/n4/ENg4X6
9PmIVEiDAjh9SiB70B9TY7xVfTkVL4qQ9IEQhiq4sU9n+wkh6UIbODrSkfJo
OoVG2OlWTQEoMBt78KRaCvjgtBiBvOKZdYk8d4g95N51yAf4ydif8tT7xQIT
Bh3P4FdlZcda/xZZ+d8HQDU1o4TxfBGF19HMvdwlBTlP6wq29onYJ8f45lDP
KJtmp0OjbO57f3BuKFQQEcFjxueiCnDvuEUZB4pWr6TT5hwNz/u273b+OgQJ
0TAxFxheI6AiipKjoGZITtsG7uXvhLd6bLd5abCnuA0VO4sMzMKNuq5G1YyR
etaEu2FzIdIkw6Pn0xZcE67iWIeLRhdw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XW/4c57hDPGLFxIw2o+/8Y3hnEyz+fXvMq9+pddsDtGjoYfjzmnwRxtzoIK8
qsWd2F0qej0d/gAqZS/MWBUK+o3GlR6CQF50W5RsFCnY00wvgVcRzb71eb1e
GGUWbFZxja/G3ed1o1VuGeMt/nP97cYXbnDyBgM3uNtzc5ZVLNE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
kFXIEMJv/NDmheV0cFYzk3GQkwsn5FOOHM6pUwvZ90/ndA1PgEEALxkKZNvw
qIBgyHHXCfwewpv/rkVxIrxFBuqiSI3PjHJYTuWwIjUP1zYQaG2/SBPvmzJU
j79H7ah9sJj9/jeiYZ30AXj0TOcC5SMm492ZmrFddtbxzP3RuCY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6544)
`pragma protect data_block
i61EIxNvJ7cb8zx3h+amnEXfFIOy2D3EVH7pd67js1ovpt3ErUDHPf3f4QN6
3QUdT5YbPM8qxiiwFI8F9AYe8w+48NVdYjxVDPugRKxYmHsd2t+IyTPDwMnx
grj6We6q4Inymez1VVdb5ugqna5HQBIVLYAoQ90A4c/gAZQS7lw6jLXrEgaj
zcLn7rtYyVoDyR+OERjQlF56ocJJScKCfyfp/nEGIgWrPiwZOkIdgGYoUpIM
EvoGDiL794RNIS2ePOWAgZvwrBp9HBE+SMeqatiugTcuye42erw29S7d3166
wioL7HdUCAi0z0lPH4jNbxhm9FafZ4VUSG3epDmTp3P2X6ZXg+5ZmirZCdZB
jA5q3b0m1bsc1h9Nib7WiChw0+YiBL2NZNvbGOMWdmw81xZP9MrpaHDTpdqv
4/cHdN5PeAlB8KRF5R/W+1biyykInu6Dmu8RCvt0ILIO3/OwCT+niPliBfOW
stQLvgIZT2HOVmO+devrWeJhyGmomo1ET4LxoF5q0/NeTgc2gUOXRSgRNSQg
U4Dyt8wD4lekla4/5SNlWnwWpHFlCAWpA6uMxyIaqE7WV2k0Sj+JraL2K8mH
bqNAh7/dHMto/9t4+8meHuvYJda2b+c2vMgRV7PhkP79ELO2BLYfR2t19NXI
EKvm/32IWH2pJQd1lF5v19vlyuckJPFwd3qkijiL7JX8/Zxjl0yJ9WrZnPc0
/uv04V9ohpBuZaEDZYKYRnQ/Six8aaNzH0GT1Uw79obmLb1vyzZ0wK1bK4JW
Kpgwa05ql44IBg2w8t/gU4/w30Dq5cqBjpmooGRulv0qa8KBtTAq8WcJY72Y
YpVTO5DJxe4cmDaH4Ye5jgxbmb6j9PlAhg6asBQJZRls8yai34oRL9tQkly7
PbJz46+LqBVCEgxDCoAfiu6ETTYFKAldj7JjDMxoInXpdnfSuzFl9KhiQbOw
ILM8JYbbX8U7R3wOzDqCJhRGj2Vl75RC+8QwavOC6UbmfkG3wyFUXEx66RJ4
t48U1CoB+RADaXClq0pUvQ39TPnE4JA+ibuyOuiBCOgxsWFiqhAIa6NPjsuY
qyGuf7yykUASZjICSq4rgvWiXKjfYnL7Pj9X8d1RQ7Bh3lkKoCup9tbEVP2E
MDM5d9wJUE8IIw2445AoCpT/sQ3yQ7gEOmJGv7sB9ybLPKXoXyIJwFUGC1nX
dqZ4N+skfdLsxPk8HSqtZH4gQY9Sq2+7JUyrio8xDi16CSSNHgMtuBLotE50
c3RChi21McriQnBc2LlNGrTvTEKXtHL9P0sTXiDewfzZ3qZQhn/XZOxClIhA
WnYd54g7xMsUG9RCq5aKdLwZzo+8/JtnwZrpEo2BqOrxZOzpX95hXfVsaIuf
04NNDwyWKLH96k9uAcg1anaSkTTbEvgN12LuhVPJhwpvgPM59+M9JQE+nZ7o
ecFSCY97NFpJPR/48XEIA19c5rBGxDkQliIE/Whh8pMJUWjf7J2ujyd9SroD
tQe1fVAk3N1wUxGBVivcxhwcSGWZk+dQ5MfTf/Lqj7Sr8VdxAncvzUDPTI7b
Erf5EOtuDGcGdMzTXOdrllDd7clh+BxqG3fO6LTidOStIi+KTqhty2lyz5VP
tJQHqq/mkFNHuxfXFKRFb3OEvuKjvfThMDwGu2gKWFpJPDWPrDpSBiKraCtZ
CotES27MO3ExWrK/L2nJ79QBCdmgZd2Nb38UABT9lXVZDKi+OiNAlMtkgEKF
OGoGOas23x4R04CwwzCuO+idBPZNpUkGm9u0xKmoqkdPr/wuw6svXvNYoFcY
f53/L4mR/Mt6NCSyyVCQWaQdCp0c/MB1kWFnlFOMcEfqhgcf0Oma65NfweNj
5SQhgd1BUI7JDTTd0P/GsDTigzgd/93bkiUZftG05qRcKg1LAbVKiVFD3sqV
1fHV/9OTyhUR83TTXKS3DmyKDLVDCG0h4gtCMGYOQPQGBysSjx4c8ghpMlw/
oW10VxwDNXcU8SV3YlJbzsxlID04DlfF23jr2ilOG8XvnPPGVEqWFDuU2rTg
xKKCnNoTHhzAF8bt1DZvydzz4+BgIZEeACT33bc/a1aT6Z3md2xYP+JBdlcQ
sJmgcbAWXzr/7qWrvRaUOcH2t2mKGZOFj886VIzNo7qxTgQ7Ttv/RB61qLrL
0UsyNgklwiGmxjTIBYZeg1UtnIj4OdpaaTotvyQCpX70yANBD20GXkPGqAVX
C6SAp2ccTmyTzY4RW2qpym+Gdtnibhu1ueRwX8krsvB4paFDjUQVm90rEwi3
nEZhOH6ucyY1Dz8B8JDPRzXtlyfxDQnlaMwY4YbffXb260iTbo/olE6ZGvcG
JG0luBV+IRNpegufgTF9cNN3xQOajdOThrijAeR6Kdb+rKfu3NrrS8f94Lls
Cmq8iO1d60awbg0zrVXoV+3qUHP0IEYzJAwmQWumRw8PbSKsrC74hWQTrKS3
TTJCnq6/S8Hhj+Mw6IBcGsPi/X8qmqjcyIoIv+pwiM7Ao4+HwTcdABFA/F58
urNfVCnc0kvFSwtNvrhrfdfLErkMyq7eg95psFsEdqrgyab6FdNza/blGtlP
i895WZK+tjjTv7tiEJSZO7BVi7/l6JVKoxOKmhRtNcNd02ypsj6FHlsjywuy
1Cj596v6N+M+DnzwSHQOI6uMx+7pRJegPYI++6I3wr9CxSdu+dyVxn4iC3q6
OfiJyASrxr2axJgB8unZ+6Y7yp7Cqp0pSnjB/QSfRke7x0XwEBSLDV4rT8eZ
gHxi7B4WLoHQK3hlRofmxKJCbbZDQALzjM8T8a3JFa6qwFWKTF3QxrXesNjZ
7JTDkOifKmjRMiv8hr8q0lt33a71Xq4wWURKXyinoZ4B0B+f8wVlNSamoKCD
mhEzFQu7ga9O4XT+7uF1REumHL5HxqJ66stt+pQ1yOTa8NgQLDDnPXisvPYW
V9cTPm34Xv3vlC1KE5DEas7H/beTbcsOmon4Pesdpy9snGrzDc7vpjDhO8z0
yoAvJwzBWn7swlsRsMq2JFq+W4NMJtHeHs+tc1rlKw6JI4C9g6ju1MGLaNOp
+4hLaedINTUbtEmAqBfYLtd3JX75j+wqjlFfMHYX5IDfo0VThAmARVKKs4e5
Te6OCtK9BMrs39EHjvXNouBU3Z63iLto/quhAA/bRqrgnsCaZ70APYUEjdiL
2H9g3miyu0YR0X8Lu4d71C+Wfroov8EVb5Ct4KonpGUTjtT5sf7PUMGRRpyZ
JR8SP90b4dNNsjZM7KcP9LG88uDAqaALd9qp+ijs1Ji8pXX+9FApyql/ZW7C
demiW4L3T7i/fZcKfRllQ13LcqKfsck6tDPINPGDkQsMIquSGBGvEnhHeX1H
6RgTWRE76HJAvPCD5kYZr3LSet/eACVmRzFNps3sGOzeAhhK/KDwU+oYyzst
sQgN4ZdjT91h+YCHpWxOWj/QP/2uRp6n6nx3qg9kzD5WJ9AQlydHxsNlSpc7
/fmyrN9OSwIOemfjVlqs1hmdulb2jhcxkzwF1hgN30ZvvgXwRpK0ujTPSP0n
ZRA9Q6ykhDOueW770WX//Ch+QVn2bbQI2oEI7xTP2HMfmoGQUfjSyPrFATe2
d/slZayk+uAW9sjj8NOk6A5uMKXq2Xx6Hq3KDc0mHtvYGxgGqxZdq4zv66qb
B4A681i/6StahobLJi9J59WG7HWRDdZUVYKeX5d7ARADibKs+a1P3sWzpnO2
ywiBZVQqcSdDtC8/az8FSE51aB/ooArJJuB/uxTjoD6p3XRS5pXIXIEfdUdC
QzUnBku0Nne1zIrb8uKSgNY9fcX9OCgcjEpILhnNSiIZskJmnArbyI92+Ikg
Zr9H8JTC/ki08UozJdcKe55fBlEeU0wQgM6yn8FtJS6e+4CEmsmAwMcY4BAj
otMeIzovUP4HwVXe3/kv4s2x2IhycfX0m7WAe7KWJdjLmWVoqzNekcL9Z2xQ
jqKCsgrqBoh82AL5L8mJRZp5hVu+kkg6hAKTmt0x7NVHZWob/rObsbzxASEv
668PvhZVzM8xJnO/nwjyzrWyy/cxg7gWK8J3xFJAlnXjRQOEEw8+M4i8Hpa+
Jgjsw1KS62dgOJZVMgc9/tRg4KEsRgGwvuBrxTjeT2VsrtPWHWiwozRU1YBo
gHp5uM1gaT4sI3h/MeDJw3NGIjA0uhtEI5Dx1AgP+IYucXoSphoD59e59kkt
QGKWGQ7InYpLEZUmE9oU3kfmdDexULsTzU+smUnGOMAJAIiUgx6yYc8GivZB
mZcEFBO6b+LlwvRktCY6woD/t+vJmn5sBdbr3q9lLqplnA+Gs+3wyXa/frtU
BmK/b7Ipku98n/EPh9xHim9Asj5rpTYe/narzajtzeU6hGOOu3ukwWjVoXKE
e/mHC3Y1Kh4onTcO0YVfnZlAQ0EU9r92tqhB9y6IvJuIq6SGi8iblTHR+YT9
sNoKdEQndghggGvMkkBPf3fAImvr8NBlwSsvyPArrwn1tovvB3xh1Ee71T0+
ok/SWaDVQkYNN90gDgeiFbui1DHClW9yULG3mqWi9hjcf7aLZ7aJ1PPw1pKt
eKS6R5xaucB02/7ZdN+dnGWtfw446nKJGy7NgNyYhOAiamukmMPhJ8OgJa30
S0w4fc01CGSmxoHRhPGgap58i5jFNKJhLWULnNN5MaOpgQPt+znOxnZ8EQsU
Jij4PkJA1qvUtGbKwLzrTuzA0prDhNXcD8dj/lBLMWicMzfkw/ugXNxBkuqU
LZiX1/d5rQH2nqN1pW+pRh1TWdW/ayjX1TJDESHPuGidA60OPAq7mBMvrDv+
egOxRaYBm9fOeywSnZPMXq3n0H0mD8atqUsnMiDJtKgJpRUq7xdFAEwV8tAQ
xbXk7mnE4xFuCaprpemi3dHslBgz5yRFV5+MtG62BzeMEef0R9WYHyRzb95i
YDU99RVsqz/hD/d75V8dpzAqQ7/uTTMy5OBumQHITAUA/AxcTBudUD5vHpdI
SbGGgqsTmSFJbqPkLwhAdDSGoJsjt2eI4R3zGLNU6b0zXDK3ZK2j4EFnc1Vz
nsujul7tYltq82x0dNqWF7dKFFPvj9nHoOdfxVBzpA/y7SKag4Alg7prBpqu
6b1csypvJ0J18WAXrB63blzBXp0nB0fgVNXOlKX8Ak6vvGGIWgKoXbIYJgmr
jCEvSCJmnLv5uCO7Es/gokpJC6vofeCkCbHJHFFDWelfJMNmFnY6Fo5PyRUl
LDloKoJadcp/+bQ8Vp8TZE+7ksFvKrKRYqTVC4goAw7oHSwGHUxO2zh/tojD
2w1m1r59zKEnGL9LxicN0sU5VPLE2Pjb0oAm2LGYE4Nc1m9c6rr6uvP4EuNx
KCU8ZC8kBnNxrV85anSq2gH6bhI7/HJrsg/YK/jby6r7ye8TcUYnktljDw7j
HofQ+if9BXMuke03m2ujiOTq+cB74zSrw4JgTeA6Arhd45Oek9LHa/Si5syN
rjtV3oekzCxmUui6+HOuVPTdGtb4PEh/n2phM5JZDGvJT1V2khZZ+JZFDZgW
s06jj7yyUdCUDa7yXzFrs+UETHmeHxhwDDemXBeg+zRv3eI0mx9z2q9fYJIF
aL+C+2iAkGYFnnwYb4/LYEDfY8CT3MLCr1IzIJrW5r7FO0X2QCndESeQZSZ9
0jzJhEXc1OJYc+3Msv2e7fBCWN8tHyoIsDjp+QScM6CZQmoehj3qyPgdvR0k
XjgA9INIPk3tDBQucpqQsSnjdn1PEfzXwjPzABgVzahhM+z61RS2oeSKov67
OEDjUBAy7xCSJXL45e4MnfW0u4PqOUw0EFY+inf3rr6k8nQPjIee+LkJqGvo
zfT6M1K2tYhstOn7D38Mb5/w0GcCYeoa3EUU7LevoKx4/rfM732Zl1+9jRqm
d12GujZTl2wq5KT4iMnZ7bOmL8+kwTvhQ/tlelXmL+7e6X3X7UNzm2A0szXt
PpIhG7WtUUESijN6iR5GX8ALMZFhLkCmvL9U4M75cM8q5w8Gde0L23KKXVq6
p/VZl/+olIWP07f8NcEyF8CuUP4BsKGAMCyt2bNchnA/q/N6lxlKSYYxKZTL
iJkOBjN4DVE8Xr+LMGfYz/roZUZG3qX80/UtgBgF2E/fNAHDqOVVjC8iDk33
Y1y6QdSoFKuIB/QOqjZRYv3DtH/xzauZV4MvuAOA5cb15AS+E2tvIF1UPTZ8
XzO653IinUVf0Fg5B6VMnofnCY0fnB5G0TrMh0tK1TPwjB5mD5h0VraeICkL
g+W1rwWjlw+3YROuHWlp8xEwOz7DYF7xx6RzpLKJ9hKV8PYuUcPlHDdq67/K
Us7KRWZvMa8VJq3c1zOBkdhicyjpPITdHRD8GJVLeU1ijdXWKoh1Eq9emJ2j
sVYkEpRBBrR6qMPHWuCC85e5yBam62wyjNQQv8Edj2s45i/Ar5c/VymeSnIX
O0OV87duk3SAWGrBi4e0KW/eTJheS1AZl7D3QdfPqEJEvjnoXFoodKRyUZoN
A6hfYQSYHA1kYB3amq4aWc5ZBjxahSu5DKG77BvTINc2aPxKqG4bNQm9Cp8l
tYZ/5dKogRLhNBNlltg7a9pbVjQv/iEsd0pzqwAy/mTkZrMqEEFY/HkAynLU
I/zmbMwwQZnSXMOtQrQ6SKx79/22JuVZx/OOlci+t3VEeppWwV4nNFHoaseM
Z7ytGSets150DlwAnJg7iPf3jytQY7ofedBphbo9hvDtdTL037PBiUYkEiQe
x7IB799rSclvhWCCp2AkRH4eqVeiIPPB9drr1/UhAFZaZR7OpvOJT0qIcSOR
htK9z4qwWsaSTx05glU0NpqUcqWRdLO7xOnqF1YCQFmXXuxEEqyuwxAjEoPP
AwudxokXGzmTHoFEuDMFfwtKa49k2MWHb3gDAW+9geKxmtn8RYJue0rBV7lv
zENBpzYyR45CmpTkG4fhTEXHPtlvxnnUUosfu170T7suCSoRaBPIrXoMHOvC
5zo3X3vAoiv42ZquW5TrPr8vCPTuB7KCPCbP7EhORhkXb5+V6avoqwAhjQg/
7hxLM/ZCwW9hABBrjhHmV8RnLhnNA0fDt9wDekY6bjJxO8U6hY8EpCQxqnM0
si65KTiY5R3eCFdx7qBvfmGNjQBeTIL/Fd2bBoa2rc23QVrsufqlmdlrR2UN
pp+v4mnrbr77AHKsnGDoALfvwdHinBPMwGbC+plijVTy7E6SLJSHDcNVQ9FB
e6tHPkHus2DyuxbwAUCnoZK5U0SJ5CUZNzdkN1LcCktGRJ32JQ2HbuXZHNpL
Q4NS+SPP6REmeYVToSkC/Iau9RrGF7hHinFUelFiGvt6nLRtfjbokYEPhC/Z
XeSiAUnMsUSSlTeaM9tuFNCI1IENisQwkz9/9Epk9ylHExI4MFADCWutk85F
Att5TAbG2ZUWzwndiD8QpM3ayzjvI83LxtTijCiBZRazrjeCUhn/iTBXG8pC
kmCBjuCuVkkgFfmUrpkFimEjg+WQGJ2RSict0LjDEHopI3fnrOpoJSGNqPmK
MfNn76uISxemOe/g2wH9xZBI9nkFd7qsBb1/Pq6KBL9haF09OMhjXYIKbI3+
K0CfH1fl9dgiyWTCCckMiJ3+xRwxWEkZzudgNwnW6u6RgG4baUsjaUi2k68+
u5dM0GIPf6rLYdQmcfAD+tWk3Fpy8yJaLeWmBLSXpKt+CeSSK+Rb2YtJh6NJ
qimGN/Qt2Wy9c2E8KUDpoZZ9S2yC2StLqr+BEu1zVoXPPw8D9YAc15OuYhLK
3heKw0mtuPQNFIoe/s4POcJsgdsf0OQnw4nZkNiIdHS6K8uPwe1Fa7uU/199
KTLYOPoUgh95omNG+qHCzyz/EgimPfIeCMkdCjEu7zh6fJ7UqWCiQGeT21GJ
tsa2sra4wJDFXkU8QnBEk8dpBaCITeElpwQc794dizMzvzcHenY+5aIClaON
V3YpPk+9eWU66hiAN6/m1M233jaiukr2Zinw6K2Dyu0igGUxg5GLW5qDOhtS
idUXR52WCnYGteRyFdqcSFjqNtpzhoZNPijfLLHIEdWeHOAEOfWtRw4VuVDQ
fvDGtSKi79Q/1jeIpbZ3RHEuuPoncSl8eSPla55QC2XusgLefD8+b74eiN68
fndLoNL+UqIY1GiyN056s/eVIM8TWcScdc1jDB8NxdvAWUYGQB3q8pY6MP2R
uLh8Q9tqmxgD8mYTfy2mzTDSKuc4ERfrM9vxSeKcb2xwoo5cyDUzLHM/0IRE
6ZWpP2DCcw95aOccnd6aon0VXBAI7Sxo40lOddc2e3HY5MRKUhSSTI6L+Zb9
Oaeay/pY4yT1ueSZms5VJ5mqx9ohMRMrFt4gY7ikf6suzGcRZ8ffiOaV4SNu
kHHZBaJ2KEvojfGtOfIb+xfUV5q2KX+TS4dOebc4hTjWOE8drWEuTldn79FU
xcjGOLRov3way/i6GmdCsFc0ZFor+pjqAThiOPM8QDxHDOzAvW9HAw2AiiHN
K7bwMzKL/zS6fXu3i79PZlh7Q79fdyrGKq3S4lKBjluSd+mqCCjZ2rjG3eNS
kmq9EmRSOOZSdoQ/VZQ/6G8q0pYFL1o258A8tg3yoF/A3O1Y6kpmFauj3Gmk
tDirE68L7WSM7aw5Ed5+sGInumwPGTF9pWbPLCPcS/Slw4FGeA6Aw6xd/KGE
XluRqxmpCNDCumjy2Z+guSk05Isw2/cNiPK9iJJbZ7n/WXcdFCIctJ+xX4A4
0n4upT6IeiLvTb7l7iFW2fDJPg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+kRiHS5X+di5VLAdy01N6UXiulpxcIX0037JVXFja4wpap0CXjd3FXIue451WGozDb6v/mSSazZoyUHkCryY0uTqzuS9XgHul4bjj6/3sySt0Uvujcg++YjyJSd5/tdSfxNI/vheE8ZE7e9euOoCtNw6SJYBcoqpNaxDqwavFF7PTSdf094X4MQgzMX8nHpAU/NQNn37KnE5k58Yxxnrq4klb39lfNVv+NyjZ7RZ2PEH/OHgfhaykJZn8civrM3IlfRKQIkQtVJ5HQlF51fNUsCSyf/LVu//VX/6chJUI/W5d+R9QGEEZeKcIzA/EiHLTaSXeC6Y2bZaIcXF3fYgAjflSfyONrS2lq0C7KMDJAdi0I9keEriDfieSoPGAL2PmpjdFBuGIufh+xSX/F3l7a3aJ4XPLzIB4G+5JVjarWBHV56gtBbVLdjNonTrBLmFtczAtIqAJ0PNCaDO2ai15CPpA5sdwWCH0qwIz7xlN0xWAONrSeFQSOZEfiCIJQ8WyWvkSLQYkI3+MB+aBV6oDQufPaGr0V04OJfobIDjy41eVzyAtYSZuCvTi85dFUyxq1hwGVvpmDAK655GzS9bNWVe7G11u2WtQyFtjuloq56wfIufYhJdR3nc6SVyqIKPTJ6ZLmzW6Iz6PlRu3rEB/om429katX3kzxkjnJG8DlEf1geZ1PQKlvgagr+k9Aem18Kv5HDk69aWtUfmyqqs4QUeSZnFLn3PHPeto/Wj9+tf/SF8BXp4TVd4xLdLO2RsSzXn6eaBYFOeovURXVwgCHB"
`endif