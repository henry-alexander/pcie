// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rgLi0H01ojikG4kbQxt/RJPjT5/XPViFO0v7q/sVw06NVVuRE18E2wuzBtPv
kD6Q52Eco1nfJeZ8ufalGVeF01xUynLSqmjTH1ANNVAd5MBQ63te2Zvg+uqh
7G7CGSYlDr4stv+2xUNLW5J+kycLjgR4hy/6YD4JcYFB21bD4qPuEW9cbqos
oAx6J/zASKC1hAtXYTY5uRqYkHhN8oAWmK7upjvaOcvW2R/VgSjXW+l6I/Cm
/b/imjfnpKT40RI0o3M5uPva4JNlp3h5ek64Y3N7K+0JG4LPifTEwNajPPlP
2KzMbUQrE8wRFd+gpBvWag6YgBesCcRrf3zaNgUMWA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N3fNmI0ZbcqNNc1dov0ItdSzeugJ5ThXBG3+w31VjH7lr8mnRUgyY9nekNfj
Eic+54xrZFEAvy3ed0qE6ubocMaDn2jmn8ZgKUEVjXF8snjWN56lZcrtIavg
d4rHdJF636rJT8tyNh6f3ILGz+38HttpAsN/w5BEWHCZ2TzP3L1JDEVJTUPg
jASR8YML2J9NnQulK3BwM3b+sk+tspi5JCkiyzQp5MLq6cuwMYHU+r+Loym5
TJwtJfRuzB1q5bjNEIfVfrouEZkQl9/lCbQ4c5d4qT7khN6OdkutLLGASXu3
xe+SucBuKw1uttQvZP31PxKBQ95hbTpTMBZu2to3dw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cqUcGT7/2MlwjCH6JlVbhgAcMuHLgaudydc7oBoQpxqdqISR9VBnI5/q5+vX
4KECP4CuGuX2kixYqUPdM9Mz59P4cnIRhK4f5UwRHYVh0kslsYYyUTOMQ93G
5ZCEQ0gGvtiN4nbjB5Vcho0pWKZLrONNJKkmYFeSZNwaFnB7n0bT9PdrvI9c
af5wQ4vjUmoEtZyTXy1kBWTlvskr2tX2OlqLKVkbPnmYFso9dwjcZJm0Ybjs
LIagTqmz1g6Zvig4KCeZivs9a9p6MTjFCnDcpnHrq4QBX6BJbWNlIuoOBLCX
X/vCAyEVDEuSbeoTmbcL7F/8MNmVn8R2kLtrAITPnw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GK9CpEf2R5HaginR0kLvzUsa5HfazhdaqpHeDFsn3q40pEbuUhvLWPGHLqFd
v88eeKL2uTFMOf0LW+2i56crM9l41325N6SPsyTo8MiTYBrHmhME+UtX+1Sk
pwb/NuxXFEdjzFiWSCZppi5KdEkJs6nYlnWCtUMLAfnbAdBBl48=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
L5fLQ78m67HMoc+qowb/snB4I97QjgeOzic/vKrgYEldU+Ou2lG19pIZELzM
+GZAb8W4rgw0fBcnIwBzmK/HbKZrhh9Yi1Z6WCnV1ha9c1ly3G2F0ytbXb7p
1U8vHgZi8YSdYHkWijAh6AgUwsr3NVoPXLn+7DmTgZfPc6/cLZd3J1eU8fM3
B8kPH57MlzAiKw05IWG1sd0XtmVGUUuDfjm5QY3Q9y1r5Jo8jEYtN3EtP2Os
7T1O5dkj9/V8EqGhc6sUKhRVYwPYiADUWFkLpNEdptHbDicz18pOkfY08D1r
9sn+xa7ZhtzirI2tw3LJqD9NLjFGC14SuybpZC9j+3TA759YFlGmHYLlORW3
r1M2/mExostWleSFDitVM4roUITlTjxsYuXUI3mdxh0A5D688MY6fM50OWXg
dNghAZGwHVCjD+MMq0/CB2J714RB+aIW56YYeKGtO4mdv61BgInJWs85rySZ
0YOssWOEOJAXsnxHdNWS/1d15NtwivXF


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
biFEFDGIxE3uWlg7V5Y7RrC5bnv/cVXFjgsCBfeA26SV1jsF7McB0Fy2zOx1
kaMyuOSKqOKBc9W1dgclKgJ8CefjhpQ8B0Opv+LLJj/fHUxCry0a230jyflL
PJD5pcNvSRTQ+XGlvtuAyDwwMOo7oU6aZ9bhVPFfGHShS90Dubk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WBUuLUTZwqADEIjC9kr+8T6kFSGamp2gtePuZwQWOwLrtn/KI92UT51CBg5D
WHIJWoKXeM18iw0SIDZyFxABvac/O137gF8ZhrMgSi1CEqqVaRwtVOSItIRv
cSAbmyEIJmFkw1RwGt4a4DP/Ael3A52bhI+WiRdfEvbGQVsIpk0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4592)
`pragma protect data_block
WjhCxhS0IDEYH2C/Z8ARxa821qnF1atRh5fqkL9w5dbTYXR9NMOSuelU2tTI
rKo5b/RSQDYJ/4OmnL4abFi8f22VhH9gCnPDboWCvELA4m4bRdMnGo9fMGfG
azWh+DGxuIgDS8CCmWjuAn6Z+FFO59J8Wog3h+Mvv6oTXjs1BnWHTnPbleE2
jNsuK879U59DFGmhHKRNqyyvFVWP39auQlsNnF/cslKDYJyk3M8opv+biPkt
R2duTtsfNgdY7EM8S3HGpWzh6EOczDLH1WVXpblSxbVRGlDinWUCSebDqk1l
IEBcUBoermGlcqJh5p2gJUmfNPUTtFAQ65Ru4v925kJEa//J5U+yGrxWEvvb
xfRCAQrZHUW4dO8ySPW2LYCxzlRUM1qwB/5OLQrhtpRnRVI1sRNZii90mdEI
KPtQFuFWIg0PWK/h/6lM492AjplzYPWPzg3aQXTh8nbjkPLQtq7qQnsULyWo
FkV0kzOganvMmmphKp97/J1sWX2LueGG5mMUAOlFHxFpp26/xcLw+uyo2n+M
IuCc4vG1afigEVzdjGTn0kAAMTsy47OtGZBdPIDAQy8GuD7lW1DMNOOiDm+4
Yu55Hr/644qbjUm334+lyQmbo9ITwWSQu82m+ugrPmenMpkZXU1kA/cYhot2
GAwZ1Hs/CKBcfGMX4UTVk8SB1FznBVhVUg7zjnufZL5itrpeq1yXWhUCqpd8
vukxAyPYAfgXozacwBQE+UyCVVJ/6Ap8f4u9WJ0nO+WFIRuagHs/AoxGHvzQ
AUmBUGdEriZEOhHcfgpwjV0I59ehTitsY9+4jhCqYbfRJriDyTcOIi1nB5wJ
NeuBImkZs15rH44c5pBXD8azEy3YfhF1qy798UQwFx44B9u9qdms8xFYGPlT
h0XYQOPUJ11gfHKXS2k9FLpQ51JxPjPBWHLZlsAN6yxHZ+G9OWMJLGPn9qC4
NggpHTGY3rgc/Aglv3USKr4OuVaYooNrDU65Pqhp5Zc7Mo4GCADzGzsWAiWr
annIE1XLtUPiFryAWyvqhc+B4AlmSyRwkmbk0UpHsd5hYibbQiCMepyVgvvP
8WIZcqwumpnF0WqWWPjfS6HvPy6waZUVTPhrdjcBru8O1xZhd6+8/lW+rAjg
U/xE3PxS5+ggS79Wr+nR5UphVFHrrfChNFPHU70KaRWVadD3OGCp5SZD/BGP
NzBpqNwDHuPL+fSMVU1RarIVHIIgp7C97QJgq7OJnhEWuo4dkSKeexFyGDUd
Xq9hUCVTm9UYE0C1Ho+Sbxu7txAJjuyPnFkuEqDApOlVbngqGBP4FvSCFMmY
01IG9O24cH7duQMJYyJEGYUpsvvnQDBi7l+9tDqvqLxuod5wNB3x8OU8Fn3l
txWFfRaameNjLjPqjRekHVtj1HKgb3r5tcmEpJp9eG9dzQq8cQuQ2qKc+oo+
YFYOCQY3/Te1jbB1Zn8AwNfMrDLU6e4YBbKUlaCG3BbnZ7owgWaZpdz0YOUI
Kiwk6KAeoijQss9KtPqQzSF+LJDjCGZB3iWZFa24fKxaYIQ74H1kaxf5aKGO
LgAutE4wOEWFbd1hutsJJdScutbb7RdbNd9dyGTonhPvsnzS4wkE+iRRaN35
B0WhbaMK8Z4gmN1mdF4kXJ8QGwPVxVl9W2pfmEeNyNCNbqP9kd4khDI2JIjP
iimIxLpyPaVVhdk7O/EjYMcG6IeDBwoQ9FNHQm8Es5hVcDwAjVslV4u0kdkb
X4o4QfurfQ9yvNdBwlNZJORRjbdUo4O/Ot1nA7f3bSj7n7oecxUxEdDfm5DO
Kt5N4cvrcLv38KNYXU3BDxkrdRg944e2Z8SHLkK2e4VnS08SsWs7BAQ2jheY
dbXCenr0IylZvSmbX1r6jxPq/si2oYPI1/kJbIA9VohQ5bYN9ibOWXTBxKtX
lCCqRccFuflw09dyvvvyhef2WluAinUYl2MjEYmb8eHshBSYxJXkAcY7CDIl
SsqCVJE8d461CrUWXQ1Qqsvvv1v/2cDyIR20D6LfpEicX4PJlHQ+7egSV85Y
JH+DMaQsvMSfnzJLOIsGcT5Hq4TpQU60EG/L0q2Ee9X5ybZ3uvgLec7u8W57
YzmrvrGIESwb5kwmGaRVNCRcqZ8DR7wRWsBmDI6M17wFu+3fgv0qQaQVuS/M
1i5XZwhFDFiSFBES51sP0eqT6r5VdOIPIaN0apj05f2RnYcKZiVuz8hfth3j
uCnqCFMidFrLbEqJKscbm3KkfDYtRSyS5m6HXvu9S3w5Ad77yyYd2cMdl3Py
HyWe0s2FJNsjKsuh6kvPwcChDqSKgrvwlAjcRGqI495a9zJwcrRQ5qf8te7N
3G2OlK9wri1tPGDzkCiPEi+cFwffp4Az2CkIGLkiIT06GvoxGrIclcNmQZDK
hyjCw4r7DA4vsbF8h0jxZcTgjfRPToJPMRKWZBTXr4zTNTqEmOU5DMOZy7GT
mF8M+i3ey2sv2UpsiwEAxQNn0xPiZ7mqE2mMIRcdsg+WBDvjIKIvse+HEJ2K
GgcC3xdCgvJ93QDyoFDhAPQEpfn8Y+EhwbY97N4A4SlxfPUDk9gr8+6q1GBh
4kyMUedODrKiUFlj5BFUJmzT2gPquaClZC+pD3bxX28itBLnshaGJHeOJp06
d/o74VpOn8K3FnSMM89F86s2pPL9a1GYsxv2CVY4k+7Gjfnos7MgAcc/zd5R
8cqVhAAp90Ay1LKgKgah2F/9hRgeUT7fhZFonkm1qJkeO6yF4a0yqm1Wplg+
fg33NuaciZfwiAloJPo+giW4HZ45QeBLXUfTJMH2W7cJ8oMWIhPJNUg9yw7d
teJQV08ccbw6iMSBVcTNmP5addYGy86mVO3H8R3fqHv4S2sV1obbY+O5wI2h
tJLh/IA8pITnHvmLPngJwRBKR8q3gU6VRmq3a3Z9bahHyARqEN7WyS/fF6JS
1MetHZN4r8X+sdZaUwKtESIe8ELRMPgO8iTD9XigWkf2RukkpUrpxxpUFG31
5k8mVW2tMHTbGJ12Ir9e9a4dMCMX4ZCCcacgC8B3QiErJ6yuF/Zlf1Q3bClF
9qk9z8Mm46XuDN8+JyrOToCzM5gF1lbvJ3FrZQTC7k4eshIAiLYzKqntWGVu
r9AK89VhayfOaWC2BlQKHIgT7496cUzJsGUXLM+Bq0uGF7gbsWenwadLxAuG
LXSkORip4UkLLkWqPIDewuJ7qeuSHJV6cRDM2UKsheh86yhUxHpEg7e7gBo4
iAFOhI2gIKEyhg6zwzEiEfhY3quZiudUpJLY2fz3SD5GRjLmArlA2u7IjZu9
7/sj8BIju0ka7C67fxhj6u4tt1sC7CqLS8OVh056nkMFO0pFWRCwMIEKFy/V
9I5jZIqEXag1vB2CNgK9OfD0leVz6mpnvuE+ozHR2DOp54rP8yAOHVwygiWo
MN/53hTmmbNo+tDzpSR1VxFSfcBk5YJ2GBzOwy9IRyTqIfL4PbBhRusdFiqh
20/NHfCBzEXavPzE1tfgMHmb33iTbf9y6Abh8LGuzRektcy3Cl03ZcEXkWuY
EXiXNp+jikg7fhHPnpWikJXY2ipxFzlc2Yp6k7Z9e9KLbmVIrE8Bq2e/zKav
3HN339g/7MFWqx4SmlcLbOVO4lDYMgNj42Y/F1q767SAfBy5LvjmC2+5Zfmv
L1QPJW14U4OmwN/FEz/ihQZEnUw2f+q4albIQ6lJmi2yMym2g0c5aCQDqeRL
pWdZzLCggU7yU9cS6EiseCgcih/ASOlY4Uwt7I2HUhEa6ZQyh0aUsRcctVEN
p0i5UWgWOhM8kV1l38GPaKjjlzYLcZqE1sKYbfB+AogZQHcJ4SdQy4W3zvUn
rWpgyu1k14DVZavUAVg2/rxKvOKUNQM4sUT/y923P0JiFVUX5rSpFtixEkYe
DJfGx7vX0g/rO1rGjDa76e14Z4dYC7xJXGjzBft/NT4aMdYxGXsG4dYBKEW9
OHYuCpYQ+vN7O6FtkSP2+o2GIezxlawPIDnbIve+b6MFQ641kEGTzxKgc1LD
5EfANxvgNq5yA5ex3qr4OcnmC/s2OXa1oKr39cF8hR0WTA1ICHIiQplmlKPe
LiEmjfVR5NCbvrlk2/YETsA7n+1LPuh/LZql3XEqDsHEjSA9d3ZZtkar+UDz
yboO5gXLjaQ5X1AJMRX8+uPbr+YGx45DAwTW8BV3cECWcx5YBpIlg58cbyqo
nL+RdyQdRaWu7TzifOMBXZQQEGa8MbFa0s2hPkq/mzDz2+51uCtmvM2yQWlD
FX8Egp4BDVND0sHC9m15x6kl1AY69CPWfwvp1WKP5ksuZwMDpUGFS4RRwJms
zaVB2edvVfPWO6HxZHjhE2dgGa4qWsEeJR4zayiYUuCp+ZP82oRONdbmAQ3K
pJf10PVjdoWtNiF8tCo8wqqy3B8G02Wo+HaG2cdxPhkIYe9UUIIlkzkIHZRD
o+4Bnsq/IIm0daYui/3ofc/ExuyaH/Q7W6em8VCGVn0uWEoevp+hSH8USyyt
gIgHhVMKMX/8E7Ezu1ejy+0MIIh5AGCoO0exRzIQ/sZWH96X+Lc2FYhgNQi5
n8kwoSfSzLB4dtRbYyzglvfXIRSDkDSAIJ0jh90h4zQhPOAwCIM4juMgFzYc
jmjRODkkL3IxUNh6S7EkgrNmbIjf6WyPhG7UbfIavFxR23mbVafTZmObR2p2
Smo1/tSd/iFMC8MBZbVeKnYlyjoNNegzdQ4tMZOy3GViAVg1bSfo3T3G7ULG
PSz5FhQutkWtT5gTprfXme/n9dyOg48HZLCiU/rFk5ERCMkxxGdY2sHfbL6G
m6U+ozSBCvPbMNe5gVrsrDsqLvhawebRtJASgaOJqFhi8DGi3fHrv45WbNnY
Xm1vYM8lEXlUEXFq5L5THpvYygCqPl96z3X4NeyPd//WJxqAvzScU04DGkyG
SJpgu5z6uMZU0e3NN0PGs3A5ZuSJVj3xIY/+4fzqqg7rPYmntv7lEHr2oh8O
cexjwdC7H5hvcMXomwO+dZ0GUHy6ta2PPquPooGXduYJoJih1qA9WDMIa+KR
ZrvJyk4fj57RKcKsX7qMbFoPbf3unHi0HWFOQihVx10ASn0DLFdNCMKEUmTD
/YTLRkFP6iQh3QgfX6ScdX/N5NBI0jOvf6B19TK5gbfot4bTmWtUS8texl5U
LMGfFmLjoheE9o79IOhI54jI9yUs/QOtr0QQDu96OyGcX0X1wGSTQzpqklLd
FbISVkpb/FfDM9MdGOnQbqZEGbS2LUpbdNMmAZnM4iYd0zChTWzzc5VgC8Nk
tZN7yn8AsKKfHFSmbMMMmHEOIPseCVQoW82ByVBPQU8rUFZ7YHAf+wTMIunC
9d2vqfTkT/nY71iNxF3IWYx24X0dA31TmtU/1lvEbtRHBUrGPsJYFVHEPEQO
nqKJxeK81elsKWX/RZGmOkD7O4cgWd89ydY7USHidw+HFTrQ2fWrrm5bSl8d
VSNiSYH/e9HyTYwhmiQdpq5y3froileRG4O2SYoqgMsTFFQMdsExQDoHmIPY
IGlhksMBqkO4O799YBCpOrk/EqJBRWzdxA80zhFDVs7s+bBA9fp7AP+wdARU
gGiI5mqJ4lm6m+djcHO5vcGK5bBhCDsmm6jJAxl/8v/2FKd44g/G/qjnKO6+
9Li97YZBWttEJlMvoIRSUrvsQH0FpwKsfUwgh7HrqEdRTJXy0yQ3vztxA3FU
6Xtm3wwyei/F6Zeam7YoDF/rPgAmHvNwjCX5m/55lw1YCg/piwLaiwTPjUuS
DMgQiI/EqPEs+UJLVF/pgiJ/I5+s/5zEBRKwHAwinE+Tzbg/GdNDDHfE/mX9
hGjxam/ZJiOCgTO9md3cm9YEgVrgdxi8FfkrBRmYGNV5v2zW0+ANwyafNV32
l1rg1/C1KBK2gr5t3BRE3GG3Fz1xiqdcVFnJeV+DcoWQtDByIlc3hhUOaNaQ
bVJk5VAyLoohyGrDtXBWhIOFlI+GLApFP9QnbVljhlT9JAPMw8PxfvRk3bjf
x2DL1CL7g9HOm6qBKXp6onFGYe/wZAuM1V7WusOXeOdj4yHi+ItQn1HyITDb
YZWCGzAjEf6bx6U4V1doYmkCTPUWeMq3dJDrd5+Rthz/QkCa9PJkOdYNXp0K
fT4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3HVvpl+SLSQTZiP0TbJYaX/BvxT8Mu5cSEA5vcyatbtVhnrzQBeCyrly6/s4v/f8b67BQU3MllPC0qHNApQCponCMBfpOIWbqe1eAHjYLySaj12qlqDSZIkUHfw0mi0mb6k1cjcJTOPhp8DReqsKllk1T4GwzACKMaoIzjEhPmIyLt8Xs4N13LpKHacAdO6O/mJcNYz2D9jOuffzqGmk/6CgH+pZaGi9NhSZ5VHwwn82396daNsZO/9CPp2Q3luTPkEVnJjVzekkQHB6YTa0vUnCfjz5JZ4LY28yTofI4HW5aHGEKStxIx2yunIr6IYOfS4RZsMrIWycnWHQR3/Wk8pMOihBQE21UODP5+ulGCSIzpqKuHnzkeY8Ttlj6imAIFvAqyR7ZhQ0FdSK2KkWZXfmkFKpZbK7i1jRDLVNo2SYxwBVPx1WnEpV0kBHNUdk6skdUxBVEfulzDH9gIZjECXnWEb6TlZsg4knddIVHmY2BBkLiM/Ep1d3JxW45tAHf0TOV0M4Nb5/pzmRN/3JwOx8xmS3okCPTFIZckhgD+syKOnun620N8is5Uh3Pwy6a8M3GYM3Dp/jddRgdETn1hYNByO8OZLX1uENARhTjZws25jGT+ghHbzrXgmHZOtLkiMXp4G6XCDo/gPz8yn0yLmLznLn2UdyQOeEusQYAfMxYDIYcbwQWuWFph+YPdf/U5hk5LJXk5hLxGzvjOLdzzrNP//5vFx2mTJvOzu37MozzXefoSfvGMvYeTs9Xmx2sbJRSdxUhaxU/o4qLn1+sFP"
`endif