// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
rmGSTRGtdfc/53ixeYnun2fFjGirChl/+K7wuHUwnCyNsN+zqEHsQDw7aoic
vt2ryWIgwAgqeT2bZpA6HYG1jmhtCVltSMm4+pY6eR6+CgOVnxf17Fojx5S4
V7mOfKww+qKRaCxqRCbQ8hn4WeInscxoniM3S6bxqvkF4Ev8QZFnSOUuNHjs
QktNCYvQDfztzGa4X4Aq92V0R+1pQr2i2cB8XSFA6EqYsMOjOSloOLdgaRPd
gwo83teMSLY93vVk8wZ1z8DOYuCmbXyaMbiiLljEOkEI7wBPeo+9KMWc5Ac2
9qbdQrlh8YT2M6J8CRwkUQYHgAo/7bMXKwEt+RYH/w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MmtCqEeiOG+SAqBRmh9dtduUmJkoYWzkGIhbpcnmJaQZuM5MLTDrk+o5csqP
LGYPYqhTHKuFu8RBU67ZAHYougtnSnqpehDWbjqpkPunYUqc+TJf0qo6yPI/
J+eFsOGb2vmZw1nCB+2A9GiHrE8/JYNtAEY+Om+6CvP8uvcd5lBdxUgXm/bm
cbxEqS9LjvxLB7KwEJCMbkiQ1UWVyzyssx/uXOzpcv490/sq1VdZPqZ0QkIr
KG+X0qEHK5YdMOeUDTxLbxc6rby+qNkor9KStj9AJR8mNPbM+9Y7PC3Jl2em
iionuf4rRysUM/SwV5p4SzpgCvI6yAq1wfRv+fj7HA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VphmeB0guHFCBOBe7xoMrrUT9Hwbu/nBW4Nvu1+y9ZVAs73m+H22AF1JmEHT
u/EJ1u7daTSHMktSa11CszZSKGiW0b0HpONStj4sNolSGygwUkf7nCooueY+
bchuaO98LzuoFlig1InFjX+hlrgLvWpneqsEJJzBBY5zb6MNvg/pqCnwAW4n
lGuViy8+9XasO6UzgIjIgdCY4GNU56DhsScCMxUDGaGTtrD8HeFyfqoEEbeq
NXigjk01BxRWDYFmRdoF8p3/WK0WflBOmMOZlK8IG8swHnSoJI8tZRfGjDRO
wqIOWTMLpCBeWxxNpKBcDGBVcqZBkzIIIW6LLZSiQw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZGKs+0xXN4vI47AANmz19jNoqQYIKcuJKlxwJIGf4UCyAe52NQhJ3A0YEGNa
z/Cc4oG1YqzupoIJYA/PvVBoo1iYuvbr4ZV81LJWM/VJJHSayIkTsy7cYEPf
TCOGBRQX/uy3xQCmEs3tbEQIr2EmHKc7bFGlls2oDtLzt33FRb4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Z3Mlu15XTzjn1tfkGdjyuALRae1U6WBPzncWaOIz8WL/rq74fIaIjopHR6+f
JBDPjxIZSafcW4Xp5nVsHa0i7D/zvBcH72qdADABc7QGEDJO0a/UCP8qYefV
IGNRyLi14ECUsFC5FGajknh+nu+2yiNz9HZAo3yv5NFBQoeBv4J6bB09+SYu
yHJ8Qb15vis98XSyUQma83MdGvJ0+wB0I2AefLemVAX71jko3xtwQRGcc8l+
Gk5UdHBANT2kdnYt0uRPV8oFQBkgLlh4EX250jUmgRLak0fyrS+E+kn1Ldo2
qLhIGZ2U5fZmTs6iGhOoeSqt4GkFRIWGcd1042h3jLkO4156kvzr0MlCvFBt
RJLIjD3A/y7T5spt8yNh1mOpgBwVQh3MLP+5JwnqTD6mPJ6HQH7W69b3Z7qn
bRh+X28Bwx3zBBnKCTdDNxh3UWFvqY/oLzJu0WRFFNpsgHEVWzAG9IyNkLRm
7Mf/DG7G/ehPj5qnzOjwID3yvATdgPjG


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ohZhzGj5DhUz5f+9N806v3KG3wZY/95Lte8bjWbZESjgk+NxCRUoYMOijwh3
iwHV/fPToCupNWctmRDlrhGfbFlfz3E4fskqP6/4GwXa/ETfCMGk/fci7GOb
ecfyfrmYdnOLnUxV1RHHwgH+JN+0pc1E5ws38fRDhN8deJaKlXM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QuKce5H8SZTVSmKEG4cATD346pExubh4Ga2WjDFDLlzSfOFuU6+pYfNPURqQ
wmjx17U2Qz+jelQs+pvfggHD12qK8/UauYeDsVjZbSRZEs+B/0Nl4WXUWPPa
KXb+pruL9TXn+w8LMbb5ZGBOlzk9pwtBqwtmjkGdO/c8RZeJI6E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 148160)
`pragma protect data_block
T/GP0ROibFLfY32wVtxVwUen9HlaQJDfVRPE6x4B9eJz9UW6DoSo/0QKF76Q
75HeuZBWRWJ8IGoxw98kK8CP4z+cFmGsAuRvqepU8WlMN511Rs3iYixJWXOz
2B8MeLrl9UzrY2nwVXRtJSUNPOTRenVN7D8MJl3LaU2wb1qtpCT2UWcUM3yq
XNVZTTWANTgLZioLJ2W4TfhYUNVUoPI/sCndKfz6mG7O7c4NhkS7imtSPQlb
j1gucWTLEeJYVB/PYwt77nGIBvpVAM66GOWNQbN7NV3zF835C9wS8Ire9quh
tfqHMVWf1qIm4Um9WKdWnRWuvKrs4J+ysgTaZVf0PUbnx++2UfyLVYxjDPSy
umA10BOIMbVWbyhWa8dRzkf/WlzEPuWprOgMnoqM2eWEKwCkwBRSRSgLOAO4
Z06sMfxJrlqxg3vDuIXvoZGX5XDgUjQtTTyonQroQE+Z4vGRZu5wwJk6FDkC
DtIvB7D0Yocw0cgAeQZRzR9RqiaNsIixi7sKw5PVz9ey10WvyyATsHLVSowF
i2t83gYGR47PTFLVeDkHbvXHeN6IZLvd1iy/uvNwvJl/2D45Atv610vUldf9
/moF71gorOh82xEo+tG6vp4RenesvW67YHemPmZwTTo35vmSQ0oAXYmsmF4P
Q/I4/A59byE6LOFoWWvwrAbCAgP9e2qDxWYWIhqCJQa3IWQKEtgT2EV6Ce8O
F/RKCl9IOLy/W+N9HESAcci5MRDCvSarAcAaeHgaPL2Gg1i8wkznRP3FAwDs
28qobdQ0E0CDyvzivNWIDhd0RtHgPSFa8lwMKmx5ol6KBvA38QSEIfcOMVNi
zALrBIopc+QzUTUVUPgfzMfzphVyg84bGz3HWyFtAPa+G8LaOxyI5s8Fsdat
gwHTYpK4AW8tqKzigVPG02fFQGsCxD0tlCCl59nOFiHsODjCTAY4/JmwKMra
1Z4SE4jSiB4h0iGijd9XChPAYshVn0buKQI0LmUeN4ZWu6BQc4uxKp7f1jJO
ujL9nyoBep7Xv3Gz2IzXoOvngmJY5tt+jNY4DPAOwj3/MV2U6lOqOE34J2PA
FklKjLicVynpS0yLYT+5a3OEspQGDu4y+n/XpSpHPdjSBBldr8vJdtR6ND2z
ldKnaqzwVRJdEBN6ibmrbmoK3jWGCr/IldC5oG9Qi1in8b/LHkbHpzdZONzN
UfOKl4qk5fbGRT4+FAqmzr6B0bCylhKv9IPUybxIC0Yo0xn8pph/NNNoF8DL
U6CaltPYXsobL00bfDKJf/B+RBwupZ28KrwKA9fyQffzgc30nS9l2kVisaXh
YBrGzbl69M39/cTUUrqrSlUvoM7hNXnYWWTw50MfIq1EjqxCIezYbz1ifTOZ
eW1GvS9svzLLFMhw6b+gFxbZYfRpeeZPgXXraqkRPwwRWevFxmttbavK0r1L
Wpd/Z39HXcBeeIvEpcdwq3PXWo21ljL1b8194WAC4zBRXfSdt99BJ38GD8VQ
1iiwrjy6omYvCDCYGThp5HPcVjSp1bzcHYPQ6gYu5FDDRPeGuPkbYKkKz0cw
izcTTyLHHuW3FvY+tpZFSCAHJhRmEw5WR2xl3/FifUtCPcJiGI35lwGLfUL0
KTzOfeF+CVA9j6oBtLF7ufOXZhmbFzxNRdvuLovsMr1DmYXVRlZBxxcJ2g/0
GSE5WghKMNzBH6paOuGcDgFxLO8iHrLBS9Pm4EQCtjczX5BIhJp2+jD8I5Kh
IivhP3NgrrYeYCAJgp7iJT4wOgBeFi7RK1xdyi5lk+zbD2ofTv3M8Yu0IY8N
l0YdOHkHVxTqsllVOWu1NjcqiflWtlYA/OsSi5g9WoUEcjWYw8x2wvBBdKPF
JfFM7zrCWPc7cUtv8FbLyNZjenhTADEFjmjhcPWiZexznDzewWEUYv/i4P6a
JiTyK3aNNIC79C7vRVmrfsZBDoh0zxMJ3oHSBKdKZOCsn32hlhUnHpflAydY
4E/N2uatFB07HscM8TrxeNVIpcGSVQ9sR9JpJwpwIVS5SzUc2J8zOM+kCjFb
QpOwKiEtucfjs8a8NQFlXMfJUH4x3Xu9//PfD4334TnejUio8x64y/Knn7A3
77lUbhX3aoA2gvdZBhlVAcjp6wTDw6/eZxTuSTIrJRBuplUlW3HQTBGVDfVm
Nyldmu7vL9c6WAQpuyiTizDVvmAr631hIu5qKUiOOyAaRHK8aVVDTWcdqHuW
fqPsUYMFbFIzOVg1lkys9kAoiu9ybERA4HhNYl7oTyNp2rav2aLWLeC/tDrL
/Q+L8cQ4P+bHIeat4kS5hofZTq8NrGWy6s3sAWsms8cT9rHO7uUk7AIyzlRk
Vw433RCdDJRSM3Q0HkEF5rHsNmw5jacxKNO9iv2+VVMBG+XJiHGQR4x66sxK
Knm5T9q4oAjKUjWogcVlT8VJlOZ7YW46Rwaorn5ZbmdnVSpEoem7lq4uLrS1
vmle+GZ7RxV8NTuCad4f51rVsMqY5uv38z5l7IeYuc4w80YOXxQsnDeu9GKB
3i/NemRU6cD66hfxJuzZN6JgpXNL1VNbeFIjx7cOwAjbjammOtqGcWXRaWdh
iw4t+o98HJ6vNLB1pk14sJMRvGbLwwt9COj7UJGPZ8p2lrvPziZMO7GJojDt
LoE/LuTIn//6zu7hlw0KY2q0QoUNkRNCTCNaDSMzlKbouE6nEU1RHArNO3Ez
r2hyWsdpY1IL8t0gmCXXwf4kU2xav9rddbs6RptR13TytcknOLeLteinEVfe
PfiMFH9Rv7N9u1kTz5+EnlAyyGq2KLpaEt4L3EWS8zPzDRrqOCu/YGdXrjsJ
xL+zerpYBZ7jGm6Vnn0bFwLtqKmyq7NIyiWxILNHtbrzOkdUv9iqm+5Pm8CJ
cuVpvE6CvASbVORTTA3quEaNiOR3wYlZEUZjAGV9xGHDsDaDtLpGdBrphDuR
lhob3Bowrg/jMVePexEyctT0WcexqUMamExlUZgLvtlo38EzvFjLCDrgm+BA
X79v2octg0Lz+flO8ZzbXNXFA0II1iC4TMV66+d+YRLayL7EMM89jKg/x5wV
CMuaCy5HWE75ymGlKGI88/Ycuf9k/GahWRTqoi2Xy8F+RJGtmqjuvbvasKGm
tS0XOOJZiskW//mDuMebLjdt1SRkpwjJrPhgnllodhZTyvBbo9nZYTfu+U1m
mPsv4/qsFZhniZaSdY3MCkPhcZjJEbcB0aLl9wfUbbtCk6inIYJUcm42Ec3F
gmBItr8qbuZHqazxAKSToExPnKM9uAoI8jYrvCw7Zwccf+RIgyZWxrMkEo/y
stv+/0ALMbz0oyBKwnT5pICagC+/KZ2FnDJ7UZNlq3fL8Hez11Hn6ykpfPWw
iUDxhxpPkeX9ubQJkaFv4LDL8YZP7h3UwRAy+jj/FFvPyzCYxTs3YR2RbOcW
9dNM4HP5j99XObpPGBzPiErsuIS/RxIuSTbVozLuE0GGbNKBj//SzpiVJANk
ENkAfY66CJ5fUW2xxHiNwCn7U5sRjL/PyGitkCGI6faF8Les5+otiBN7YoY3
dFvCwUyykvR7YmKetTLehwUD8/TkGNMzet1FOwGtGS6XHhPQtaSmGCnyRseX
Do8KJmAtykVMkZgT2n/Z+qpw4LYs5zejXvg+r+czJh6+1IMu22qLnZ0YlKT9
b7Qzn2a+5ACLyhAEJnoN1JQHOFwuJYoAj+uWe8oXfUwYjwvMN/MUshxiXDHL
FeRoYjFGixJnrALdHhMzhkNzE1VMp5B1PA+erwOJvWZYThoobevQYF+MVujs
JToAy0V6sjcJdMUn0gRFKFqrhlQwPuin6cJV0hVrifpfigVlZvQeD+x+XLsj
s/nBmtNOzg4UpOTEVcTJiONxmBvgYAfVsJfp71Aa2JDMN/ggnFiHasmyMr08
BX9wDFt4muNbOz4e4DTqi5XLlBHXwEhDOxlvx/BNrRhnAxiZevmxxb6geUD8
j1ISVSX45DVhq9ftLycFKd1vBg4wstWLkVqUQ6QFRd4kLoiaR7l1kBRC0lAq
MOSB2N2u3xgSroU0O5uP+jXS0GGTgE27kWtAbi/+BL69Kqvs0gdFxfokBfLr
XTtpYAYoExBfpFiMUIbCT9WwaSM+YIr8ERufup8+h6LHtRUdOkYZzZjzYFaG
ijdPtMyBbHx3S+r2BWSNmN6Sbsh0AP/FtBRB8nLCZwjdVIQGVVC4C7WR3GIx
wPl5oExxUoYWRmkefE6Mm3jaMkPEFgw1wchuQZxqkhmwr4zgQCTyxW/22+Nh
oHM0C99DpvT2NJYcETOa7495dZKvlwErohYfPpaQMf6muX6EedvQ5tShecAg
vke2W2xblFsio0ixES+TwbgWiTce6FpV1R31M++8TR/vJzXkPn8vWohrhuBd
AtBFwLk4hc4c7gSjT/zmvo5anFJxlIyjHMb9aOaral2AxgPgWzXHWhnRM6N+
FhBi+8EoJ7GDphgqYKe7+y4TkF+qRsZKeGX2XPTRZz3XdkVeoskRAzDJHA9t
W6SQfcTFDj+XCCuB43DzpgwMjbm0iGd6nCGq69bcJqx1MdORnrAES+1ifa18
Xn7+QOSx2QR0QU8ilyt1Y3kK1wT6Xndepc2wrrFAuEtu1qOKHdHYE1LlJyhv
+DJxnxuUtU05K72NS28FyKInNDMyCDlU0mpKuCV8oIZezjkJRsOf25mJ/8ep
go5PcXFt4OXzbUequjv9W14FaMqciBLJYWktjz4cSI2rbHPiYIx5hgcDxMJC
Le0e2lypLxF+5oRBrMXIdEM+G6BK0NIvUMeKYyrhUKXosQOyyWcYMDH5Ef25
hSHzMMzAUZ4bfAlAUO5+iFYUm6Zd+zfqlMQE5oZiG7nxYCJ+QJGwxH9tAnMt
ECNftWnVGIT3pZGMbD0lpjTLnPoEGLEbsbqW/f37OulPNC4ybA3CEAXeDSmc
1fcGccdUBQEG5iPtHv7yIOlvsKjM2oXAvKkIVsTRKzyDU5OR0dmjkKy0mic9
oisDKeIQsZKajYSEMA2tji6Wy/gP6Zhzj6vAWhXTL0yxsA58g8arjtLf1Edu
RvgOEhT24qi9eQMgMoyEExd6jdz1YTFEcAf+DheRcINguOaqLKRV6w73ULem
gXZROcwAa7pPE7iflZcZPVjagnMtpiTwltG8/PPGPZ7EvlGilZH5Emm/OWmC
QxpCEtwsUIBRJMccvtCb5KwF4Nqw/6Uh0HAN0tfeVKHTSfirZ6ka1TB/TOKz
PkIagvVUfnSTABivS1Gwi+UVrmk5lBm+pd9m3jqgU5ILVMaQYOg8JLtXcqhD
GioI/zXkMdCWYpeTsHFUiPPYGs0rB4SkFxys5xk34aKb6QVhBV6Sxv1Vva27
Z13lbchmQGWMiDYGvzLWwqza/x/u0/EfF2gLdog/fcNmUZ0NIGoOhgrt7kfo
mjv1XPJo318lLKA+b1zjVaNQXE9bAcONDhe75oSTSXez7CJb2glJSXSTfwfg
y05IpHCTJihYqH8CL1L55fKCIE8RLi68tzIO908FE4GZ9DqvT9RWvLspJvN7
YMYGvltFAoP11E32/QQOn3sYVUJUUtx/AhPQOW/L6m7W3LmEMwGLAvcCJ3Ry
otye8Nrxau3WDjPV43Xr46Y6Es9VR0pxL7hwX40guxipZ3+yjD+fAF9W1TxK
sGnpmeuCJaiioixSgBFjit9f0d0M8AArmd9qNc2ffgaK8Y5DSP/Jwhqsd5n7
E/8a9D4JL0EzFTutzNAShvmR7HPEPPls/nTTXP3Ll8/e0w+H7d8YJP5uhqlu
JCzx95Cx5OkAgMa1zT0kNTMHC7i9ANmVTrzLPRi5IKmAOK5wE3IM8VIGUfuT
E9gZxOGpeHYDYr3wVtNDpD9xGEXrzdnstTPAzDjT6hpy/D3LXLBjnxM800W7
7o3NSmfg01qUBurAvHcD5r+7XR3UDCObdD2uxG1hOu2AJ6EIEuVZ3hpFRI1m
+sHgxtiGYkZahVf2O5YuRtVpw2wDj8CqmHMxwyjewQI/5qcBGSdI/cawYutp
cWCSPHT2J+h6+/lOFXx4g0/Y29oRdNog8VRnwPDgjVOrmZ2owejmDM1JJdJO
OIp5DwtOf27xCrIBQcXqSu1z0caKMpaoBm/RXp47sqnLf7l1E2futXdPqyls
JihfKqfGBEAWitS3ZLBke6V+CWhV1GAawTJ2taEPuVMrYZkliroBuzqwL00F
guKZQFJK6nFyxxYp3DqkXH7D+UXbhyehhoSP4n4AsuDonBVZ7onvnvp0T201
gaDufvPjMCy/iJmxDk7IIAnDda1I1Us7Cd8W0bB1YuqZRsg1kKowzjBpDw/S
VwhXtKiR26G5ZK/vFb0ouTZUKvTB1D4N1vcdhB6Zfqplppjiw0FmOXLxsxDo
9e1InEeNpRDwcLblwDtPPUi2/8KzBLpwWqmTwJlpIcbM9nBj9ccYjf7HWdm5
C4Zv0OvFHN3P8U7gcVaiRTO7aPBTn4HdmySFbLF+06QUMn5lUiBzQqXy9ejY
0lYaoICVgSY4lBLhlanHlySgZHVBG4kUdXy3G12Mg1PEiHGjKzNQrgu2NryO
HnEHcPRgqYLWx2Z1a4oTOdx9RI1rK1WyzBhWXsX+RWdyohKJYvYw5UBzCNya
G+Fui74K0zU1R0ALV9FDyzdyzWz7ySWuR/3B+Egp5UKyyqv/LkIJPukUkQGm
MuPuY4Nh/BZ2PzFOXym5j4tDzWziiyJna/4zqmSbJHC/TInwsjTFiY9L2EMZ
bi1V3HkcsBy9dQn0AO+4nRzvlS327j59aI4/Nte0LZsLoIRFGZcLVZMBqsSB
Q4OBSq9dPQQJUARVJqlnmMNHjYNjaq4iTwAH6uKzb3b7DVY2tzdC8oOPFEc+
LRTETUhCf5+tLUxhkVVdWNCird7f/WVyxn+gkyjGXtXBh9zXvn2IHr82NIge
i6v5onBKAWVSZU+Vj5T6OJzxmODa4nnaqWCVNuGCKThC/SRh/wI9quDlUeJM
yWgV+xDW2PqbSUnRL8p3CR/1B9IGJpHgw8OkYZHhbnwZIk9y3eEn3RMpd1np
Ap1lE6mHfPg+FKbPlciYAXESMVM5mUGbo1oGIqnnYA1cO91hwgHteOAb+DgN
iHyLSFPsNFKCsRtLPSBHrLLengROhGDTzly47GEM4qz6R9Zn2lW3wLjBBZqx
OC5ILoq4MGcws+FYz90zfR9PXVMdEEsUaI4WZ/iX2ON3rMu+B2C0ZyKIOqup
++NInlA7GDJ1L+0EF2P7srwhfruDWI+TBWRU7hg2R8gFYrAU0KW61DdlrXK+
YmK0eBI3RND9Cco422tLi23lfIgEiE5XSS+cPOFxxgyzJpHGBak2DeTsoJhX
7iKVgDgLgLzzSNTsgr6Y1xiDjczGwlAfNnGcNJq8rZDHYDW125wnE20SRDmm
n/luFdB9wV78358L0y99OsPcfSusPFzpHxSbGs6vi7vjAJwD+Uao60+xd9Uy
C5vbDxUtxEXfeKunhZ3lqUhOGds5ia3G6mJOHSJ/fMvxFSA7gxWBoLwjKljT
8iRY1mUxVwIiKgTc3jImt5beOW29VR7wk5MXa1720rOgU3BSZdJvdregpfkJ
UAwuH6CheoskrXqPhrDk4i7WRFLH25UMIBXeZsaiHhwvjTZrFFs+Q8/krAIt
ASVkve91IR58NgP9FKEgNln/+Ab/axuLGhGB+H3cPVuDkay14Db3uvC7NOJX
L7R/y1mhYPbNmWj872IGRAUt2Pbfs8bREr6aOPADqpnOXqxb1ZHbyDKewLy2
FkYHRwbHHyj2cTBaf/lTkBdb9tK2ZNwh147nbBvc/R6M2y3OJm1V1Qb7Pdl7
GUJPu5eISJ6txfB8P4Gj0T+qdf6c3K4Ma+dQgVuHTGOgS6RN3bwsCiZi+PjZ
dumExBvLvhWameTtc62IWT64i2yTU6uisH1h/KzHrZvKGPhGXT8BOjd68MAz
KkjpeuRkPKFg1OAZquaLQfMlRzvY0blnPDkFzgzMRTcRyi1TVk7M9pV0B/rW
kI7fmLQikFgAnyuVCSBZp1qylLDXzgjE7yZ1+C4ZymYsD7dSbN0X8hNZpAIC
aXvsQBy67x0IvKTOArkyuIZfQVHU0ea9kqPs3+LaZs/SkoQhz7/Ole9M8aeq
NLigVIHS20bKUhIX3okXGzkKEFnQPuq0G6tZ6uOqiCutE94jyWZ1osPRT+VX
GpXSGcLdgaH8YI3QNEm4S05OwcHfoAjbsPa9Iz8ihlkS4cSzJdPwhFR1ZItS
guNovDJQLgzitWR2hXPL1X1Nv2Zwy0qhes+bbQ5bkDVU7boNKkmOsxnSYOUs
5QoB8fIZ4gPLIbF0Qg48ej8N4RlX0R2LICU+l76IDdJHRf2pkuApVPHMHODe
OBXBvqys2h94BjMdWpxfugVbAmAFI+gvsdpXQTH3jD8Ntkch32+6m/r6Xkaj
eS4vl+6XBHjINtl9vdN7MjO9uuhlFh3nHLCxZK3vI3ynk53GsAD1QsfCt+iW
bxtByYaaPMunXjVzCDVsue/KPKTiGmuDw9VSfvh1V34/hbeH235rxBdx9bB3
EeN4xwKbv0LcT/zuWWX8x5JYKiXodRkwrx4qRGnX8mcVKpCLsaSieEMRpzSn
+3hWPcNxJJVmQpp1YQC9cbcediJvqgpdPZ3XHfN+KXs/7AYIm4OH6O/6zkai
pLq4nkeqHT1rW7KETuRlgEszInDZ4y2C9YAY9EEoXZ2umeFHCvFjJzd+oXgk
aDj/565AF7gNY2b+TmYrvf6EBK4o70RSkS+Xr/yXlBjdU+ygOLIObEcHcgFx
uLBfncn2tOiLScGD+leFVlr9kaVK6TZYGRUQxcj4NnQm6euOK39CDkdEdsZr
/zhsNTWAX3NOStTQhTGP/jSvl7G24rqfevxAw43c99vcp3O8pjDrlWgXIVUk
VfZP1pG2hlH9/mZ1IIvPpq38BL0TxesOqKUUl1Q63lnUtD36ESzUJxOepFUO
3ji4Q+0wEGQymrVE5+vsJEAGEy1xarwSl50RYF8xTH2Z0xbxVrSUnNQb2XH5
jtnBWaADV1OTa9FVgiJ5Mf/IlKRh5R1HTOv84Pm4eiaVfJM9a4z8+meGdCYp
feQXiGUfxUp81hHow5xiGfdhmdGcYw4xJk6SsPjDIqUqliU7bT+KoXp9aqRU
YO9feVfoujOwPfW209NM9VwQ8exJ/9lbgxpxhKJ7ybrcfw939Gq+JtjQkPxV
Y1BUXUSAQ7dhxLxxxZDLVMUakeuZUU5xCjUw5OGqO72UD5v81WzrMBT2lbdW
VGsQvdJc3sW4Pdp40VBUh8ms2/6/E7QrpcUnub43L6tdBo2fVH15dMLCt7HH
8UyEFRpxkYbVL5bgYF3o9+ae0M9ir+E1yz4nwcXrC04WVpn5qXUU84OUg1Ym
8W1CowXJNxL3Axc3pQPYo8cK9Jk6EiuHdqBou0abvcdbvdyPiMP6BdqzgI6U
Ou0BAuxGMCWlFRONCpal+B3Ji2ApPwp/C/rLirOD/NLf2LpbIIxAX84zWMoO
NXeVgJ1MvNSDw7/cXJvaoWmEqlIP69FkFpjRS6HyZOPlbWnGNcMvc+l9pv/U
EcxoSVQAAWLRIfY2kBc58vDLpuPkE5CKdZunaU5TLN4JooZK9dqMOvOOS8Nj
0fLVjSFq/G0f53Hr2hDT4lMkb6gyDbyFFIDxH1oL/w0tfdhMFloE5EMIbJrU
eHOfjosOiOnL2LbVNx4IK0FDWXUfbsQRuW8mnokU5aIRiN6ceQh2nv99zgDj
f5DgJ8puYPp20VHhU5j4bMZ7j+FSJgWTAKNFOWz3agPk/+5m5pk+BTm7DyRq
9FrCQIWsIYlzl/nFlFsU352rjoxFcFDj7KiMjwKFU5zOMMpbjwQ4lOwSOcVK
cWHElE1qPDPA4y/3KzlBMi6+i60zvoxNdYm32pbGu77VAw2BDDb8Eu7fc7VD
EPlUL1IfHm3IMq6tUs26NODKJ7d0UOvR1XdjBePG7PpuwB1f1sjPHXMsl+6+
ftOXYPFI2TGwhOyE9dU+Uop/JZX7XDCO5qEcL/mnvgzjbCs7N+4SRl9Sez1Z
oA08rI9U1N69HqWvIYRzD+BKvxuoM12uSgP6NOX3PplG2b+sv9PoYC53b39O
6eir3ITRBfKbj4e/m1Y5RL5uzezlKNB8m3hTdR891e+7DqMrd8l8u37FwBFz
KgKEsfN79i/JhDwqlB7giXGei8pligm53zPCRVt6ORs47J1zyjW6vZCz8ZjK
JYrSbdKh/qNfJxNPS9tBTcjWJ2+CYFHn307jSAAES5MTMg5dy8vtoz6HDFjW
rrlIDG6NC42dtlc62WdBOSK0w1PE5O9yZbD2f9A1+rIca2KESrjG5QB/KPP0
JjTJruPUYBK7CePZ7WlBqWDcLKkBE2m5Nqas+xQ75Da3qUfg6foPv2paClQm
qWYidzJKm7bgvg59BwB10FlbzEyYcwz4Lmx98/CdEC2uL2WFe66dwPO7H+lm
bLMkMjnxWHeSZL02Ij2+Wxx8WPLfJSqoLWDFb7KFj7RpX0l6kQ0C1dFKqtXt
sCoJWn0IrqO9VyKbAeez4QQHMuhsVv4+gfXN4pfjPx887VkadBiGGLqfd76f
vrvr1MgU31YUqt7BOf718054hS9CwXFydSJddGVFlHS1fx6vhW2mmW0wmin/
6E1BcncOvf5+uuH2HdPL+BV00Mc3WngpBHcuijL24zVY49nX6+xGEIYzJHA5
dN6WIuRj87t6jvsDKYbrsjSSa/4Y4q0HNyuQLubmw8mr6qCfpDGqTQVvrhm7
ksAgR0dRnmE9OjVYoh6JcjjQ36vdsOxTZkzTmPH/DCNftwhQKwCf/gY4uno7
L2cPnxZdywlt/S3Ci6t+ODWJiEMtpR320DvvnM7RmFK3i2SglP/amKn0t6HQ
pMQT4L5FsuPYbyF17OP0ftiekiPbSErzZtVmEHn8XcAfUxrhEuk3fPUa5goO
wweitqpKK/BiMXR3KqjtPeyb/1LKVw6tbvvAZiOUyVcaD7pLQ8Uetbp1fr4T
T0WD3FI4tk/gtLF1Xk6+pDoRNd4mmtMwJV3pympYvpWAkjFgq68XycrcrDqP
smScICctyadCVEWp9LWGev3IFzYzaI4+A23FOel9Bo3+uLBarCKGLx+opv+i
Ha3OpcuBE+x4MyKoEsB/eL7sfQVRUnL0g65OsnNeZvPMRft+oJpiF2EdOOyn
H/7kgtnwmtNVSpWS+peDF3vmzU0eR+7uIPSFjR3cOfWJY6uBaoVFiEFAcmVC
X2iFiP5hdEK7+Rif7om0d5FGZIVvZY92ctO49e+p5m+79pUygtSzp0Dbpbm0
KQkcCiKZfCSYbWDgJjjDJVujtxDw5vFOsveftZNTiH+CuO4Ra/zLBCecWKFj
B93+ajfx7SsOliReRF0N5RPft98TP5AgLoiiD1v+PvA1Jw7BO5PAa7ALobfy
z0JOyJmU5rg+M5paBwsoMx5tLOYSBKAidU5eYDG03KSJqYwaU/QOMIZowunv
V7BE/wsAUlj7j7IgDNDyLiX9cTcg1oxY0zl6VIC9mJGeXH8LzPJXmhfycI29
ViNq5jeXoGiudfqCWOoft8nLxQ8s9Kv2QActzcqrKaJ4eytiuIF22L9jvvWV
0zGdvraLdZ7UHgTOvJ0440vPrEOj2WYgTGIsOMwM4suRK7NVDEnxuPm1Fzhn
sy9tuK996nYLMxK9WTDTcTJDQAR52YlYsMxq7QEr8IjEbM5QBf0NifwCoccR
KUZYASaFkUBxgC8gbJX0FtmFZ+QvJJ8SEk5dHGYYz28W/wHiBRIlpXDLbaOn
9tbo2c4GxLbRSCA7RY/Zi/oUg1v8LMgf+JrK2wvhZkQh6twcpwCpPHwrUA1X
g72DuCx75tVQ2DR6EVmWcJgve2pxLrTQxd8oCcFoQw06BdWFKO9XABfte66A
e4A6QlsJpcX9sa7Rv5pjgiqe0FMwtX23tjhXxhDJ63V5jH9XbnsKpHoF05IG
zNDcZhoxrJPO0qXvB5LLkF31qgQdNhTiS9DWxX7ZkD6dKaI2GjeENNaSH6UL
vVp7PajMX2L3L8wkVwMBMpHeJV6QOOhrNadjsjSjaTpMhXf6XdKHgtOY7rxP
/p/mu2fWqsD6UMhH40OFE8vLz+v5QisLlVjbUiGaqaFOUwDmJj/8BTrwqD/V
scVoF09CmVXlm5Jl2FKal4sdIdFSwj3+HtelB16UaxZcuFdSMZK3iEC+ywrp
s6uuZkomUNq3zNKj56he9seCCHBKdeeCpqNlKxXWxBWktfNybpaIg1nrQRgM
LxfVobmPK16WYRIw+UWwaj1xDRaLVZ2zkwGYvo1kI3YOy7lzaZB+n3LvADl4
nzwWOzjAYJoQIAlINH01YDBCyKAYFEAm8FUZM8TCqxL6xXINo4GEM09kM3uR
kD3IHRD2BnrYwfAqrwpQ/Slqb7RsE3G9LmuHwUD4SScIQQXl+A9q0R1/g+hr
i02opr6Lo0AM+flI2GtUVYx1SH4DkCrY7owmTcqo7HpiGnhCzKMxTHK8fuxE
4TzCsuc6XtnsyKrtO67cS1wCsaGIbrR9WiAauDL/KcZ8jk5Da4ZQrLjmb/mH
PNlgjI5JrdqF/SxMKgezxg5bjEXYTOW280a2DZ3UMUROG9+dLsTe+Qba4Gn/
vMDhvICF5FomN0jhn31MdeaGppzkuTWUC5GW756c8Afur4jCLWtiXqkShSbG
9b+vTveM7CmS3k96M+64BnKqtCzdYjhAVThnTBi6KXwGOqhOJVr2dOS76mSp
b85o3a0NNZJmQp5qWLU+kQoi5QqqS8jeoqEeqzB5SC/5MBig0u2V0qxj09ef
3+fNFOoXkm3HNu4bQCTr50QgFwTVnzbmBePlL3EIZWaomeCnMkytLTrQpKLx
E2MbqVCijChvpMDHgSKPYfSUmsChHLUax8SV4pkdQlgQEYjIoNEt86+qadUm
fe23FgMT2RRgE07fdow2w153LBXRxP1OyXG7S1FRsuuwc1juNvklbie5pFGh
QRY84766ZxlfOKBCGdVMsboCVhbPJwZaaIOT2ILxNKBCsV6igdE8iLyo3Xrp
gOBGmk+S8VjckuZNvITWEcWMw3tvsu3mIYgGmkVqnkSAB7f1octZ841UDKxg
Kgpytq6Ze47RsAebMfKduw5nUGB0yTW/S5NUrwWh8118bHJq8rvBYSGq+Jsx
TaLm6Qq6lHWolY9GDkPWrjod+X2X46PN7wXDzEhROP7DTJT9+A7ovpjMBX6a
YoLt0Zg+LzSIq+DJ5jTOoXlbJyN1TfOnlXCfkgUJ9C6VHNG5C1Ow7hr7iAr5
DYAsQH18OTR5K5PeLTT6NEQfGQOn6/asdneO4iT3obuM8oKPfEmApFStYoqL
m/3Z4wNcKwnFQMiU+UzBXXEcz5SQlrAgIPTM0zgm7NGFN4nz7w1uyl4ZUt7s
CdliNXJI30is+hJf/zN0AuMczR8fq+7O8du34s1zjqacSsBm2uLcB5CE4a4n
E7sOUg3pKjbJXM1zs2HjFKLwEl1Zv02aCd/ePvH5EiPz7w8TD0SAypk1P02/
tAN4MqXLZlAegg0H8ANeHKSMjX05QebL1QiNQA+7wYMCOmffEoZoeaqBCz9h
Lrt4WcFRYkIQwEjy2AOAhP/yX7BJEWohbiNlY8eeBLdOUDm5nUrcJAzAADwX
3MTQWNbv/wd4T3xT68uDFJ5rHazFAOltN0O/vP7r1Dku8NAOLb4+O1fDwPJZ
J8gkbcobwKcO2mFU9xj8glmWDZZ3BOJFrxmJvgLkgLOoQUCgElfYKbve2jLS
nY4Jmgjm1r0ZbgJGVdEfw5Cf3WLD+pbKG6z3AkHrd9CqxaNs8GsdD9P+kO7H
WpmuRUcROuwooMm5SRKWRw3E4H7C68Vj+lw41gMyUWJsWKU07LBgFvhsRJds
zN2l9AxvS73Cct/9xkZj9WCv9DcJ81onB8C5BJ2sfiudNezIHv12Qiz8x3V/
YN8lWknMpSA9DqRi4GJCpXB9dnOMqFIJCyaXwRyjeVI9M87wFSr2+SLPO6Xa
vbGngQDtRQ1HlSKA6tCRjL/X+RdjdEFVz3rjjdB5/jmkE19CDujP/oajrAQv
yzuT2wseQVFSbIZTQB+hqtQ7J1Na/miAP9hszchPzCoyiY/ZGPjEfee4OAQ2
c7qu+//oo/dWwEQctDAS4JHka58UU2wkr9UDSuEdmBkqwi6vI/RRptMVKX3f
2nv09cvKQMvXFqE90IPD4Nj1q2NnfiA3qMRcBLAKlmEjCkcyfqghfAi2dViH
jzcKU/EM0bv3KI+GvzgfXV0OLzXGgn6wE+Kvyq32TtJO3AOgGxn/TxI7UnQp
SwUqjeU3kym1/v7blTYYdTRsRBYRJm+LViNtsUFR+zV4nDg5wAzXPHDqCqfJ
yWsHYK5Atk6Apf4n1OuTF77kv6wYqH10lvEeOVezahgdPa584WWGewZt8IfN
4LyqpC3Shkf4p4Sw5YztEkNjhe1v3rRzNS+kSBVZ7Zp9ai2w6uiLx4jWqqWg
8bFBVlD46iBMWrDuxeAjITC9MMon4MKh8LTe9XAHcGe1FQbGvhGum1y2UhrF
pdlYWLze+UGo1lgmgKqyMTJ4Y0L04HgqmFeFqJXkqqV//o88jltcWjvEuVNY
Ij4o5Kyh1mhZcB5qLcKME6DAOVAHkLBb8/YCBtvU9YCYZZlR0Y6l26saBg9Z
/o/nGwf3sNIv1K2qaLLBXh7F2FZHhTwhLvGD+j9xG6IQ1iKmksWxX6+ozQi+
jlUGO/ucaA45T78QDP8e3kCxd0ebI7OQxXyJNYHoT5s8C45RciQC1mhivwnF
xE+lzpthTvmpjUk8eEWq17u7eDjUrAiG8c47CuCiVb0WuQNRqQ+4QkNzz2Dn
LaWwuI4Ag33VrZHSCCaiVsFlQGRkA6dp/yCIu6SN2NEHBkrrqsA/PYOlDwI5
5+43QGcxUA+j2+AqL8N6jBKprpxPVrynDFe0CYeT58S339qlFcVgXtiQJHMK
/YsIGfvAN7SdVEI+Yil2Dv5zX12bjDt0izzyfzKrUKrgy4470VtN4mdEM/o7
nzADKCta8iym64eoMkyRSGVZG1KuiUi++qwl0y2PV0IVLG74+PeA+aM7TKEI
sV+ERaz0A6SobZlgwkOzmItKM5wMXp4PuqlDux6V0HpQaiA6JtGPyi1RLmcG
Uta4sb2sHkjJHYe/IAqo8d951o/45Z/T7xAQlNaivMIK75yMZTWOdRsc2e5l
wNq2Kt1zM81Dpry5bXTKresIdma0vTU3l/UWd64olL0L/UTgCwsOWfQgUV2s
VpY8vD8xwbM54XgHxv5v9rsKyCHJgfOziq21bLwMpWcHmKygSMRYyCBegPR0
GMJdykXcaAV/Ljpa1HPJQ+4+MVSAzGxooz4wfP//XmrkZqGCdQPPwhTfyFPx
Utf1BKcJ9gVNrlvIrOJYaWzjLlHWjHzJ1CETD97HWX+aMeorajo5gISb+zyX
JwBSB73j8m8fHtW00cw11sPtOzUFYfrJ8PRxxKdIXAjGCSBSzYcSUtLz8uSR
l/8kUuidzr8uyp9y4tRdj/e2tKzllJD8mb1zWyhGvZGeh2PynLpsxtOkcUer
j3HofoSfknUxIaziFeSqWDX/lVdlZt/VwY3yWfLywcqMD00/VsMr9rvW/5U2
uO4RaTqbYlXP07xTdQZhWXYcY0o9t3WR042QJRTYyku0jEpmX4bHuYbLefJl
ziL78/Lq0mFKwTxw2O6tlW+CneVI1MOY/PaGraQOBcdJx2BN7HF0/svIv5ks
Tl1U1Wz9zsEqEDR2JqY36UTcWLOAsGW1W+Y1kheu6eyDmJcLWd8bnnlKyy2F
zvqpChxopFqqqmvcoGXG5DiUxt1zobpBhH1JrqRz59b18ufVPBeDWlm6M7ef
K3sEMYoo6f3rF+jKAy1SbXmVoHG61UEso60uQoRL4s5loqqqeciYR5EyfqKe
8dJEfUDV67p/gqLseN0Ib5sIzd9J67hV4gevBjZ3gCF0JT1Q3mZNzf4Uix8t
IV2lnUVyYWxxstDMRniXSgSEDZJl0ot18txN36a1xrCJHeNHN25WjteDuKuo
fLOu/Y/f/yCn2h21Rkf1WE2i/m+2VoCNVVR1IxUsGOGtLPjcvM0g1RJJaI5U
cG6BJxo52z0RnIqTghAQXNABLRGAG7vQtvSP6VIE12Ogi/iqWLNrTI3H8r05
UXmejAMh089O6KoCxAu33EwJUElPKO0SZE51PXJd6aNRsJtB3RlD6t63nGIJ
EHyFRzL/BrT/jI56KQ5qhEkRTwhSKZAcZbaHvrY6Qb6TwSKj7dcgMR6X9x9H
6GDl8LfBC++TfiZPRcRyB38fvchRfLmvzZM9Zr6YBQIggSVjzmBDi33d3j1b
XeFCNL1imCK2sotpQS12GiW/dvFtoxDSFzc1x1T4jAwCrqmvoVLLhocNSzo+
Y3Na50CclziXMDRaVYtTZde+Vu1wjdUNMPAXFVnyu24XpSO3xo0BKczje6hg
fmJBJMe86fV+lK/Vmu07KPM9kEg9XXJCRoUZoVRjiIpU+AXY716DB1EFegRG
jcFmW48wNX/HlbpXgXFGz9JI3/LVcxeTTCrq7mNHm5AxvlSuXJcQpiAxQgyI
iM/xR6RH5wdFqJeUSWn/GTyRf63gSOzFX3Mcs/mFvm2epoJC8M2LaAMfBp5d
XE5TEwNxaWu/PrFJJ6gXeIAwY6Dm5opU8uyp2qTUM6fea3woHxa3UWs6FZqa
VeRKWJSFbOhTl6Q742BqRaHFAmZJkXb4Rp8dUvvAcXjuZFr0bJ5WaSlRyvQp
JlZWX1jfI8zneX3rHkEBnZHd7AmANgm8F0vByQRSiAfuTb9wet4cS4k1Vbke
tdPjEQy0Slk+VVuMnqVoxHTWykjfMm+ey87pPZXvWCEEKmItXW3wVmoT9Ii2
Z1G5kF8kXcF7NB5oY7LlNavhHMH7yTot4YnV+l1br+yYFsyljHhDQObMhEEk
nM060ZUR9OJX69+gBnAs0l3XtoFCR/L0io+HSuuYU0zX6JBk/h239Y+ma3aN
MJGFKKMU341x6SRLPaL+3lFDFSVSAaNktR2PvJRvpe54hi0GAMORr/QSVqUI
zOk/yujbWp75afWjH4DXa8VGY5fxKR4D/6QkBYuSS/k7T89PFPy9YvEOEJrr
Cjhh6HvEfzwHkuNfeZbjVJITWMzPT2wmTcu6FW5TfZiQPMWfOUba5M1UMzYg
PomSLyT4dr9yAubjvEyXQjLWZ2oCgEoRaTXBJnj9pIPWoqI4DKZ5I4DlYVE2
1oIL44Nxr4BL0yElUWVOzshbmMs9oQlrxlxfpz7a/J+wzhB4rb2pytaNkDt9
VnwWjJNytWeosmgKez9U6InaOHNDWH9std91Er5rK7M7142mZFwZGBdHID0e
fL8pq0AkvlijRTuKgFb1cmBpV16JrO1W0TljTLlWXFQkwzzedhUaxBrIYrpq
L+ESCVl89bLuFKrC2x2bjDf0KiVJXeYC0BycGvUpohJprhLlH13X0CGNUsZ7
KS4aiK/MXT9U7gAZQuDhl3GH1C0KvpQ8d7t9DXDvYf5N1dSdWFsyXcmacpBB
lONA3Mxt0RH1wyGw3aLY40pQTV3MJPxoNjluc5ubWo4pJCydLpMz93Lai1yN
BC2be5LwJLnASRNNHn2NFKzPdl2zz/dekCGE++atIQl9Kg1eKZhsim4zZOVH
lVzwdA+ii8jrOhEDrimYOYjx4w6DkuP9XOjGr9CnaYQXykJN6hGP1lGUn/g0
jbWwin2sN8AnIg0213St6RSs/BLnE77ByAgPIQLOpmlhNXZpWnEjGXq2dkYi
fIbTSj0OIVwO1nA5TSb35uJ4tgkvL2PofcA6Xr/+AgdrgAET2ptp123PVXGj
h2osXukCknNpBTwAOLdXMNuyoiUG76Iex9xbkuMv+jEiFGu4c4+TDYpWDtCN
RtXoiwthk58H/rLCugcYd00gPOpDB6DRSgQBU+HDKEfNYRxJB4DXVdva+1dY
U0go9Dyygz9wYBR59+7xnk0VYqEjx21DTIsfoUz7DNxuOYx0DgE/swz+dz/R
Ji2Ofu01MMq6t+t7VijODldk4c52yveHKCtAqxp0tB8sQYfHf8K35o8zwUdh
UPB0rO1CCRWDTqB9ERJOhmLpb2m8O5Jk02/zYcQxyUSuKim8Zqt87RUqbvta
PohcXWcmYSm603NWy9OMT4mthP41XnxiAofDQOhM7ENPL3sNXkYl+mN38l+i
xQGPoff743+sEYF0Uf5IYUVUga1eO9cFeGf5JyRuZQfATzGIy5688nouYlKy
C7BwbT2HZQGzIp7Hp4nQjHExnA8mX80saOcGdATbPaNu8JZ3vSC2nNlQavIQ
hebzoi51bXwOrnRn0X/rWE4qPCYAGyRlgBy6i7p4BxatdUfMQpyT6Z5by7Na
agjjAnGeQIMsFT8A+awxO8B1N6Y7bTKK9Dp+lu5OmKa2q0o2CT0Yw9E3zrlO
JCtIeNC6MN94DFxoyzvGlJJ+Xfc4VpPLpgWV5d4dsswC5s4rJOnS2PCPNq2Y
ol27RPfPyWfPSiClXdKzNwF7Ht5FooPoskGqm8RktxPgMeaxD/wO62UXttvf
9xCDSZUaBpgqI3uEV/IWk/SUIuC07bCxxfwESGomd0zw01/RsW+DbrbKuznh
QSM8qJYAmuojvnNfCw+jif5E297K5Adpq1twYgchfeYBPNn5FkcIapUgm/Fn
8PJpV3OhRjcJMBhUkjhix49WfoWSuLuQRVqRVZc4lAP7upWn7igtBlZpuwLa
/wC6R+JGEoCHsvpXZWPCIk2G4iI0+YCUfBCIB0Kp8e3tK/k2UlIAtz41lQpd
r7ZvAR+dtOE8FwQjqWWVRLcFykFU276meGdNAolf+AndV9ujiZ4i6OWHh4qX
T155NejUb5vSWdWtEuhNzMV7iP2BKRJ4XLyu4LY9B7za724RcgkTE3pE/tLR
lseddfjJ/SXqhxy+zfyQj8aq2l6U2jq9X2rnXBU+omcp6XYpLFNYjxW67Kkp
u5jI7ZsgAyfi0jtDszfDYG0C3ljFyO/LDnURuxgEjzMEZKffnLZOS6wRpWLS
BKO6jdxrwTdWMXL6jzVbx3GQOVwwGpm3aIIE7l//A89Kaw9NFm8i7oNfHTzS
+bbVUCEObmHxSLHIWjyG3hBRXtl3rnG7VFwG52UfVtmw+5Xv32B1lv2LH0Rh
iV7lyRH9Kh24gpbzz4diDE/DbR70MUM4B1Gkz7j7+ajaIjI/XRx6QjrT73wJ
p9x1PjH5FUvmj6arVnVEv4vPrK2kqU6Ci/+ronIIfRazwlnQhcPAhMvl7P0j
WwkjxV5KJaFVAhutMBRJCkTGnafdQwPK3YyjliYfTbsZDKgYPBBVpm+/XYkz
BkaXsSdLZLazCy/UFd7GwSlbNNxRxYIShtHmpJXYF5wpKt7QXgn4LxhPUzyq
JmM2Men4JDszVzowBiK6OstcrgT4QZ+YVIPwcWGqjq6TCNxFXqhZpcMwkAJh
Z2uWCbCG7hIEK3GldI0WvPWxRn3wx5JMg5kGd9rYZ3yZmmU22qnD/ZP4N+6b
hsO5nl7rj1OdvUOycLthObjcgioSdAXVzlMw7dW3R7QAaRckFtQQ5lVkaGqn
ddeYHH1VT1OjKEHWJbHypY8kF7CjtvluWalTd2u0U5M9vOJ5f5t4umQYm4k6
IlZ1ajL0N+uZTA0nVch9YEu1hv6z/2NqxeozxWz/wAzkaumLaJgUEdM4nfba
LSMoImCbzXJMxtoZC0U8x2zylEYggfd2Ddw3AK88p1sWJdFjjaU6vji9jLiQ
ZSM9xVcYsen+beXdSS83mZdbwjLrqiodWQHZs5n+my6UbNxnL1ydJPrKfgEH
ReqgmtLn5I+kG/B/mjvCiaS5jaM8++nO324DiVi6za8pylQk5OpZl+v8y3nF
dcEnaJqSra76yLvg3se3yz0xKp6hAxsyxVJJ2qCoWnMHXyVzdk6CcTQVP9Li
ZJ+QebtfLtA9u0zQhILlOwLqMd7dadmJb50GDSf0wkW3jKm5DOkiQiQMVZf+
bvn10AGUJ3pYrb8YnKI0oelskNGFA19SXyMcB1ZAs5qzpdadvXC79q8ewX89
7kusF4lLfsggoMtZxCTW+X4Tf/7eYCvEiM+/8ap1PWB+1eJQFpPEzvG2VGZx
6b8VOosO7OMphg9JJsQmMhl+Yi4IDjcSYfNxkwUWork9OmjiC57OaCCeEiLx
aT9y+EHRGNPVYOMG8LjXdROaLFBwA2ZBck4wFq9UVL1fAvbA2lbBYD8CM133
nZcbKP9C0g5cqaxCD5N/OJP8ggNm5jMO7vNx/OAvg+cJgJaXezKXfh8bNiSk
lK1TfWnOlMcxOr3Hl/RxHH6Dmo3vO7GinV/WDXKeyB4QKFBXBRyNB60paVoH
fSgbsufKLJ9THQ4wgtK9lu1lUibIp7inw6ALHlvRM7jVfrM80QIh128nPQSd
2gzEL34cThkhb6zVB9enaBr5R6OanoOwW7Wtii7DMhzdpKOuHDFfCJjmYEkQ
X7NCNrS2Ys5fDLi0KqKZlibCzEVKD0U7KqDEpXUwwC8DNQLC4WxFXYEE0IJq
eI2PklxSjTBGPKLZsJzTemOibTpmaHEnUqtdgM7uc4sIgxBahuolQWdP9XBF
M25jT5avyHHkhNiR5UZeEZlLLLa2KxxpNC84+ENlhe35jjKWg5hx8U9g4pT3
0a4FBFYkWzGaeeWeh7f6BO1vwKMLjTVUs8re9rU+xTkW8H8qJllOg4BwIsCI
r8FkG9qegRO1bZ6ssgxP/OUaVvf8A8e3ieqzVlqVewFj6AagMK/ylpq8rrqK
WnrSMt6x2EquX1mUpBpGH3sxZ8cyGsiqggHosG58qvXqA+S/28NXITNhe0E0
WU+91IKwm7a9Y7b4QtzAsBIEAfNuxknEfpA5/QSn2d69VyDHtyxAlcGX9Qqt
57A7taNlEczUn+M0THFAtDw3b6qbJsZ/Tt5InO0sXndhF/mnS+/4+jf6CI7o
kEcbnP3LQRwvCTRgYtdlupHlpV1pxqLgBd7LFfjXDXrn7LApJdsquHJD/Wb2
iQ6UciivopMegui18U94bvumZGIyloP8kV5LLw0bLZLPNY6rQypFnae89oX2
Na9Wy+9yBLFGqEGHdlPbOL8YLqJpe1YeREaE0G2QyL5JzOwk+69YLsbfUKRi
CbfV4CYu2Fxw2PBgqQ7H6U6iKPY91Rde5JKCQ5KC8S0eMN8Dvbv4suVtZVXt
6fmXZqef7D/Ni6HC8zP4Y5QJV5xzk1yMQYgq0YBCcXICrOhDMy6gc+49Tt5k
U/fxw7/XVkg6wsJ0tlw3Viui7snk3nyPma7uMF+PAzi16VxS8t5H5HId06Uk
JJCUZF7LCL0CxquQyJcr1fUtojoqhljEsGzfSfsTh8X4nzAoLgYYCqtr5087
pJ1xc3BI+yefZvZ1Kb8OR4G+Wn4ae/DCQIC+YyfqtogJesgaL7dEfVIG3t4U
DxFf4q5OMZjHw6gzUz4Zqqw7epOZOyeMabrI7YvJQpfvTs9/F4SvydvB/VN0
zaYjxGwsGASsvbA+ASa3iV/hs6oAoLq7r7qV0s6ydyw2bA4YBVLlr/yhkWoq
BrHuzybcWEmjpvHgTVU0wYqBpkSCWepKbKmkzongUkOWhvKwB2R8fbSqN2KL
nm+uCGvkjHxP3uirERzr8RNbX8Envh0HhzIPrrRejf2VnF2gAInTzYelh6qn
DhrzMJsUiPzpkLvOAD6OBm8WHvouhDmPJtuDwRMqNR0sWPC+km3LitNaOFqV
ECFIiEqhe+/bXX6eiCueOt0sbbPxGYhgRwhGG6GkK9XDHk5lX2Jx/QCn3UF2
HhYV7kdTUqAa/5KFB9KAgYlnEfyd2qsAxPdfDM942qHHby0SN2FRval8gMNU
7bhC6kE0PfJXcXVbBZ2nnsCUJ23qztQSl3GbU5hkVDnam8T4aZ/73E9CX2JW
XdddUA+gQ+YDosbr7C4aBHe/A3qlA+izSit2ccK88LMfWJ3tEl9PdTXc9LMO
NP0okLul9MXTB1LPSOxa8NjrEuiqBk76Hmo7rZmcVwkzPjWydOUIqX0x9XIr
e6jowB1fiNX0msppWfIEzSN4txaeStT9T4gORcsNIXlFUUlxOiMU2zL0INUg
XkejatY7vIfDNeu7qeBONTvsgc8n2ggDqkJO7kRiaT9kcD05VLdfEp6VIcKq
U9GyhV5DbSLgpwSt1fM87/W6g7w8dtTDZE0tPPz7OtVH+uunQfOw1s/3XRQ1
BxzE7FJ9ausIp1abDhhAkXPl60YlvtoPcFJJky34598q1Du/OleXGnTmJeMw
Nyb9tHG4sidy3vgwxtYtexJQsEB3eSlizylM8Du655rj1DAhTPaqUPvP2m5v
FQrlUigY7AHDpP3F/VNKpyYHZgneu8mOo/Lj+TH58io8eCs/hAAUeUv2wAUZ
wQwi8L6sk8tBSJR5q4zEZzRou+S+cXStDtxe2NEA0GaSzHABlbTxPfcXFIZT
SjknaLTQ4M7H2GnVDCgV6mRzPRXfTggrEuX0MjOvY4qu+8jO+VbRHLg3YeyV
Hb3hgeWit2mPlNSX7HSOSTOIwlm3Foh8/bzHrSsaFRnykwBYu/lMAyTqnEWa
7ETC5dokh+yEqT/bGt/S7+6ozu2P/CZ0bhoRcRyI6JA6eHAMEzlxS2z2BkD/
/c9WJ3HuNDnv2lG87KEHUmxpQeJDq/KTqENj8O/84KMvrYYSYtLSd7jAUsUH
P9dJnMm5HCqY3ozU5/xyuKI2khHPDS6duLF+m9B6MWB5BOvAjB8pV9dRSdgR
nS1KM1NEeMvaZUkEsq/63OUpGUfl0ih9jiDYG5AMvMWZpEC/uGR5aNWjMHj8
saak6PTGS6TiJBSbsjGZahKU4iPi84N3CYX8XlBCuaTl5JM3C6+NQPnJzXBJ
HL5c64gTWld/ccSJGITNVR2aXtAz5Oyvpl34yM8AW5RcNVXb0nu/S6+qrdiy
4PuUKPRfKFIy0GUw7I1MZQmsvz3g3qUI1IoqpvoNqAHppOUmO+pKb1DqVF0l
OOHziAZhQHhhaJ28POYGkWQOgoOJptmTZnqKuq9n9Ps4cZl9R6w3DNcSh6nZ
RyQz7jIxpsm/yXytJ3upoMDfIOtW4W0p8W5SOeiSoLSXbRzlRiKtfltu18dO
1gBNOV2FGEGjkMXDk8VUcs3ZMwY8l44FlnLpc2razSg0JyQlsoDFvWUONIja
umz10JulfJz1jFQlv/8VeV3tOuzFkYwwVCe3Y+hdAhIDpgm0KXPB/x3bmIrw
3ANGAO4BC8dCHIAk/t5o2ZJN1OqQH8DHpDZr5NOT2yaUfJDrgiwjx3YOinFm
2KVq4JRn1QhquUKt23d4GLG0LaZsPSxhvuKY46TkTHBag+KuRYLhCHV4GZ6H
NoC8ZZijmrenUf4fAeTZbkcKnQJsNT+0/dr5AwBIG1EFi794KPT+/jW0dyn5
ojnrppJQ8MjOlczPaTJLqq/mgOeRqqQWTjywSxSRA11I6dIOiV7Dt/JjaqLh
vTRwSwVkvIbqKdPjMwpuD/bUtKVRBmjIHHJ75SPRx1v2c5osbrtldzKx9Hfe
7YaZ+t1mnQP4P5qUmD+AD7ff9iRBFd0ZsJxkeUjj8lJ0m5VJYL/WHoOIbG1i
4RzoIvjQqYEf8gUlpC9U20p9B4KwtPb+V7sCDaQBGwYYtFYy9fqzRJHQ7ecU
OfsTf+gsl6z2uwg/iiha/Jsn9DQbLuTMOTyAcD9IVVXR6sQvmtlI3JjVGb9l
G2nqvqJKk5mi1DK3O3rz/CYufKHCqBTSqa5wb9ItGkEaXTd198E+DS5reJV0
DFSG28/yzNqzuNb3q93yD+dpigVzaYMGlOOk5vovykGW1DroM3f5klnMGzaR
c2xspZHkFUWAszK0TcwzoM9LnZEE5LgkRb7RTl8L6RFpKHh3gySBFuEzMJHT
TRvROHZhtMFuUgLyoRuhhdnepWPsx00Pwpgvv2bB6Ql7nuroALDd5mzq0eAR
lBL2NEQ1WTKoF4nwFXs8rR9dYsQHjRBdmwKPOwvNOi0DjvF7XD9q8JdCuW0V
8oKsh1deJXmaaB0J8zN8GaMMhqWncQ6UkG2jbbAUg8Z9WJDhPBFyMuKNnBs5
53wjp+TQkARxJ+fdNu8BwvrgI+MQHfIBJ+2F8bRkPVhlHWhRgrj+iOWotGAT
HkmbytZBuaDbGjI2IS/vlw3rXk7uUFn7aL8Dog6DryLMLzASxcorHErx7abn
c9pVUsPW8mgecmlLTWXSwDEPd27CCzYerKBIfqdD6x04X+l/4XTcbnIba3sb
0Uh2/V4T15IXqlucW7IVPNDt2hw7USHdSj/ls737NmpnNPaLsejnjyX1ZDl2
C16KDNqXiK+mebZ0Nzxr4Tbg/NVo/szJr5GH0epFf+ORpN2VrSK5RY2E5hVk
joZdRcL6H+t/G7YLCCLxs1mO/+d7b8v2Np3rBCr9yEsl198DvQvy4qaQGVl9
3n/JWZBvIKzd4a4gAodDU22w6zC4541e/X4lm/hb0API9yNyiaYMmE7Go/9N
qv2Yl7ATox2mnxsPRnMX9S9QxhF6ob8bG996Av55Ox4CPbRcR5zEYHV+XW3N
bVyfKYUbHGX13WLTTt+wZIQNgwbseH4aHeeqzJNAQpuW6ojNnwg5wiLY0Y8s
f6WeEM/QT/67yfPeLt0JEItsLqbdhbYq1N+B6GzActTZHXgJpdIhqlvog52x
Tf4pJtIQH6AMkbPYymDt4es9kPRSrrBrMIHhV593Ylm/F27qyJa5ub/j/HI/
cYif67dYztZyxs2FRSK4VfDiZXBhfSshCUDw93NTiiTC7VrrGSAZOOzX+GCr
OqvFTzmQZeMzz8z9adECBWg6azAnk+vF6YaQFO+AczhpXj8RJ93ZfDRlulEY
33NvvEO5Wktv93EDCSCOFWTn1EcESwYBSbi6qXwuYTXG0u9kA7fmvXkwsU4q
B+30RWoEshpJbdrh5I29Bd2jEF/0q2PLfcgr6BWTvncs/MpZEXCYsHE+/1ph
zd6SiPt/GhQ39+BoxpyzYX88EPDW6VtFW822knc63BYdXFvrD7kryliMcOUA
9iiq+oCTfcEjRVOJwiv2ohAfxz/BLK/cwfFSYStIFei0bX+zGREdxiNFPOB/
oojRze0UswCoSvlWtgs/7Mw1qH7jR7N4SRmazNY/eDUU2w1BIYcwl+9DPnIl
EhcGAH8klU4ggHFQxcn0aakQmr21i3uEPmT8kpn5NYnDZDDrir83+6Ebzz5h
kICMRVFZWonsqWudxOfAEFORHb2ixO8bcxANg68CYVgRq1uuEfX0hIAVUgWc
60gFgMaHpC0HL2fFMpZqEQ32UCOAwNyEIGJ6iqY4QAKSasSQZcz/O3T/X7Bm
LRpGHVHCZr0TIM130gPvDyXepHTTMm4XzP5jE5+ArAhXYGa6bX3wztDs3lSf
PMSv1D77VlCPUHaUPuyaoZn66UoErDl93AZRLZEXr9DO+/GumAPIFUTBNCzn
V4Bd/6SBQcIkYnJo0S1DGpknbpyYCGxxk2+kILkVEOuITBKED5eCobZ48tjD
q1nHzkxOWrWY4YkphFLkpfqwQE5OVKQfqfG5O49mjfu89YXSXf9CEZh4kWST
DjIGJ1rpbf0gfREEQb3BUtcxFyaKy8050JCxXXCaErUe0AExgsQ93cVj2yUc
Qv49GjNDCrGtm9TPzKTNyyt17ls+thNBX6M3uHakrP3K5YXJoloCgbFalVrG
u9/ioO9n/kg7aWl5XR9CXiaru2I913eWgrOse6YKIj8QmkTzJ8YI+5f7mkiG
nR3RgMvk94hRo+fH7zkOjjxi9deHF1h+Rz4AoOT3652PTtcKjEqa2vITBhrk
9jEvFapUYlOvOaWMq3K9gX/YNiCNYWvjvzfXX+5ioFOqyO75CZe9I9DviHHM
d1xEGnwVd3y3urpr53c38WVxzamDlcZWpPd80IdPX1Rv08k1RqjhArHZOv1J
OpvWgeo/cOWhgok7yzCKRriktP0qIAicW87La3sz1NbMjLR1EA6VEHrlC0RX
ljuNFrCZb9hNpXUlXjCw43aO2d8hdLw/PEGU3RlwiTQ4kccihBDdEN8xfiIl
pc+81KPTezpRkuRBZg/7Kki8E82fX37xk0J+/QWhTTj+RCqF42dstpBzk7Vk
5uUI1GvvuD7yKtkDN4kVtlKJA4qmqYpNXnjKtHryvXTrQw+VQem8sIwYBIQl
6Fu3rRoXO7fUG0i46Oq9HD9p8gD1G3/ycvJwQT+kJV1dtQG48wSMYBBIRZJy
Lb4u/0+H6Yg9djmpaSpjjZFe+uO523DhDVZD66LEsCQKvHe/zHBHaXfChgRj
9CB3d08tPPPKwTAqFU8YdAd+3+2cw+RfKiG8xTsPgJihN580IgzlQ4s3gChs
YCNiU9SxY8hkbsB7H+YLumS4hONT9J/2LuiwLDoPqbiD0oO1EpkDXULKbb6R
L54O9A1JLmJNB7wEPfGKerHdl1g8BBcSf2FKMpQ56rk0SGPtNo/9Je9ss+8m
J6y++IuXJ42C/3oWU7+9MsIm0AIVXcxbwZlT5En5GZJi172r5GaTgK4MQTRf
JSkin9VIKsKlUH1X3ntowzm4lcFCXvIcvGqMiK16HIHaEd0LaEetw2WApQpo
pZUq8rAEYYFf78Hqc7wvjri/3Z6Yk3P3gI2VeyXC0oiz+WLuiVsNHlE0l7Ir
r2Oj+Q4EFoH7cJjwyNnwnZ+CcfVcrYxfUMbCBXVmeUaH0THdY5nX0KLZkwDt
YqYLKTGz/2PUzG+WX2YzZXEwrqdl92Q4w4RKZxKo3SqWPzy3zmD3v1az1wkJ
Y91qN7Zqd4s/hCyH+XWdpQMNhlaAwcpxzKKHzP1eGpAvfSnAWizOp0mPljXY
HPYdLatM7cRuZ4AAwFPvED33F5KlW1JhtDhCfzEJKLSG5th1zsQhVAE9Keao
SpFBu2hnH8A9EdijevRjZbHteT6U6g+l+5Jr5WkF4kRFXMapjC0QefvKorgs
8MQAFACYbD2CgtX/z1VSmqDr0d7Z7hOezHtyCQ4IOu1aEbBhf1TyihX56ZWQ
2S+dzCOQpCBRhjVDNQRLL00mOzXNNuw/UPJ9LFZRWAD2lAPG5OBLC5Il3e1V
lTvSeXUk8ij0OBgoHpohAF39ethwjsECRCvavVjg0FEtOziXXH5bMaS+9/vh
Vf86WcD9umJCpiVGMWBrsmUY8zB+C9P6X0PSWU6xOtxLEb9eNqz7v1AAMApU
4Epsnk+qOWmwNkQnx5v9s6aUf/ThxeZK0hbVhsgAptv+dFMiei/LtOKyyY4q
3qWqAatFDiZCQx/8y2+9aR7DMt445snnRbFC/ckGEVFLqp2mfT0pZ1VyH1ie
BMgFDuc0sXocSJYI013Cth35sLMTUKCYis+gODOZpzgKpF9PVp2uUfT9IF9G
qQEUndffNxmsmFomUJP546Kit1A6HuI4cw2YZNX+/c+bWhikdiJs7wZMj1ki
kkW1kfljcmMQZBQMj4rmy2DlXEwnjpU++CFxT4mfaDeTIfr6i/WSeKR036EZ
nO9E628nQHfuSr7KdXZwTEK7IlOm95+/mboM0rvdLFJvcnqQZ4ICBrHs+tRQ
J+3XfNqNmihV7ttm41g1xJ8cmsjdc7Gjmv9n8YlttsV2eNRRY8wmywB0D0ep
GrdYYCF4Sct2zkJ8BVlQ+ycoOQAp3zRAtdb2fF3RJPUNWyzqYOQH/Mx8uUuO
rEKEyqKBTOxHekiaJif8IHCMj5VLRDAzF21IwIp5YLEDFP/ahmMOZuvtzFK6
AeCRcV9aGJsd4cgjIShar+hMkVuS4p60LQjH1VxBzWtWUeK4MCNNRWe3hgiS
kQfhQQXjEa3b+oVD8VvnHEejK2w3pV2fvsW0LUTMWC3QGGmSJDJV1yOoaUpk
2N8uSbPA3HMvxacW+LBGIU1eIQgmHlguo2ycaNLhcUOFclQq6jRNgcdneLth
QPikFpEFx4rJPjYyYbRP3BP2h5VrF3fbEi5OtOi8WzeT8OtJhT0MM0tJr7Yn
i/+ucbMKFpMnQIE8OC3yb0H0L837a5PSw2grD10vaALhzeGxRqbFjjY34xeg
KSGuZssYhkutBQ40ua0/WYvDgAK++vfu1sGP7ltE2a7Oms8KsoXjzi1x3BHJ
dTV6sVPlZwk6nBr7RJlvfoKs6y0pZQvuH/yhtinHlmOq/0B8hSWHQ++i2unG
SqwRH2p/ICPv6Bsg0qN91s1iJ4rqMZpOQ2jWYgMPbthWp55AH12ZlalABWzS
OplG+xcCx+dfDKcl/V39aDY1j81ZgNA6vZuyv4QsfWgVzRf2ykQxyWrlh0Hc
JXISfDoOm0+Sc6ZXfx4QER59ekHeD6uGQReXdT6G/Uy6tIEKwbGvZrqYa+Mm
35eVHq+sSiLwEqKPXMj7FM1qmbyk40hwZ0IMBH2VrYndfSjf4y+0T6f2TpGJ
CBjIEHnXucU47STtRb6PcWgzqxMIQkXM1i9eAYTi36TEmyGXIeSukigaBcdl
q2+uhYjEH/M+25TayXHpO41n4pCQm9kBtTMV/9LQF1ZpDeUI2j/MGDfhzymk
sWPLw5vAfX8rlOkFY2h1qVVMy445AlxhlkRxrQ6l2utPn9EHRpNf+B34/yMz
oOWnJYR/oh3L/2HVnw9/UuI7Rt+HSGXP8O9dmyYN5HcjrRWiGc9IhZLzoU5B
0rZonhT7hQnOR8oLZ/vDSUeovynCw2nO5FDwZw9Kly7GnMUfv8moMvMUyPPV
pBnTJtyTuYVhn7C22HoLDSAGAjAMBXXO/KmqerU5pPr472ktqiMHImz6Uj43
rDeh2gyrTFiBd9fInxWd61yFMCORNEA2bJ4e/rsbETydePVuv5se3gw/3Itd
i5mjX/LnN49fSMeasBFI9Qj1UIn1Xu1WWoC3O8imwq5pPApmyM8jH4soNO5e
3ALfjdyEFbKeFhisx5TfTMUsuoiPAmX8peDcmk6b7aC+12rRCIdXPBGJ4gAt
sA1+OrvDduFgK3f9qVXM9Sc1IWFvVv5x2akQ84ieQMhydmJMPsExdEB8tBDA
BJ7sZK/Wry9HfuMmB+SMwMeYegNfBl6btJUHL7uoMFJQKPRXKkeuxVJCyj2l
CxyC7vyX+/y8xoRLGSBv5E+9Ui1qn9O/JlRGeO2ph4/01al4KT/yvBV4S/1N
Xm9TxR70iUTV7pA+3SaqA/vxmichk4L8ZxvqCqggtqUGBvwh8Jr1RcdDDzcR
iiMi4cnnlqcX71uJ69ZNTJh3QNwsHtnJgyhSSB8UoR/YJdwLttIS+Es2z2CZ
1oyjUsxDndGJTNIs3ElqMw83HlfZA4uF5CpMkm/vf2aCTROTV0bv/K1C/VZq
BWlBPM80pFIXxYOLjKBex5gqZLJHlOe4mTRCyV3/yDQ2i29moRJmtk3wxO54
2vLQAXR0kG+/TfR4h7owVkACQ0vRKI5IlcX9zwaBiq63ipVWG7EX8Ju1BHFE
4o/J79w22IeG3Nt1RmAPEo7uiF/+1IBpCRmK0DZEoZoceurXO7Mzteg16XTC
yCegjmEUj3AyGVpV+Hnllsuuu+Bp35zCsUsecNL6/GbK3M1/3fUlKpHzqXKs
olJEhOY44zxJCD9D2rOQgqgxhBbIEPfQH1lgP5vQ+zPhV4Ynnr+OLyV4eg8L
mXFDgyOk/HO3rqQRAw4VzeLORlAaImjehCFJ137IBmR7fZPPygSyVboHN7+Y
WYFku/it8RaxlzcmLnC/OEj9PCkF/AexsA4mukF9LkrP226r0E5ivDrAE4UO
wm/nVgTUDnP85bSBGa36k9H+JjI2fdzl+yfwt3Yxri+RZRbgEQR5Y7Kp9JVg
jZwzRzO26mPCsztUMWRK05rlCvn75LC/Da31GYuRSiCIp0LgnZ6mCqy/2MTl
eSnFZQrU3RnMBzJxXevgUr/+oTI7eO3kCAgdMmKGcnLoRmPPcqR9MSeKiBpn
dr+HkPjUUi8oiFN62TliVHMB1lStOSfecyRhDlR6uylNFjzC/GdV/x7jEn16
exUc2REd3yehtuKljLFk3JxqiU+CANpiufZQVcY6RzMGnS1zT3UehBpkx3tC
r6lojrLC+WlHS2DiN8jkW/IL1q4IQd8j7Lsjk1LXY0w6DPCAmAi1EVzSjexM
VMnVmX+s51PJPFqqAiSMRtAWuDqw7ZyqeecxJaBO1rrwm9UnIEGTi3gVRPW+
sV6adR/Y6rdFj1j7fbhRl25D7/tfzjagQZ8g7kB0avBxR2e/oAfTd4hTib2L
P3+uVfgOSrBqYW57XfH6X3Oj+9y6JUUB5UXvdUSGxfEr89H/EkLcYEfeT+W4
WKWIPFKzf2zSvMoEzkr4K+5fOgMM1ntWEiJmw1/sMSfrfRxJiXpNfC9HI8Em
/U6irBK+49zpRDEQq+0tWlOTrVfdpmT/4rxrZineMu2dkVVjc/ovYN6mNquz
V3bkYh+M1l5nzXaxEKxsxSEouMeBtm2AoEifoJ+F0alaePgaQO583mj+jyVq
WZCWsWr2ML8+CUZXbxZs9XIc5ABKoKwepGhTCY6pWPs8QJ5KJY8clY4GPWVL
HVp5lQBtFpYhQY7FJtaJFMtvMgrcyQ4XNjEZEN3GH6O/OcZ7sJIAZLVSsxXO
vaUJx5z33Epm/B6q9m2pkUANH1oDszor/ntweEzr/PK7V8n8+0sGH1qZX5iN
3Lm6f4K/A7dPCuNrGimOazBWCHPL8iQnnwAqfeipJp3bx83rKMWzEqwdQQxB
AukXRuUCFfHNyGptlQdio1nBjL8dfMYwuUNB7a+bT08ylEkdn2dNEn09s/mR
zDw87L2bDb2Ebdoq5hLiaA8whlCPLW/ZjEcGVECrJ3xiDgluDrPn1Qxj2swJ
ygEGrJISegQtXQt/vpPS1yvarec2S0QZjwKup+8mA3IvDQa3hBEVaBQLq35g
d+ERZr32aGqByICL2dcM09cI420JvGT0gJdkbC9kc8sfhh5/WXHV9pv0rS4c
IyiXiLJeAe7oRtB/Kn7QXLnTY8HscZcruk/smmT8DBy1AvWsyE3FTCJniT3U
LCVCjsFpCj3JSZPq4SfN8i1ZQTe9fPlEZEPP8CGsf8loU7CNZcEOo0S9EkLu
Dl1uXsg4MUcfEHO385UweoFTKbhPzFlWevYJ61UCbyWmuut1ZEMMngtRdELc
qfZDeQyCjs9HkwKPVs72wMO0sHSEC9rVjdsJMdb5yoFDKANnEF7kgSRPc1v+
NK66Rb9MzetnR0dIexMZ0+WAp2Zp5SFnlmMoOJYDo9PvWX0UM2e2AfzLa1ll
yPBHUQKNkJ6OUzZO+F70NTBnbTr4wk60wdpuQr0icWJKT5DNysU5uJ5dV95/
61WiLgLzOb/M7XFaLE7HU7WIJaOPiX/yJWNN9POnYZoW7LVUZkf3NT693kZj
GiuP8vebd8WNutIBiTrw3/FhB1jerhuMK5WE/2Bl3fRpEhAA2htRorbKggMb
cDjQb866Sx4MGZJmj1k8K7JDM+Rs/awDNNFf2e8LTaXnCcTe/ry36OZE+cnt
9gvZSmvIDKEKc9zK+bG50H/GMJ5aluFsj5RKyhDWoEZULb0TtYVO04f8mZyp
h74O1CfXJjKSqkIBjhSzec2b0151qOPDBnAIPhjtgfknBMZkNXA4XfHftBjZ
7bxs0uofgDQr5C4lw8eO5vynM8tpTMG1bL8BDbpWsOegtRQtRYaAJTScYVYQ
zlKcwg8SIJU+EsHKoOFqRFnW4D20gfX88uKoJIgypvDKEQ1QnudrNPD0eX71
wOJHJwCYtmVBaiIfo7EH/u/I42ghLUho1kUFyHnVnaEXxkkB/aaYwc4QHEPd
0REAWEhFKtYYB+D11Barw/6ayHQ/stYOE0pvuBvEr7g5Zq+oOHSXN0gqp1j9
jf0W9/5qz4GT2Bh6pIMhvZs35bO0YeDgykqtg9pht73hGbyvxAwMAPCrw7Vv
oOtmKaUTn7jp1PQtoWxpswxUNmepU+JQtypHWAY2PWqO4sfyJqTV/hzx8zu4
cIsCsDdcNHsi63lwoYq1oX++tXopGeqYNB2q2OOFGK6zChjE0WAsFQJWD5rD
HnfFdvdJhWeHEBYOm71YyoH5um6p3ST4EGIzGdYOZrfyR9ACy3yXs5o5/TMW
sxLxugGTL3MMMoFOhnMCSnG/hTOimkgtgyMBc/2I4jyNHv4GkmPQWi2U2i+T
NmgJt2UccLFKsc7O2liB5Rq81bu8drIB3jtoAmPrN8gK3F51jAnjXjh4mT3f
eKaeXfQJ1c4DgfxSSnQTlwJBrG6HXPNp0FTPhUoEGGG0EGvuHCFLe5N+tqXn
kMd2hXJWXxSSyTIwfVTYmmokHRn3lqFsTSZTZqpP7l1vcFCPHEjBI/2bf2dw
6cwBaB/2gE4b+y9V+J0ZqWQ6F9peYkbwIrYrpR1Y+0XKVFwyRffeiUQKBs9L
GcYaS9j6LECryVzLMDnja0gEACcZrEkK1iZMOdY+rBOn+CzpkhdVgGPSUK5Y
FEN2YvZY5CV3ysy+2WjIjh9JRljROr70ZEtDMaV6NUuBZiDx7i8BoFXE5MbK
5WYP+bhf3s7xJIt91oX6tPAZaZj41SD69Mp+gHe4Y/ugL2wVEG11VOKmTLmt
9qZPl18zY+ewLyn9euo4T2JB44XqXU2d3fLLx7eKV2EdtmJBRprkt8RgQ/J3
1P6j/+zETTRm8RTz59DVkF9wRI09aF6zpUIIebfWJp0duLjS+y2X+P3WqaTJ
wkpg8B7CAQ7wfzZFKUMx3of7E89n0PPo8Hs5LT92sVV05UcqtmzIKqKjIX8+
g7etg6D7ZG2Mhr9MWfFtaFSRmNoJlI4B3PemZTLdruRNVgNMlQGC4pnKlQf8
4SqnF4gH2nsoFZ3/ouhh2gWjHhLSxnlwtN3luKu9QJAaHc+68CpdXz7tpntS
da3gmmAqxXbZBqcDNLA+rrrj/nyepyCqU8975HU0H0hcx7YJsThxFtWbPd5Z
kas92Agj7jt66bnM6oUS2qu3C27DMF/KGuhwmDzPDd5vO0hPrWXHTxlFhfOp
JOL3v0+u9JqVP3DalKNTWA6v6Dy5BECEa7mrkj8lwmfVWJVZ0LfsSGCh1K1P
rHrTdywaNGqCzQKkoMhTERcJqUWQi8RccwkxjjOKJ2s54ui5LStnyf1NnnQu
uiWNZJ4jCFbI1lTipJvW5zoNn6Ri9fixKj5uStUJsJ5vtw8ONSHRBrehc9ry
Em6kEQWfv+vn89vWdiPX9eAJevc1jJOiz2XHxll7FCP9XgMorYU0PWtwNBCa
nuzfd4LxisjMw04LrKcJBbh/bkQRQZ07WAdtTVALFOOXTW+U7QzyDrAx9vTJ
nC1NpDvRin8DkRcnqFmsN5sGHRNdEaPfN0LmyhcCNmqtVrlf7Rs0u76bp9QR
S2Xc6rSVFTXyt9FERyjXM5BK3Pb2MZUMrT29lrQvYS6M4DnQdCa+Msqv/2nm
+w8gbH4KEFD4H1pxQ+e3x4A3UIUoDr7ibKnXuWrymgYHPVRBF22+bIGmfUrv
xAP5jQGTe5JAtNZSiL4urjBXgGN/vRXJJyo8gqygcdimHPwDhX0qgCESl7Aw
+sqIV0Mn381dEapDofElQZhOKOCFVyD06wZwuZGjZdb0qE5yFVpBIX7St7r0
8jtMncZSMWqMmqJIJCQpo65oaS66QJBldkt3bnF+SyiZzcLFHqfs/U3TtaQ8
sPzUFHX8S2HgxF3xYEvbw37R+w6bnNEyd+/TQ+BGduyYN3kr5lir6mII2NHu
rnpHCsqHg2jfYj2Citg4dnIJDraa82pFfiihPMMU60KgkyqX59xlHmq7bAsU
psilc+js5i7Ctvw3gAzCz31BzWitKzDCTRpJkouRj6BcLNPNS6h6rntaWcss
PP5ktOX3WTmgsRiQ6V51E17Poo7JAvZ2aSvwlb7l8fARpEr1wjHRYamW57cw
VqmGhfGPXdE1TGy79WcHF6VB3tuHSIpFOVnfEGk628udDnb9fmCReZBgwYhv
x+vOJ4W09jdprr/K0vllPCmnm81dAx6fl+3xRTtw0f2YIH/TFsGa97SIznWQ
QvyM7uiZd6wXPEXS8q7nVs4OTy1Oux+rAZi+jI5ReiLksj0gKvIyeb7+OIxU
cWyXKevau+82HRB8KNHu1ZAlSdi7FjrEtHqxJstOEo+ic3BpuSZKxvUr7yrP
EStJ2n43TVD8tl5pURR+moeT5oyupl9efc7AhRDlL50+W4Ekk+4JRF4nt96U
Q6Jkn1+DENWuZu9LKd6l9AUrdjENJ8qVyRSr4NyxA3KxNsBRO6MRlkOlIuV4
4A9cHC1n1Nqmk1zCvYEqbXcjyX1MpxwxY2fcCjynl0Qzva8SRamLJNBsKtDa
JS+XFD0f6PVxh4bUKn1t7GlMVzIeWyJtTVVgSisvhYvMylPf0BP4v1D1PCyW
8KQaEiUOEQ1YWd4AMgaTFXrpkKj1phH2kIFkQ+MxS44lizCl/UiGmUQV6sSB
BkKx9k79Uphbxlrw1AU3ii0KGGSCn7/hoet+uwxQZm435BkbRGGgJo1FzzfJ
EkgrCBvLz9CryzMYqMkRyKl+uhrNUasgTV62vOVU8M9Pu6Wqt00KMLG6LkOq
O4AURbOdf/GN41TebFd+EgUnvG+xQR5JEOp1xYmdy1i5SaQ9gxKcAyVS3Fqm
pp4hsQZuu9icjOn4DgetcrU5c3hZ7Mo/FJ5CalAsqBfqgSaZ3kD/h4lROHkV
BBWZMNFULxQbWt7EJdUZrTQkat8ACuaKqotF8XlSwoUjtiZNzPDiaTrVFn/N
cREO8VIkJjJZb2o9n3taegw6ZPIfNXzKqhTUcCmAZVPCe9d+U4VDXmgslT91
XqJXOGuTygSAeD3nWvF4bzSey7invzfdGIWvg8c+pG8BRvKyg5pu0lHA1PQv
Nnf44tGKNAgythZ21NoYHGUqqzTW79rlitKeVqKBe3ORrPvPbQFgiDNLjS6f
5u3h1no0no2RrrUFdJyIAEOSK8hEcmwPa8d8X0CIceMlYdiyYETfRXei+Tlo
EKJnIb8OkvTvPQVZgdpdmHyyr0FMHNl2D+eV/QG/KVzH2EW2gcqlJQEepnBL
v8otTVrkzdb0L8j5a33/mtIatazIR+RYfeFZajoOMSusUbsG9CqcwiYyAj3d
wW4YJ8t8or5AD5UuMd4p4EylY7yBYf0SSx9NwhWifTMJR7ZLThshlsqO1dXZ
FnQecQiruDihiUlHWqHZUOMiojHiyWnkKznzp6yzVVCIcn6Xme3dGZDNuZve
C5BNKSbaPbs5mDieBJ5kCRduVXGLBd00GmRF1/u0memaxxWDD5c1rNRAypDw
gfjuFDdtvsLwFVs9G0X6T9qYkGTpfzfTMsKqXIhpRea4Niu0YhhVEDezJUVG
sVGCe78ECiqhUVer2GYRE2Ev/bgeuBBm7hDTUhG4RuuBFfcsMjvdMa4xtHx+
nI9DIMuw0P/u0RaKDXHwtHOT40+UP2rjEbtkJI79BucpMu0tz+G0sXeNW/Eh
CY7QFEsPNsyOWcuobXxu1Nrfd/5HxxbwWxyafUHOLNbKi4mi50KzXrlOBOlj
J+I8K0YbVGH/K6O/coWE8OPMjmv2RunsgqGP7BLkaunbvUlZrGat6eynGqPI
Tc22it3jonjnYNlP3AOhac+HXynaxB+X8FBYgqE3sBeVWwvM1Yn8sxfQqvAc
CD854YVZbiUsILNX8KXzQPAZJh7tjg/NeJwYu4COj2T9prIWKx2FnYv/f5i5
brBvxgZqe00pq2wZaIwiHXi6zNKwrlbceHK85ppvlRRMfp4NE1Q7pQo5YGHZ
pZweADdGLVVFKlCIH85I/vR7x4q3Y11Cr3u8uWrSa6P4Q1msZSeZDEaDlBDe
ryh88qlDipEXugeEH8rzmrUUs0oHIpuFPqN97ZtgLNx52ADk5zG5OXyKdI8A
hO3rFI0A+jSXBdHIYQfdpJdAg6bE30Fw4ZBICSOkOkbBT55NQZvMlvYYB2bq
rD/0UvvYS7CXD3c82BvNooMthQQaXiEjImNxkHz9FrD1s2kbUTTBgyp77CPM
575rlfRgoFQgvCsAHl/Kf2nDBrJ+J4InJ2HiKgRTRZEpVYT1+kfBewoNSn5W
6APRmJ3GQpD5vKiRJV6VgxDmVsFIqRR5voH6S+zSeTodWxAgQ9C4Yq7VyjYn
eE77mvW1S+8MCOIhnG1PTyVEk6lmGuWA46XQNmAt0U7EAyqG841lxaHUuGZc
7y23pHkTxEO2w+MooZNRzxlNYgPa/5OyNW+yovYo5ACIDLsSPvRq1HXcjFgo
l8tt6H9cY+h1HhIZIGR4Ds6xus8S3eEXsQY64iDyVAYcXCRjf/U8E4JHG7kP
nIhXB3sQuMdg51AdzLa2gt/C1iD/BM+diJ6NQ4yq7QMyD6172jgswAK3523w
Qm73ZZdnr+qXx/k2alLYi7EzSqEcDanwKWSNevLX3tSuPPBKDF4YBK4uedvu
bwZLT9FQFOsvjEd42pnG2b45gcfnvRST9eI0QmMTsXhxLd2Rv79ZAfXIECc+
t3jIlg3FPIILuMrKG8GLmt4eGt5h/JhBYEHjpRFMzJVU947YW98KT2xGqFqy
vCPmDj5urVK6qSZVXVL19/J5CQqgZKCmxpJaIbDU1K+PC7Q9RiuC0zSMJE1e
MANktnPLgzIpcvKsvO7plRIvEFnZODBBhryqNk8pslZ+Nli39SrwakYpTzlJ
uMFSJ+9JeURwLz3WKHKyat/+oTThm9AMNvc6CqGPzHdh5AFhxa0aoG4YC6mG
Hf95lFe6lUr5X/TYTTVK3V/kOuX58R18rpGqsJQyV+qD+3awV3jqzzdSyvQJ
kjyg3VoalL+AZCXJcCeSUXpRzuCgBeSAG3LPPwjRXWJ/G5pJauWp0AUH1coc
DJK91p7jYYqV7tjFLBXFpvdg5Dw6YpW+0wg7dkEoVSVozX3tMuPqO0iX2BZH
OwgxFG1LuqHVLrfmcXezP0rAfkf26WvKhGMieNTGN6WrSK/Til7N8UN+Ic6z
9nnc6kdVWZEAS1kDZ3DZiVFtA8hOfQioEPd0W/4lOBNn4Zg4soigRjItEu73
niTxSqvLZ8vGgOt7rcSZJz8ppM3suueunyThxiquxjBqdr4TjWaJqBY3WVTP
wQI1UXmgsY9VNkN1GKWmkZ0+h8tF7jgGsMoIgRwS6qKMlH8o3fRszzh9mg9+
7jFxbfEFLnFXv+qJKjJS21/tWFYzrvphLS+zzKpQ6+aYnNpYP9o5fyrDDC3q
D5N9Dm2PFdzfe/N0TdGsxnin4PY2FCfJZxaq6wD49dlMn816yytNl8wjxxli
uzvNU8t/4wuNPT7MxRaw96s3xZu1yyNUx+KV+35+nXZDOWG67R6cpCj78W2D
zouoXfxTvKrj+SqpJZHJgFDGy9kKDAhMXe1QQMJkTce3HpGq0EDats7T+Tcq
09JsXBvwYBcn/BWYs4k9Tqx9TfRj8qzHSNxPPhM7aFe4BB09LFt6Yuipg5RE
3+mdPeWjBkZkFsODzRqhfpATPK5H5Noo6YDHgoor2jmor3GFJyeGqQxp7Oge
1FtGExG8+w5oRoBp/pcFmCtgccsV4wWXaMkhYQjRs5LDtgVGpK/3Yl/aoKFI
Z/ZhnEUQYgaYAWh4HzZQ3NXdzeSQBZ2w4AkJygpagthFEQRkFVoXmdNJHIy0
kCCsyNjIgzoioK9ouD8sKYl6V8kV8WM0bpE9ubd4nQjx6l0eyU12NGE54Xcx
w/uG8kHQfZ0aX4od1ggLHkFm04iRBIaEySTkMJQrYbvVHI08459vHr4pWtGc
9kLjsXNC4KmoLQpyyPobbh0IMoSnFZOu5cHBAcveKCiB+2Uk/Hwntyz7nqmq
gHyfqslcHCbND3swyo/kWRT8JJXBUBKbjsKnybbNUWlI5rTNyhXYrvAOEojm
e3KL8EnDz9c1GHv537xcAHGBjPxeULd1Mqwqyo+zxmqMOSDybGgfjmw48JAi
IqYonr+gZjEEUO2KzCAVUkNQrt0sQkblQIoxgXN6Slz7uoNrOCnSd/Yvl4yZ
9cmAuuoLSKenIdEherVhN3AjhrUu3jrM9rVXjlx0SYgVgtG40wEGu6mMq8Zs
jQR9oyOPgOqYroCn/8Pi0PTJCugvdehj0ZRgxVDXg+UmJaEAZ+fCTWhCYXnm
BuC6mfXWtFb8YetObcJvOBNseXsa/BrAJsCiA8DxMhojjmJ7WO8uKJu3jbOw
2URAWHuVSzPZCpeS6Zg5ZlRAOMGKtvfE/EUCGT9sHo7miZOBqTMaSRsnrgU7
mLnF4eBPEzpl2xGdCHXn+ZqdaMliYvhDl1pFCY3HHX7NOClC8WFsHEc0LYc+
T5mGXtjm7aqbmM3zTj3NO/SM/I+5ZpE6GGRQv5pA1enCydzEb5NtYa+LVhSr
vmeQBiNtbl+gdY6Q/EnCBtDD0RsWILtXoWCswj0579msoy4RXWz8DqesvpaE
7jSXWiKCdvZ5WChQwA/U1KySQZEAr4PU4KHbaMlr+Zp82CPSLM5p9H1OMs72
KPoWLJJRuu/iVBi8j7Fg9/uWwiQWX7hMuYAZk4hK2ZmVGJt+n3m8NJ6gqV9y
JHFGgvwVvtsog2s0K49FW4hRIY0RrgP/Ckaj/tKH0yDJdSkA3f2sUC9tBg6g
DKHQHbpii2q3f1oM2nammjQ0SG9rXMLk34ve+6fboE1ILd6yMtKE0jF70vHL
EYsm5dROYs3yksFMBzF2c3Pq0oPxZ0+fIJ0Nat0RQM92sLalkx4CzbOwKbN9
Py62JpGREsxg+Sl+mrNGpoi9cT4c4PSC5yWkB8C7esT6xGrIU+Z87o+rjGxr
Ahp9F5LjfCYg65mD4rJNJvUrrdboVLIdTIILlRjTMke1WhP+JCEoevK/TrAN
9US9bjxev9o+DTGKSp+pURHKYGlW0XM9F1OiJ5qogPAtdpuiMNSwy+AdCchx
Kt1d7eG8aMfuHOsbkQajpJ8uQyjUBnaG4RUW0Z8P/KOd3a+R+mylyT7ABbF1
RD0GKrFRVjM/3SXoTEggYYVoFnkBLdeMwgaQ3lNVJN/AZOXNQWRk91bfioad
ghyHuDUwLw4p2dRg12Y46GMiOZyFjKYYAYCbG4To7QBhSTd5bUxPrJgWSFH4
69Luamq//QBVUMmDYDuniF8XGHVcEDg6Bmb9ZQYBpwpWqPPV7O3mdCOVqUIX
8YVIeaxxx0xPs4Xn1J5AXg2ih8usQ6/UKtshVqlcDMIu6DfNPHa2xKaSBwGu
McbbBdrZv7WGqI2R2MZlUjZXlW9GXOA8Jj+Wd0rY5MvytGZfQ9SMb4pjwgsf
+vY9SKX/q3OrQuSHkGtnFbAFxO8m3coACAYx0D/I5UucahVu8rK9Nvts+5bJ
18c3F+imZaE2GRLEXvwPg9EY2dIEAApET9WllDRnQl0VfrdLjp5fE2aGhrGy
SjPpegxrWT7BSdlvXt1qjYbmdINxMmlKN1qY/Zk+hT4IjlJ2nMD2sPRuUUGt
40tjl0zRGv9lG7gyaLsAJNN8tyPbnMMYgYDj1g7O5jZg8lsSO3cu9EtADuui
Xkhv5SdKH1jLGk5EbKxyBJLxy6zWYGPWj8MtaujXKNmmpcaXPXtBVtLNTkAE
1C9li2nEveD0rbp5gUzxQj6Qgw7aF6wg46dI8SMJdEJ4XyIwhVVZMMyc6wF6
R5QgJ1tSO+hzni6ba8LAb+Xpp+Gffy+vIEFMF7YxozxFwF/mqgM5wVMKAo3j
oG5YLfQSwgVGq6oxfKm3JEt4G3NYPyN2AkPiOZG1j/aQwuolUo5QljE3nIQx
49HMPwNbB8KMlX0fakuOV68qQ7gYSpqGV9MIh8gefFPKnJDCa+8B3f4Iyfnv
sUTVHuppTRtkU3tymOaNn4xAVKHIBfm6KEyX5tySk1Tbu+LO2q0E3NWCv5QU
gK8bGBSocM6V44J81j292S7iPspvS+4LVAFkfhquLe05CGSXK3A+b/6exItC
ypnTb/LP25AaaLBFUZsBlqHd8GrIV8j4BIb/jNLSB4NH9LlqxfXh+rGEAjL1
8Ojk2J75RVzglXJYMF2MKxksUm1Ng/jmsJ0Uri6GnDQmgoX46dF/v1G2gjqd
te6sTVx658sfEqkZSh/s1/QTSKQZHocnmMMYY6PcJjuszoTk8uBW7AhPHqJJ
8ZJXnvzVsmOYf7Rge19Hv+CiR8g0u/RDW8K01PlkAmaLzDj+FF8uCTIdYCc0
bccDJhSvTl2I41WwpH+yeJM9u++PvuvjJeFotOzfpGodKJZRFq7Lc1aFyZ3D
FFHYmJk18tH5Klcvnf/aW1m7f1pJl/CVtUA+AS0c4WVX0+eo92pLWbDcxkXC
vERE40Lm5d+QYXrySP8SqODPK8sB751qblua45eD4brb/8AY1e7wruYlBzvo
/VtZ5EI8KIr2lbt5dhsFsJ2qv8s9sAiGCIKIEPPZyFTHB2O76zQ/YVKhNuZc
gm4PVH0LuyWI4jq6aQFW2I9yIPRq3yOco5OYVbmB77TIBWIjKkDkJmkIyy2R
ujnteBlioFLNkrEDlbOCDBKt9BAHKQoNHda5n7/rUYJomIQPv1z/MXh5XZcJ
73w9ZSkE/yF5sHyo4eMoyJAiVVC2AfUo+S9lLPc2t2/umVa5NU2Je5Pi7Pry
Zz3eh8C08TnQJ5tmeuse/UQQOzIeZJT5CgE4b5lBBldIRmcgkekYRjP6l6e/
3+8hA/Z0RBrtXhIQHvMFr8skdfIPMFvOK/HjRYKQHyWiYLxxZB5MvBoPD/d5
MixVSbYWb1ReEm6mgsj6NeXAb0uLPzRaSKb4F3qO7L55l6NlUwQ63Neq4obm
sicVn4rI9SrJ9qjCBwEYfz+7pbLLpYMhaiMxdtXRUNo3R8/4as5LxmF0c1ye
vG0ATWDFW0ahwsKEFAfx/EicckpEcHy21cT9VvYt06qEIzlxtx/onBRGeU8y
Rm7O/Zj5pRuMzRK/XYDt4snxFVX+Udh5y6i7e5lhFVPQBucnuPpDroip1HFP
j0tYhsG9sTs6r+p3oxfvcfjnNSro+mwiU/15jcwbEiC8By+smhdVXBR/lFZY
FDOiVBslwPX9Eim+ljGfGHs9Zj/rARibhix/Mh4sar46/p8FRuVNzU9T8EJg
JuvC2SBb+gnXhHF21u4UeOvIJH1Oad+8SMcfx4XjS0V3zt1G7ANXDTr/myjD
INmRPSBV/NMny+KR7TmQYzsQBF7uhu/JkK9CW+oXzVDGdXUJg0XEIrwqcG1t
xDVx3JJS91ymLVMpzpBsy4/7gu5HZxd8Xa9NmMEmZQWOtXT90Jd3MSPpoKHm
Mvanul7ZFpwCA+IIq8RAp+7TNcFfLP3pFV5D9h80duhmbX+NBFHPhdmbl1M1
+kpkRLbCaRMD1zK6nnTyRmXzOv2rcHfV6x5wJdvRlGDttI/ALMMOo1cTfWoR
dCxTg7U36Jl/jdkuyM50vhDkLGInAw0IIWWS/x661OAfKhYf1q0ivqZW96cT
+cjqZakQ57pAG/mfF4EFbkCoG630BgUzC5va2O9xfjR6tdceKHoYnr7Ri9ai
I0w5Gi61Vazbu+uFkIbnIie0xmOtRjlTW5PWODVz4Ql5AidsIxP6zJBilSkA
kUSiDPGldAXETp9Amq3JRDEXrYow+hohKDIPgKC3QlEJuZG47m9jO3LWCfs4
CdODbseVEbRM0fdEqr82AbnyVE2/sX0FU53XL9fNesp8d8vnDG55o5VNoKpa
txMIDbDOHu6eLiE8Q2WNas+FKK/IiFJDEh8iXK//QdLAKRHwv4pbf2u/WPAr
CI9LdjsjS3V5SIDUH49fdXS3sAn8qziuKmJJmd7LMGaY+W/+j7LMXVG2p+Af
71vV4RVe0vpLIzfA3iUBCQdiYyBQNj9WumZdEjxe3ZdlQS3GJcE7mXqzfH+I
hwVpgLrWyLsj0HbE8JKXtBeq4fqTDtgiuS5/+PXRm7yWVRfVjCjdkJvOPD1I
Gu3FSpjk09urfnAF3j/bPAynJp1JlWmq7Pfv0kE9edLiAiaBIuGwGCmr6cvn
CvXWKIhBGwYHVIXnXvyQ5cIPB2/mRZWbVmb0PouS8hZGoUogdub6TPYl2liT
TcD+eryhlR35T6qUJRcFr/1CNVPqaQs5lG+9nB5l283nmNNJFwlrGkcRD9rB
b/t6v9k34NEJxKXVbfXeLqKHWbOjCrzQGZQy/TvdrndLWu3IKAyZKLAfa7Ym
gEDOArUMoDR7y2d8wf3j73U93JezT0Jow9u0uAdPcgSdtC8+5bISt2Qa51qb
BN/Xxsc0Y7ftJsxIu4TqysPfuPV50aLu+vmSwO7t17iNELUTQWFScjPr8zZ4
JNFj1JPUwCfT+CjjpN/fSBiZL57Oh06tmIP+1hvlJVsFBHuqgQm0ASMICC0x
cdPI1VNmqm8p4p3PKb4ZbiHR+kCndZSKkfMjiBUAff3mP06KvfEhgucHofxm
fd2CjG0azgnd9DRss2tWJRwqHe9d9Ck/UZLsB3XCd3WtQXLIX7RPsjeDKjR1
xMgAPC4KefgEgSL14Z67iRQ28CdZVgX64dqHVcV/ugRgcfXGJObEHXYcGM3y
K6yH0s6EdWf8/5vS/IvhxV9OV2ZLiucDuBeaOvg1XYoo7U8VrA3c6uba4Aev
q4WdZQRDnV8YHxCH5PMWW+9sCgQkbfHlSK131VrmZvmqnYYxwAkpj9+lQxSQ
RdnbtRyoF9qT3Z04zRMigiVayzCzf+jDV43PJAiy1VN6hT1Jp91y1LZjKvt6
UYU9SU8XgS7Rb/MhJzMytR4MrkjzZmELSdIyk8xCwmY4BIuI3uSLCkGaBHm9
b/61b6uisqdZDPc/GMN0MBf7dyc4ZVpiM8Shj2PaRPQ6jA+84n1pclcgsMHE
v8xRWbLw1kX5q3sAF5FWjAiK/DWJFtHCEhK5axfZr9TUKSDRY5MKLEYer3Nm
nRN3jCRul978AOCvOdIO61DlwV0H5ySMQWDoMJilvk0ZKyW0y8H+GpRPxYdH
0ylJZgRU1jzYyuJ50hQ92WH+K4jUqkCXGJuKIJRZi4S3pKW1uwDvj0TiDcc5
WJvpHHXLT+fltJnUp3LSKjVd1XKB7iMBZFwU4bsOqy2hZtIjKwF223noSIJB
7RQa9BUHdsexoDl4THFqsfnDlXDb5glZr8k9w+ZpNEbKvIktHSBFObl/SO1V
FnovJwZMrC5ddLifC6yimCaaY/dSO/ddpYQ/LXOmhGUc9Oc8Qu0JMTT8qzc5
jzEoe2viz661yewr5yL5SEiYPIVhCOGEBp34hFIexOlo5YL5eLoLuFzyGqPh
Uqhib+ObQOldcg5+DFbLC/lxnwNz5+YnqsZXOvQWEl0W/LUtD9Qn/RR60Zup
bnPV6P/AOA3SOilUE5vlENKY7pdKPB9h/lap4rCCg5q1Rq3Xa+iAl1vmxdso
OyDMgwQKUCsGFwgN90mA9unM35nSN24NLdmpMo92efX/y731fw/jpFKepMk3
XE1fP3bveUu57x+33Nnfz75ZsabCW2ylkUToz8stMkPEBZDDKdPiTDXUBmgi
S14Ei9rM1b7JlHDGjwpiJ+QSFBg18mJsZBoA0bLI58BXg9GH53GBTLvht/3E
vYY/MoIgdPM/cFKsjpP4qk8MoLaJDi0AbySIBP4rG3Zd+hctyB2JsM+HpV0m
0d3S9k3SEq8DDQCeo3KLHtvl3Vl4N70Hc0rryJIXzHLgFjnAgc51AGZHdV5/
MCTt85uhr8yB7HMoX/pO5AFIi1K49OMccV1RtY/V1aVg8erV75OehJb8J0Sd
DFEmmg/IsQnXHn5cVKvlq87D3nG5BGmvOFv8SSbpJGVSj5CpvbXqKIgdtbZq
DMx9mWX1A4cwM66roJ39UAWFn4jgMSChDccGFiZ3pUAe5ihPzGz9m2KWAIjU
+0wqIuTfwmWjRPU2d/5K3c1Lpk+yCPsz8zJanVHeXM+GBY4gXoluLXhKMlYi
d1Kuj1eFHVJOpoNUH1CaDhZwY5GV5ChyzNoMqK+FvcxpPk+5T2S9keU/ROX6
9z5LIue8rCi3AQEQ5xIKf5YDeuojwn/uJ5FB6zzvWA+hwUf8SnsmztNbmmRa
CBgzEFt+m5IerkpVUN3K/NDSuJhe82uyylUvZ/PHDPeCw00ZveKEwPhauuNc
rBXaHF16+LQfpV+wS4c5XCYr3A9tt8TLAYyx6+K0u82jsOP2zTMfY92jGXxn
fZGhcVIHt1r7s9Z6Go7EwpDOGFMOFum/bzgrTrF2C/938F5yvYrF4fOkRuip
jUk3GxIV2wAgIFuWMooCDAUEKAxDd9P3vhcIV6TBAyRrLoA9DhJggAUXgIXt
13QPvGmrs0BOYabdCBVsgScyjHLqY4aONFINJmrOkgCHnRGhzVmcBIELgNVB
QznbvUn74KPGoYUy9qWEZeU+OefS8MXGS6hIUamNQ2JaLRNsNVAeUrfgHihi
uhFxv5LJrXvjsjUbVd8+7kXaSRGeJ5va+gk4+QW1ZKlTHRd3no36dle53UiF
TP20HY45ZKMQrWkOHBviK47y+b7W12NQFIBxr4jD9oaWRlh1qrBQSV/tGl9s
HBYo0fOnFmDbXzvRgEYEdS2BliMnZl2rgAFIT5NwMHFWujNSiFcCNjjDqgKA
6qNPauPQLbkOoVV+/pwwk073H1gySpGVVQvwkw1O2LEHWcrZqHroq1bVgUwP
J4Yh+3lV532LirOLfzxvzMXfdbSvPEL2H5/ZPb/tX1/DYoD9ZN0C+Z74YknI
3XWXR+w/0uZad88RGmJ7pOOQ3/EOTw70VUcary8OQwbCBJgr/ORbEqooxDxW
9YBBFFBoPkswuCJ6BHJufwDvAzTtB2FeYv3YMSvCtyqRO5yDzoZJmuywTM+h
Kio+Lf05iG58+SudKlDwKPIY36wQfoL1npi2RPsBnRk+QONTEKxnpsSHIOm0
7i2ZMcFC25fETcuEuNcGVRA4wYvorWXzEjiYmO0Z759OB5GoyJ0egJ4KN6l5
Wc1EaokH9DHcvi517D+tFE9I+kjo66IBG74dzz/Ww2maZWRqXNcC/7Hq29SF
LtDdahbOxdQ2vJCTq0qALahPRCNalZho+urvubx2mlfiBc24nN523znvXAd/
F/HrgjF4xBiG1Y44Bw1Pnjiopi2BTZYQEHtFbhiAcv80vRn98NrwDC5tGJ05
7nbGW0ZhD7N5b7jvidoFsW3MRO96IRxO6ReQ3JdLfHq2dyeW1oz7HDzC80eF
E2wlO9qPcX37qVodftEAmEvULW+epOkyDG0VDDYuqdzW0/TGg74gyPi7OjYH
JGjk+lsp6yD377e5EDKn5OOldPNMi+PT+/2mKxjbgy5bPeDasdUg4Uf7pIr2
D0WzoY0K2+rnplIdBdZ7Ec1iYcRIxdibRpn4a7BWPyXSgeeEIUsqcRwevkjr
5X9AQRS63f8Vt8IN7d6uspAAoWLJW0YyTH5lU7wvDl81mojUSAEIQp6BXeHQ
EVooMbKbfAuOKtquvPFn33hTr3k+JEnFZ8anpUva/mo0SCEKRimo7FpMxqJs
g3QNx91iUKULpTvoHFEZggluDLjMUzhLdZy+pp0B3Y3mjNtQNHDD0/7HK1dF
5zHil6k3Zq6laE1UjV0tjpphPsiadCwL7oxxDuY8XlyvHjM1cYRi9mTevdWn
SZawoGNDRFRGixgZ+bCdvTETW6kmyPKAiIFARYEUM2pQZXxaA8X9FvHFH6FS
7A+phX+z6hCAB4yJlLXaX2Z0nSLIzm3nl3M/lyD1zQ9jGP3DUG4jHfISaJ4O
z3Nz7gnfVP+zPjqo4he9UnW1LwQbDXWcH88POtBq5enis9GJ+a8lZaF+pd4q
dLWzBZZbAPT4KWI790fc6IEj1+bCRRDafrmU5EOfotQmf2UMtGrDo880PVhc
PhobyhVzwEtIKKcKzhJKQ4elGY6AysJlPpffnvMieKmGY6Uwjwc+Q0qveg7T
aX+/jC7lq20eSas7PNKJmwKvWL+Ag6dXOaOKv3diikOqS+KOQgwWvm8I+hMo
dycvggB47LFGa/qJaM/LwIRUfxELeaO9Xt6qbdXuIhcIpYRpnHKbuYQPla2b
5ynj76yaQAsbwO3OlYx28aHFS9Ellq/JnGfRZMyjuvL/e2gs7CaFmp9ZcIqR
XW7W88xhvxBUZ0CvGKBK3BSFmV1L+ZPH3iJI339Hcma4Ahc5zxeZHKnRX4Kr
cJdaEpIzSfnV0rgLUsX9rq5pgr0eRL/5UD8u5VlLixk48QKo99AUzW7oCvQL
eTbSULNjTZwoDJO5A9RFVjdUYMVAhmqLXgbz+crTBOHsOefYA/FW5Yw57M+k
Yao2IR+kzvg5nvZPMqH4X1EZVN7aoKOej6HbD9S31jlmmtmVpnq79H75YnDG
pMwEOOWIKIbdq+/oQBj+R5+N5PADSgDebaYC5Kr3D0+ayb4z0zru6+3e+dJl
kmlHc1ZxmgiMRKZOjZVtwpyZTOMJeAfPuyoc+53XKigbLxCSnRE9oX2AYNOG
6i2jkdAEN1aiTFLhPyL0CJkH+w6Rkw+iozHuYEPM0ZNNVjkjzQjRKz8jexfS
VnAhBUrPRUmVyWK/bgpWWCnXpWmMk1Oi9C0AFexB3NQbts+oa6R179CBkk2L
A6swv5qskWayxsZHuHcN03fEeafIHjnmN027auzKfO2AFwLUcQ6vC+D4ZOVV
phZlWicOqor8OEtm3nCA52rrxgV2c68QazzmEA7KMPBvj/0qGh8mqrq7biPe
9QomZAwiDqjUujmp4r8S+bmyI7A5AJ72QqgieAD5Sozh+sJHtVkA35kDk53F
U3xpH+yePVh4q6IAIKjUHWTOs4fLSBymfOD43VUu1/rY8OAWT29YmgRYBj0Q
HwE/hv+DQtZ7Bu1c/LHtCuSe+Rdyc+K3GXxq6TFmkXjriidmhSN1xjlkLzb6
ckDiklBCAlZZZ5kvdOcZ7KvpI5LOlaqOZc+uCqmgnFwogSvtNwjRh6Txh8UK
Pok7Rsb7cB65nkFDoM1SlX7h6SexIYd0r6qkQf+8icG/51ULD9NQHVKMIzqT
b4lbazW3JeloqzPm9v25PKsSYVwbbKvAA4sleZQN8kU1EYNOlPQHwx5eOUkH
q6tSooNsr1o7G/P7ztlLIb7jtI+z8kX86NqFjHSX+lFsfxKSQqMsmQqsvy1M
N4amTfk8zhxQvwKVcx7F8wY08sZunT4F3lrIx2PbRI3MjLdlH7qDI8SqSgEU
oo2YLPrKmQbxG/I8yPUP4TblXuJlWXy0NC5CkdrcRq5NBYa7evg3NMhem/IH
yAH5fAHwBSJ9Th/icIpFp0Ve7X4zBqeMBSAmWH58xHzb6jDbz3vpIW0Jj/wx
jTvqCyRfRo3fhGiUzxdt/vdUaqtOzylD9JwRaaPEVrNZxcdegOXVmUQk5eC0
76TX+bJLOZmu9e7maK2ZJr22ju2qYMO8UPrfEH8SFIcV4Ms7CndtbmiUtD9Q
XR3htiLK8LiY1PEbteGha3lxc7JlNiK0EDrSk6rqM5XwFoHxdxeJW54CRj7X
wr4WESV1nUpcdyr6J/+yXwGEE5um28d+smpm7f5Shbe2XcfN2ziQ2/SKgrLV
MM7Zp/WTr4dsrRSw1TYQCsPlo7EPeqBgrlpYxz99T6Q2B+J16x4MGP02m59X
OmiUnqWw5cUsm75Wack2A7YRfsAH6q68Wd6fJbQsgIOQSRMHSqg1fgLJFzvt
d+eijqhh1Q4yG8Llqe2ju/mT+aa2EKrYekx4Rk/D1ert5pMW4eZ+KbGcHLSM
iSud0WYy65xtbZlmeu+r9bFjePFRNiSW8volLMn+soUWSncBAPB+MPbVc8Q8
oDYWyubYojHDYj3KrdgNGdYUcBfpZPmQhdnaKTRztjcG1ed6sVDbFavAl9bs
G0NkvCGky0RcZIYBVjRoe2aORFuMzz6I0GfrRkllx2WERxgtnvU51FEvdYMl
+HKv9c4GwtwBmtc8XSqYg05mclrqRsBOJf9imP+t187AF2AUuCRDHddjXVbv
/GNaMXa4REBUlpwTyaQyXQiZ0sjk5/IaA0WNbu9ev8byB9iY0cUNnfZuOvEx
gvBd8dcjACKl6PySG1tAHPrTrPKunToDiMW6SDIH1DCRxavfAkPB+c4GWJqM
96Q4MIoF10/rC6q3YCs4qeDd0RnUbLs8cSuxMFcp41UpJwe/r6qhJ3r/elci
jBdcxlpNZoc3+Wo1C9BK1NMGThK3F4kUdz4CwhzN3cgV9icpnC6jyhB5qlLW
Xq6EwCP8Vj84aiUhv2Ar8XnrQPGyNYdhK76Tpq0Gw6ijYTbi3eBFucbKop/L
ffrXGgok3qXAAYRssyrpn9vS8j96Iq5srvaa49yAmMQjlmT905y9A1ZSQANK
aZt0OMfzsLUVXd8eloE9jWNplavnvoTLNXq1IPBVbfJCgau2hrY2igf3m8HC
ZnnM/Sy94/kvA/M1yZeUQUeFbhgmYMVMGV8KoRNGc/rcdbe0tQrz1EvoyPt0
OKKaF6QvtptbaXfGpaqH0VE6EzxVMQb2OEefkInTnX8r53h8vnutucZMw2Ev
jL8fWuzXy82f6C2NxsoNo6lzkb89kudmDnjzWsP9q6ajdAOl92OUQPCQbiNM
9dlJzD5guEK1RjbJb6jPw2oFdVpE9x33TFzURjM1VgCMMiidsV7M+2ebfYcB
2p182XJmM/ZeCHnLSMIw1J1J2BG228R/5j1KONVquOm5jm3jm9uuKsWWek9R
4UmxgywT9KSDpSdOof3Y4kEP4rJUjueOXk6OkF/mBbCVlRHbwNhvesKbhF53
Gc6Zr+tQHgr/ah8atS8CIF2A944wTodm6DL4p89nRc5AKwVOFLTs4hfZsjs4
p0Stf22z6sG1Hg1P4x7QoQ+e2J6dFi7voRCPwl9RYgvjxHBnrx6yuXMAXpUg
NU/V1zcK2/o50ltif2XMtLumk7WyPsYrEUNxV/Qg6XkK9gBQPlYZrwiS17f2
cd/zSI3ExYtQbWsYd2+/BBM9aPflUvoHYrZ166KKJuwkqlC7oVI0vjKu2cdw
UMGOy6jxcLGHJ2nTDchDxt4NFzBKq2Z+RQ9n7367BNV64KCbpI+/9rEJkjnE
aZ0cfuU5np2T6uZCIJnmb4vQXRNAs96O++bvrFCxjF/Uh73SyKItfWFnkzHB
0QMSKLSCw7mFxlWS/cFEFbXr6N33z9bsAQEPbVqmMqjqTUXh/ew17bvSHwKC
L72fKRIih0WiDTgRTNUkNw0UH45GWQC/ZAewiUkSbqaHmqnpR/uKqQ69NIRT
oUrQp8gFnm33aSX5Q7vwfwtcxCtZdfNYYQ/95N95T5oYOJWN0KvWDoi4245k
hpCWIaO4NcGE4vU1KIt5cG2EarEcFDBH2/OnXO9i+lDAuFMNPBS0QPlYOkzE
zeI/e5Aa6+A9xjKX2Iv+NGKQUDTGdrv7pA8TTSOsazpGjmeZZyhNGLXu6LGx
DOBnxISWWP7/79+k9KU+XdYKb2boA1XW6GVe98hyRYY9mm29A3Pn5EpYnI1u
yRZiJSdZmwpS86DeRoekfpfVEt2H4vjVr7SCQBFCkHyqnaEUBWrl9uZe4T0e
IYWA1Au0D6cE+SmcTCEVMYWZYht6JGDTGO9aQQLL/Okq4CiKAxukA3MkBcGD
JuKEzdyPL9aNcZWYtgWmcr8lbfGff+N6ADyvzesIOWozCpE9wKy702kBOp3s
erAHuJjhro8RD9Ky9HFJ5+ou9/NLfPDd7hbXFGTQPUwCcEFiYX+/DEMamtnK
JYhZtthcZ5tXCJryKRhMhL7kODg+OfdyfRMEwWys7CZX9nsjcvfzJoJc9Gb9
GH2HTEZOQH5KiOFXbvRfR5WXU/6+oIlum6qozkgjsbXaXhhbas/HX7vvINvv
ekjtw7TEAHMQjn3AA1HsbIeVkUi4Ly9swSprf7JSa5C7+vocrcvENeHOQ6Xb
glQ+myEXH4xYgjkDuXo1+mB15C3Z79TWSoDXsJHBwfdm0UzwO/SBFfIRsXSQ
6QwezH/SkwDoNThYSMz0xAz17rsNa+rRVRFkmbp/e/C++Sw7HVYlv6LV7GgY
BUHBhm6TomwbPNmXaVvUZ6/oKKKx33IB1D+zMPhBDpwHRxvYSUWjjqwxeuP4
QxmHcjglcnbWg3xn/TdweElNJWZWYOKgrvdzXjlHWeLZiS8suQ/CDNqXPhr4
StCWy71MQsPcC5Y0dwL4R04fGKXlqJbHgerp6EzNyBDGOUsphjrEpP9QqWyL
yQoAr579mpaM6BO/OpX4aPAvImlNIINpNHUUDb89jr9RNJ71IMZOwLW56/vw
vyqNdIG7T/5SN4+lsdZrRLIsRbg/pkf4TP/IiqqLMlqvGVX1nVDSenGlLwKT
m/NDjbHNANrNsLNphAC0yjOxBPa4WiRw0dLAptNqxRaDHRmSphR5DdkoqpLB
ToiaCe/mSZ6imw4XtRD7U4wvxZOceq9+vaA7cv/sjMbmrU2E3Zc0G9E7qlja
FmN6Hv8s68SnWVMvl0eSJKL+VAm1j3iVJYx07PF3ADL54dA5l62xMtVjnCT8
W8zJjMN13eC8gMCCihi3bsf+VSd7J8w921w8A/OfZKp9ZXIchLbbLww5BlS6
Ciw3Eza3vJPlq7ndUVw6fyETKmCZe6gwHeZ/IKL1Sjrmdn1iyLq0fthav8fY
F9Ckn7hwENOIVgY90d6UC7O7p2Fz2AUDFRTABAqE1rxkghB6zj9Hn2wzsykx
jXqHmmhh3YXmkx4EcXOUDXnD1p40puEXNTirVmZYo6PVE/l4XKn+yZaMKHt4
n9lbVh3FjFapTEruhlHXqyNRLy1HvLukC5ro3SQbz2rWjpSJ5AZnfgY3ZV6L
hvxAIM8pqS2ZfTZAyx4HRyVbS2Clckiu2LdRFFFvEST9bhN3t2QwE01+DOeC
WuaBr1NGSb9BFBl7f/wuyjgS3KcgnI4gelEDq7s3zfuPYBMTh+xqlvwHfnO4
cqU/2xx5U3Bz1KuyUovprMjsaAA8jzxqeRuIqt6FW/p1+y5dSu0flLba8zya
bc/aQPiT6TX8UWZY+aQ6ioN69/Kx07QeQ/+bOmrhGJH0+JtU4WqZCb0boz6S
lJpUMKnrQMtMPYm5FHxFSiIM07dlK3h4zadQYI5ttHuHRMjIKHUiBtu8FwWU
qL2NtFWDjRwz0FkASln2Z/kQIpCoqodHX91lV68HaV7tkT/fI3xfTSnR1rmm
BXonFflIF/LeTrg6hrNgWzK9Pnpq4YvvKsUlHTm8owrrTvuwlIt1vqTijfpX
lofPV0uNnqX4esyT1GCiivEZR2VyWDn1Aobc9AXSkm6xloVDRqZTVXa+Yf6q
cgRzVeFCb5HCkvMxfazdaig+/ZBXEc0kEiMDcdPEzXZ1UBw2QRDQFOAtYiLS
Ev01jx2Zj8FIYxJvObfMjR9DIcVrWhzIBxkCarErHnCODW8xVbNjSnQ3RaX/
vdFrSXyMvhWaC0ubbxcSv3PPsY9xdKOhopSumdWHgZAvv5kQJvOH1VpeuOUT
UE+zmr5czvhyAjLQqC0pqkKr4qS0LjLIsI/WtEQG47vy7ptRpktKyQWW7K9X
fDe6rBIRz2wO+gsgfc8YxRjyHpwvPBufO2t6OazO8k5NY5kEXqm0b3yNjXQw
3IIyD7cFGdYdGUmcaNrrRIJpOOtpTaaovHXydtTTyKpa3rZZ76EF79zu8MR5
oCN8w+JdfJLsdxFnI/0K6jOSEIUcYcJd5ATNKhvHgqX3qIPdvr7DCyO+OncI
SL1vVc9oszJWRciPtIAvHz5ZtIkFuCNMfBFvuhMKLaM4RBp9C97+nbyAJMKs
GweGP4rgp2n6x/pylYw+0MKmcU8DTjavjOl0noOFHFToxsNzqinrs330NVZe
UzpQkb9wncicLxtEpcWDYziHsTN54nOgSpIdV7FZvYqZ09TLaBUNBOOwB1zY
+GoF+u5/RfAQfRs3RmjycpgZD2dHlqIyJABA97uF641XKu6QTTcGuwdvuigD
dixqaBBKKLkDQ7/pDWy6p9bvqkyuU9BnnukdVrQoEmJ65vjlfcC18CqD/zu3
kh030gmTnmjDJHfBdX0Fg8+8I4fLJAoeAfy6F3UCiSEcHInB3EEB00eQh8Qp
JcnvHhKsm0BWwXUcXYpMxzB2+o1j6J5D0CtCVdACugDERLs6u9PB29x/IBS4
NshDMj+1QRcNadHcgXZoalCR8u06uVLFKIvmlJhsDTWhHZS/rgoneNiZwg9l
ZxdnZDnf3j8t3GsQUCFi7KYUVmnhrR+qpblSciyk8dkqOAdkHo81eCSyy04Y
9DgVR4YdwsqDYBhNFWZM+pHmsT6eH8q3VvwJzzE4hp16JreQjib8xgUFmdnQ
WGaKGODspb16F7wBai0vZyr3k8sy0ZBciweFz8bV3TVfNu+lMsG5hIhnRkPg
D2wiheK6OXir4875HM+dOloZAmVaoxzJvJfbOv94wohvlT8BTy71dg3WSCm0
j0yXnBmghbhJTD+2ZjiSPIpfGw+UjdTuIgARa+hIYSnjJTR9aI4B0ZB/TsBk
h4A3oIBtD27KCvW/C1lceCk6SzuDwR4Scg6etL6P4OK2TQp37UQnTTsIRkNd
Fs2H9cFvT0FVucWe0wZW4it+2jizhVzREUJpxpQeQvgt80TvtTnn4+cnpKrG
9fm/Flh7IphL+iGe51q90fSHyyYyK4oZMEL7KgifWCOoyz91uvhtl+NKjvjT
wWnI2PzVMWeQywbV5UPBcMQ75eBpIuDIok53CdX5RM+6Bc/+iap3EvUC9L7R
KwRxLuXbzgamcaqlSYJH9SSfXiT5zEUywbwCwHzHsWYH08HZ49OMb3+dr2jc
PuWcfUiwqXKqoKvuXP1nOTJViz8Gxvm0Ys0mJniADCV9Lq2SFbakZOeuvGfw
B5924m7tWW1asVUu7mWTZX/h8v5Fft8RoXU0zn1xOeB/gaJPBOd6QJn246wU
R96wg2BCyeGj8r1Mrd4oO5jrRr5EwhUm+eQZSM1YAR5Cwi4N7ootbGqYlE1h
TvY/Rcoi99Asa1i3cKKd6/dl37vxWibLSywBCIV5DmfzizfLe2e7DCO8/ugG
/ZjG7649FLljEGgDvE0a4fW5QdWGDgCmecajKOpdlbcjkCqOKvlxWbRNooWw
QoRWyiUJ/Y+bMVuLPGtd+hNt7fdJEPUreJ8Swxsjif49RoaDgEvRtTw9tLw7
103yKRpLUIQj+dMatJSvm6kzSf8OyC5znv1XSPmUdCeglM57CKRl1TDxP8tC
4RfjbsBIfGHrRqdX2BKk3+fmPCwGVXkea+ESDKkDrTXjDQL7g5JVLLkOjwdl
9udiWMRGik7ZqQhozyr2gxvRpZ2jaESnjT3i9eFrde99pLMrdAQGMKAqZ1y4
9na+fzfDNx1Xl1Os7C3FiJwzPSypKCs7wWFjVq+KAq/4Gmn5KNG3mFPG+3ZS
32q8hqv6/bY3grUEsXgKqiK1Y8yP3YT6LQVxHARmkaz6zw5984oYzzXLI+SU
7Lt90iiCwQGnt5NWRnreldSrveokaTllHvCZa+eeUBwUGErPV3t/Ne2LDArE
rqnZlH/BlUxzuLnYYTRNCAcO0CvX5rgpQUibb4yGFWVB11FyYNSDBAi5sxvE
eJpxMDSHoVA8qGDLH+y4oPRMB29gS2jQzZIE0gAPRvcv1M51H4xZKLKArnyI
5V0zVE/9Vb6G4EEYovhns/CvlBqqg107/gUHBOutJ8mcqsT3NLJn375QgA9f
gSVGClwIF9oxSNVEfY11bLkQfpyr0/4dRTXZfdXnDmNTh+M0N6Yaph58QFDR
89uUKExngOYuMz//1sjt5ckpm7ZvvXbbFBwNZ6/i+ZEmgGmFpxoIm0BsGYQn
X4rPnzw2MW3lMgSwy8Kyfaz1/D3KjD/nAYLq9pbQrPb48BwJqTsRln79nICW
D1NO+6QK+hHMInnDcyGtt6t9/NNUDWd0M9ds+fq8ZjqdK7tHkOSbqKxLqRBd
/vhPmBSTQ2dWhnoHwRk5QTyVUdYyMZLFAAtkd/SQbp4IYppM50y9Lq9KkLRr
FzWwfR3vdXgBAIzsCVKxDfPDdFrr3qIh5J5MyQs0EDoTh5xywcvl61kiKUdy
KrOkjbapSypDrBsKVJ1bUj4HAAsp98wgt/AJWU4wmlnJyQ6PKyJp4+hRs6ap
XYX7nqadX+bqiEQ6jOdszH3y0Gq7TTGykfK8NbpdLwN/juyP1c3Y/yhXkLbt
6pB78368nt1ZCt7PjjgY2+pt+kOneCE+rQObCVi5gXhLeeM1cPLkg9wKrOLx
cS2hokydge7Oe57tLyx1QSFk0eHNVQuosedJdjYbQcJbCcgKbxXRUXnYfvz7
EX6Z0tCa1SVyMIS2GMYH2tlVdOp01Gptt5NsITCTxdsl1MWdusM69llXXEGu
33akAo8Yp7MaDOzOrYzWea7yTJNxLN4zY94ldCPM0/4fhZZ9nmokPhIUboB6
9L8B5ixpg9GACljJ8j5qU+jc4M9ffU6AClwxjXJJevvJa4H0iqNBblHUgFJp
lfTqz9SkRG2m+aqWiRoZIhV7w7Hqy+WqxpFu0T9Ud4lm+JTzOmNVWde1w+wT
ZK5GTpkqC/iReqHLJetlR/BeWOZAXf4eHuT1mB11kuV/mYXiKFt2EgGJ76Vw
SOMaPmgeDejzoJ/qhoHCqoDGTwGOS6TF4X+vMNiU8HU+IaOWNiyDXV1SBhyB
srz5HVKp6Zg69qYcuf/z1RorE/LnNnDba2AvWh728+zIE5281dURN5ZNb7/I
FEsHRnjNVPzpj6N0pRL2+AYQHL7I9C1HNcx0+eoCX3QtXtIHd6Y6ZZc92kco
W2qy97MQ+jrFdK5S1cZ8iBraODMogoBRC+b8As/e8rnUQ79/vBeuUPPW/C18
mjOpXe1XhgqIqwanK3E5istK5Dz+ycXkiMUHboanjAZCGmhLWf0dlFBgLmbe
vE6bQS8jVkgp5lOclq53Y9hAT7+ch/JJTrkaGZUDYOHBemMV1pkVTAi0Kvlb
tCCSo6pNtpOGH0ukClCtrqVbfwFXuK/RC2XWeNRKo1+UP/VezZW/+LBb2KiR
9sOklfcf2OZLQiNgbNdwi4p4OEXJ7z/WP+5tMCSsCXt814sTWmRMUYK6mE1C
Bfs7t37T2f9+wP5tpZmGUvAfkE8cBHzlrH9GEIVlNrwX90OEI85oj4RDpw75
K59Ic+o91xCUnvI/F3pIjduYEIQLeLpn0xQFsjh/O0vy0BDo/1/dG1KlsRiQ
DllqGBNaBT1VwW2h6NyaPSJZY+IXwU8TzWp/rRwl+aHzXnKufMCpOwF83DfY
vpHbYtOoBltWv0TAA+6YuulSYV8oUJ9zaX/mkVI+eDBvWYZL3bw+caf4xOGJ
8Yjs5CVux6mXf9oky4FjdRGpHeaOc68NY5XjajjR9rhVFPzWBrXoo1xcj458
bwGYkQ1iCckQ/6SjF74wGEFiuJiM73dlFpTwjV97eEzXwFcrNvMEeCgleTB5
i7hCSjcvbP3Lr6ckWp5NKqhrx32p9GIrriMUm/sUZtvOK4QS56e95a+1EOR/
l2mbEtR4OWyxQrdz7TzOe1ESpBHJZH78M1slN9ZqWdu8P0vnejyjf2LRkPaI
dBjjusm4B5W6XCehzI3mZ0U/9CE6B1JlZc0vZg1YzqcjUAQ3ocqiyqTY4LND
QKs0zp91VqVDllzmlZq4Tt8H+/Um9Si+VRW5ok5N2esVkKd8/mfSFA3PA3iS
1VI3VOZyq+7gknl72al7n9atwplklGXXF+m4owd7eolnaMEqQ2QFpbhWvXrW
t1Ls2rh+p/2loF9YISWMQMC9IojltFod2+VbwFHq/YHbf2wJ+jhG5/PUMkKm
f1AYDcATvnhpFE65ogUAVfyzWqe0dkPlIbozTQOqDGvLffkS888RHp7KrhPU
C6pBbZIZfzR4veh6VU+/hRoMNTKA54QxdTFEo6oT5SISLOX/e8b4kAGXErqt
dBCaY1uXIQ/hoQK3DUNbXmC8JKjBl9cF5Ltv5ZyUqJDaao3H12OATXov79eQ
IYmlGNF/8oyS9nc1eWJXqrf2dHliSYZgisL2I/cOYHlYsBRtgdKmkckia7Cr
8SQA2bfZMUGnyMcHY3BaWgD2LffmtqNOLmjyI80xVSYSxs+vt2XB+F3CT5wx
71SKHSC7R8y/kQv+CoS3ZJaHbH9gxdWDb6hI1Z4x0uTuQIEwSfHhtfyZQGWz
vOexSRu2yWMIrNTJaZY8OdGeYU5THytRRTYNjUcbZw50cp0PTAJjGUawPx16
231iL+yszNjoky1EiNpt9WunqWTg1+HKKQwosaDQ+4OvI+cSVszEv5NjNo3I
+QmESCP6O0U3r8NIHicqwPv5jW05kFhr2VtF16IG7O6gmm1hXoIU6xDHxLkn
KacqRyDORLYvXR+lZmXnSosMeb6p+49Ola8BdNTgKMGZKYjs3i/ZPpCeu5Sl
s6+yp64rYAKPkgr2RQb7j72x9X9rmp2xnghPQO4GF8ZPGcIOzyMh6FmBr+xV
PVlcfQLgv9mTBReOFK0D2l/YKDcK0gq9AY+EsEb36PIk3ULIMpg0B7mCq4lq
b+2a4fZ0XZz1CYFKl+U4AczeqqvTcUwEGw9QmkM9/7++FNZvQNZ/YZaKSNr6
IBoNs+pp5y8reeoR2/UjSJ6mmdEcnVE/2bHzFcrcd2jyzLK2OzdhC+5pKzE2
sSxHpRNKwC7JTHCSnLMil/as2nasOGA+eyaMdvSx+BNxNROP3WbKb7k/1DRf
Xfuh+nqwuYlRgCLMFBYBeR8FJlFomp076QDmTw9OIG7vuxvlOU5sRthAz2q9
4Ywwd2zw3co3RBlV4g62PNwyjn8mdLbNa4UJ0j7Y2HEQRrNM+AUjdJhKj8hP
xGiscV3ijbtMIxeT1DAgBSKZqxywlblYeDhdsdVuj5F1X13Ofz8K2UtvKvCT
WuR/YlNH7nc6JfrleNZU4gi5UEB1VSFOF5X7gVuJbSVRqkX0HeMXMhS6pcqY
3ViiIYWVsT87ctJekXxs58fh9ioN7l+3XAtHIVIhN7Q52cSpP4LWAK3dbmYC
iLVTo6rZwNIO5x7ACObfHJWL+N79/FPncle7bqf+5GPMH9HJdVQCmZ2iTMN8
vf0AccaB+CTiQEOw9Xbz6o3UK71Z3UCkogUj/WtkMzIE0KW1B2kd7sbvyhO/
t8NOpHg05w/uCuIS2UeDikqIb1jGhfDbV8r7wB9dzGuSqw7uiXaGCAYVO3nj
CMKhdjvFZCdS35Y1TDBzmWF1hmsMCXzviL1zfFAys+8nwWUFYm2txhCHkPxH
FCCe2hRdrbjBjWt82pZ4E//zjWaAZhxOJU8sIIMlhjn0bc2MuH32YFywzSNx
k/JBV6nEeZzoiSGEVMZvy4LkXE9TI6R4h0AP5/HqXIuAOrbAiobVv31NpeKo
tCZwPykEu5ZxTHiMNTb8GGFyD9llaX2igDPA0AcG3dAuR6JeKzHAMBwJe2AW
U4Jy/2KHaDBLw6iswwZhsg6nOKGr80+mkjgPL+4mabSqYCsddvoLfv9IFVLD
4Zl6h0oHZZ0YEXMj3+bwj838QktsUtaRaA3ciR6+bTz/Zh44u5Irk9Ia6OBO
eCNm13lNPm3gsMjCpHS1PozMo8ThghdGh0yfqvbvtnQDE7AHz3vUHEwH3kAl
SwlvbPiPSlQ8/c8oIWor3Nq+ErIq/bI/fl1lboPQr2pes5o1e0GBUYP8D3VY
7zGv1JL0tWr5245+NoCiUYHzxwO5hTyLtsA7Sr73gV/3qP7vj2WCk8Fh1RQG
SICCnfJok45asIdsSzzl7QAVMyfoifmMoi8d51VFHtcZaWAD6Mv3mfEAtUco
9Xpn7Le0Gm1rUvTf79h5Fx3++At+tLD/UuB16aheoQXEtS5VD+9qwZuluvOy
tDH8SlaTJxQpPm88r9U0fI96NOA7fuHArw3J5tBtDzVpy5NegEig4VXIXylD
m7rnfLNqJ0iJEPpWbiIW6lbBE5g14wlPycSHD2miupWVbTuOMffG9ClhB/ui
JKrYD6dd0hZlEdFiBeCgCpkKrK3p+CkV8cG5MgsBE7+JIZoz2ohxXFVoIcNj
IZsI+rq5oC9dj0GYro6tR+AyMDNu53e9mpgY1cvrkiowAphm1w9H/GE6/bwE
FaMQmuhV2OVmLyx+Jnd8joJsJJ2MqXmsEsMz6W7LGtJVGRRWRjKQPcHY709c
Gq4beHQpz7r/YAAqNFHCkqWtj/eYmxbQj6CsdfR8SERukzG15gnVM6A5Fugi
EEgKr4IQy7vZ5wcvy4L1AEW9xh2HJBaQ3bJp5/RF6LJLYQfaWStN2bfsY4KL
MTqfWXDIBkqb2y0+mE9jn5naGhYG2w27Xp5dpRBR6FTIWxhZv1A4FiE1GP35
/e+UuAl1oC8CoBZe4zwHBN3EgTnpzTpw6g6AZPX68SBblyhy/hYT4NYuezEy
0JjoM5O1QaROYFHrHKrFk3i0rPPpj43nzl9QJ5tb0QFxwYBXwBtsFxAWsNNp
R8fMTR7xlZP6DN/+jd1MP07Q62Vg/St+ZtEFushDJmELp0f3VMUP5D16xvpO
J4eNchq90EzZLrhsik8GRfQRhjc+jAmBQulFbM9RpMDkQ/edf1fmgubv9gtu
bBCafwRmjYbLiH2Z/fRuvG60uuacB2DXojKwajasOyfhT8IbJC7oM8PTouzm
mmg6xnufEr+H3HehEvUXH84Q2H+oZkEi6CdEQXWXC+y1o7PuKiNjPQZXCqrq
fEyR7sJPxQ1zDghLt1J4QwKszg8MuKshETYd+p1q4jJqUU0EJBullhLdoTYq
HUxOWfWYQw5sOBFRGSdoUijtik+cDqWNhRlL98gUNq5scb35FIEYIDQyY5uA
L3/YHsO7jA4GQUEuYvQYUKkbDE7RA5NZZ+6c75ue3185+g+RyD75mV3JKR6V
BVUwFd96q/UDsSjF07mEU8WP1H8OHMqG9x2dYCjjqr/UUhcwg4QI42+SgLdC
+Yb732buKJJuAPja5mmIusPlZTTRgT+TbOsXhEmjXI7JL1j4NI6EWDTuzNlJ
q5xhs8ROkpX0NUK4FBgvzIeC0EP9SaJ1qOMokPLCwFVhWaj7igJs5umZiSsw
kUVA+d0I9VeMMssSgEvHx78CKVNlBovipJnWR0FKNB6kwxV+HnKH+OQ/9Sc6
39fg9LvU+ZcrvTUfsty5Xx4fJlyjlaHf9splFg4jUPf2kKXcQHzkF/fszgDA
EYietp1qx1f5CohoBhoaIUYRr2xOOYIipgD4VTUZxIiIzc8Q6bnCIUMulyo1
Dc0Dqhtf1JwS8F90uuju9mL1oyjT5OPoScxfl/hbjsXH7BhvoYEh+W97RR9i
PnZLnO674DPZb6pa/kp9MzBIT+TSYqW+zhAbx68N13tAsfHFd1qh93X3F+JW
53ThJVyTzUDE6YTfJwS4by8Yf8HmV7ETLS/8BxReRvbP0ttqnDLvVx2q1jyw
sxCz6g8buGgm3ii6BLJ1h8h/ZpCyQDQmwfJPu0Pllg5I6xHpxcXoau0iAN2S
epSm8ctHJcy3R5aJvKjrajkJ/515t8nlA5mKTmpy8oiEUJWSv2kFd5EwVXjx
EEAbL6yeQ1eK1lrJ38QeUQOmBdurhxZI9g+/qoaJ9lRWAOREluwinsTAxupp
hPQnZC3sxeqTzkFIbC0JcATW/+okzou9QE2aD0cFTvTlY+QFHtuy0OD4xbH6
TX028FTYe9UvNAdaPFY0f3cLPmrY5ZtlyMsP2DYWdHJgZvI1EeyCNpzHdxgE
/YazY2747Ls1evjVMNp2hF4iKbuaU6EQLbOqxMtmfbFdA0tIwYxk7E3Hza26
Ba3Um3K6qEe6yrXjAsvDZNwJM9ELnSYNjSHdQY2BtUKGU/qiuUB4rJZgAVFy
43lwJn9NSmGJg7OjCgSdP840a4p1WGNdwNZRPSU3MCNN97SC3BhahfPjgXfn
X9fgqqfEGfnpU4PJlI6ZrD0DiAJm3QJvuNfFlfwBpoF053AFL07xVHYxOI71
Izw1VWRITQPKQsnlnU2wYX0EKZuY+66nw19bzFhKE8POM1A0otne+TMAp9jR
z1GLrNJhgvTvMCh2xLVEADIKk8iWAeDo51PCpCF2WzdtRLd5mJOCHovUa33p
+K5BsJ3+l2r0jyJ3/G1u5hNq8UWMeyCCGMA5fX6P2KdA2Snd4bDzI+SJiCqL
xHMk+KfyO1jy0AGKM3axEufS6Zdt2qdix4h3n3n4b66EBNM4y//5jJDGFEoT
ebK17qlMqS9yZi6XL51UHFLpb1P44GGpANAHd7fclrFVsYr2j9jKCAW+IsYK
vxhxppExRUfrK6f8Ft/PYXSgIvh8vBvOaxjQUgr38Zwva6jOvr3NbkzCnR/Q
qNd2mS/U2SqS1Hz5cpCj/PoNsONdElRXcrykEZN5QOiU6+iuvk/vTG07EuVC
N/hZ6t7NBQ6h1LBV6qeiEPaC0KUHc2UXvfQdZzga1wL5tMYRaZROnjt324og
kLQgvWeIujIUrqguSZb4710egnBfe5KGvE1x7QXJgAbeLs9hSa1gW4M5HHsl
5FnGRZrsUThe1Ydc2TCHbOpUb7UDqkxbLefd7Eyb+PJfN4PJRaFZ/NM+OyQ9
JkArnyOXtm+76cFCzqJzbY6HDNf5xs/bepk1oK7fboFMGXcC5SqsZgtXhBeV
w9zrn/ZAmeerrbev+8ClSomxjSfud5ChGFz0BjYRrReqqyLbnw4ad2pr7xTQ
XnR6BBvQz0mjva46WDCojBgyP1/XmT6seCcEHDOjI0BxL2nG9+WyNQxTO5rz
aR1PlsQjOuOMoto6hZ4M2XNafObbWdlazp+OvQbk2TkPw93O+uwfnDoAlkN9
3O2h5dRAHnrYlVSwbBzYjfOMQPj0cD9HWCeHmheaabuS0O+XhtcG1MnaFTNr
CP3EIfim87E1c2y94exAo+8BxGv419JumFIJOio4BxgZSASXrB4FiYijk1iM
snXM3pEMCPlVi2G/i8I3nWG7k2PvFSXdcINyfAqpM8tF0577wu+beYT3+rmE
81QMmME+/AZflCNiJnfAgMUBHA+uCkKq7yVij8bqwDb2ImKbHJesOdt2VTMZ
mLaoqVQsyukF0ZsHUHOJ55myRBtD4rvEwwlQDYxd4IW4bNA45AmzHTuyjpfM
9Gho6/nZnHfTXoZrGCDXHkg/yVFAR7WXUVDAK6EMe8QZu/cqxJSZfb7ek/F+
bhUDjm0EaM8owWWXBYBkFW9Ld4WKVO1306JKnEsEyrq69UxMXoh0FqOWAXYM
rhfx1zAxiZTeHO/Dl7wPer1Rog4TsYWLfinL3nnbPv7KLyH/oS9r17OPVbuT
K+eZcbo3o0v7bPd/j/KS+lL7hwSKamTf3YtizxHs+51lYvrxz9lg/p+0om0I
IUYD/CSBNQ697W6tINoDbRCYi4F500MAIeLfpKbZZU73oMLmGJO4hnMNV3aD
D8eAbFWjrvENjfeS1DebZNpZ7Y1laTUWCoh0MjLk4KJc00Wr2PLAG/n3tyjC
/CmyAR2+C6twCR6nvT1iUL8MhVseSHMG8cmCxc8/xzRCmYCurEq/xz+8l9LB
j/zLq7sgz1zKmzPGO0VezI8uFPuCTIHJOplhSNI8AoNj73I2JVM0xvmW/jrX
NuIGf1p/Ses4W4gAyX8XrfNxKVsjfpKnyguatyyS4DoiuA2pvclsEKIPL953
eFOYVgxg5B1cTeBRyGJYxebdFDNxXyw1QiBN4/1Vy3sOC6i5EolPbffrw7Cb
yT8goz8saEOaCN0XoEnEhByY2CXbUzSJc6rYoMm8XE/sVuonDsDRdQEPtNL+
ra+Gy8Zd/sDiAemQpIQxiE57GSp6U9nAZdLhCJ92k4NKKsjHWZB6jCWntvZB
ZoF6G530Sm5lLpeV/uRMYwmUpVKHex1cLtDRPzUI99jnPzhL38pjnD4COx9a
XMOvbaZecduDRkssja6K5AL5PtIbj5CDL8Th/qiuegBBu+WYvyHaCDWj44qJ
oIRVxS4s3YKrTYQsk0dPHizedwax8QGcanSTwMGv7J/d7R73iDBneyNt1wU7
lN817oreU65GseGC2NryShsrCn8B3+0dEAeaTcZXFU0mgu6s2LJtJtrN0jGh
/MKY3hkHNt/Er+95JakmbYu8t2MHdwhbpE1hfdoF63rASo9H37/T1J20EpRG
Vmn0Kx8sdIZCC3VTbFyqMCs6zp6QatqS8QKTJZ44FAlf1FJzW7mNayf3OOtH
rvOAdTuc4xZ/nFa1ttVtEBZaJ1ALuYWtKVQsyExK0k0o0oeLTy1IAW8uOZoF
ivriOmlLH+1FFE7oR2bUhWwODEgf8ZVTDp9Lj7VGCWwxTCPZFJ+vp2u9PNvp
W/CMmfBznJc6l3VrGnzgCVdCQIngRuZDiT5CwIgFrFRXMHt+LMLCtXurKWCo
D91Nohx9VJOLOKcTkacWWwSoiM8LxYcRra0L8XaV7IC8VZh599Vt9nWkISBi
VxN6HwY4hKwtbdssXDe4FZLh18vb8EM7IvPxdwnTf+9s5O0aY8meuzYpqq+i
8/4Glc0qiZUx6cm2xVxabnfdGMdngd5ZxC1h9RnFS6oOFJO39JgAqtMy1iYQ
KPM0XMuuVli5Q7KBAFAhMoJrYx51NMx68yvI+ZupKMirYdYDbhgTBfCEJAxO
IK0fhkD9tmDXWTTquE3tEyjFSsavnT75j2ipKByAze7nKU9sqUyjB8ZkqF7k
CiPHhWBTPtLv9RbpI6AGX6HTodWevL4Veqy3MP+7QgRFVn4MwAwoF2tCyWmY
5jB9IpMpysf9oFt+Wz0UucI0vs9uOIy9mHUqXxFzxWaci39+OpUS3pyRhPjV
VuJUDAemUbifJ0nrrFckgxn2vdQYE6CAl6i42R3ADfimIK8oVepcwofiTtxI
IfVtccfKtyXWU9tcIC58vkSJLYEY78wFf1S9D1ZSeDJ+AEul/t1f2UMakHQl
yr8cVznq6Tx259y5vS+4xIFRG5ugEah5dHEQrlQKqjCK1HcfLqDtQp7/ZQ+5
xHSKC8c1CrGsAvXBn9DKCzZvrOpYV0gYkwNw+Zw5/cQj5qtcEdhrTeKJJo1h
UPzCQxnrggyqusOFrp+9SbFNCYTY9B0gV1xQhzIkjGI9rDsFuda7RHBaec9s
p0QuxcXyduNAYufgQ5p97kuvVT9nlMmy1GotI/v/5MZEVigemHmv1dYwVVMW
VaY8I9B5fobKffryjLy7ZfPJ5Z9rjh2MWMXDlHcPAu7IO5unI3BQ4unSrwwd
BNjnuTA2PPOFCmjpfgSyZtMnS44uEBgAQEGQXrqoioqpa7VAh+2LnKoyK8bH
RWCMyIpSJ9EFq+DecFj0RPweVBVN5MkagYAkApOP2wJxzGiwD/C+yc3PCKG/
Dr87vnHlxJy1gtQglcofIVuURwXQRfzB9CfP8OFMJikWsKOWILgHuRO+hPRb
pogwA19v+zLFV9TG0cw89CLAXzCAgW8iUu0jlL+X3D2CL+v/mnENz4jvUGdg
rSs+5U8WvNPjPEqQqB6LRzj5H4i+T7zNhUpRDVdxsFWUPW/ZI2gVs+wWpGft
c1NFpVEXH4t6hvUJfM1kUGGKrA6yjMndhUNhSLYwAsJKEqvGfatJ+gExvABv
Bd/wbtUkbfq92SrSboONY4px5+NgzlfwlwRm4HwFTAn9yXy+1JyPjcIO75FR
HaxkWZNJg2u1ukb3DStmVuHXPG2VvKbn3uTa63z4CT2o7ptmWdITju4uxJwe
bJEEagHs8Cp96ZWFyUdS3NqTzL5tEhNEHmHKL2i7bmgSTxKaYMwEZY6f4IMi
V//9a/opHG8F9+bYQe8zQhaLdrTKIMKqBRHhD53mQi3Hr3cHq3mvUjGSQnvB
Q0zLv9QmmVYgYqWEUCo9FL3FMeztc6UCqYxPrysodc9t6s0ILdd1DkwYt3De
zLtp5iUkwHwoZEopv3Af5iVoo2mf4HuHspzlx8lYW82Y3S8EdbXNONgpmqiD
QfNx+aG6WbFz89jTOi5vVEFhZRd1d2xT/bJMBzV0rm0ODcGIh6pemB0S9tb/
C9IJN9rm1DVI68WL3UB/yiS5cE3iG+oOFFoNd945StiNH/ZARRNal8yRlOPV
0d+zWh1zgIjaOquzYbxbj4bLB5tAuNomF5AwwL2k3L2EqD+ZJfw8GKKISlxs
w7QjZG5/j08CZDYQ4UdNS4RmwtRQJOCYyYjvQCTNsxhUR0bC/luLUmntgrEE
7ANCADr0/YNvtyExrYwHKW6thsHg+rCiAYFGHxGkHpvSRmMn2d7kjsalTp/X
vQwQ8LwdNhP5AmUP8uXkqpgEMqQq3iDQxIoTXqnHYO7pOijNzne/rywwFJaD
z1vg+ymga5F8Y1XIa0PCBO6kNQBw0z6wFKlmW1SP71hm/q7bKcc4MbxdQJoX
uHjWZBOn2/BoSWs3z4I5jXk1cuB2pyJIeWEFEQVBTxj6iK7Byoq2Z7pgefzJ
yJwkSLcjQmjvP+9ib6whZK0JWDqSXZYPlIrhZou7ipWm0r/crarfpnbkUe5r
uKTsg2HvN2W22UfIXBkl+nFELz9azs0Uo2F+PV6tv8JxwCAuUFiGCd4Ugs3y
WKfzL9f/ReULoVmmXcZ7SC5BFWwoHpvXSOWu+UoALJGozzWht+o2f+px4buN
56vDd5j7t95B4K1Z4nIwN906nx1/g5aVCxefNOkG7HSqZbhtyqKsUsBQi2aZ
w/vZJIUUPmbAPZ4l0573R9/8J/s1sSfX1yUWKvig/sNg2gEJyqkYA1mE446B
saMOiKMBzm8ukvRj5b/UnTwDjabbm6bbtGmTd1GB5ZLgo55Nk3mmNoT7W3yZ
TqgZrn92mcRVWOL1fqvwAcJNo36gZijkZUjLeDrfJO5qCSjN9r0gp4srsayO
YHlJnHnl/y7WsTDTtnP3DFefceA0Bb1lKtjRwXv1R+vKndtYcW+kfnIPHJnz
JSPK660akcC6dB+rc3ioTvYZXN8SMqXrpce/GIIDopaFdTj4kPclzhQ097KC
f3tzmqKSkWXkOUbWH7ovOBXg30iQibN7UglMZlWCSMJU6SnbPGBx+Bi77Sri
PusBhWB6L0D2NcHZSEFaHYk8gg0gTmDY9/64Z3DIjr9UrO63sCeWYiLA+ENx
qaAEjw58K8P4dsbMFMDI32M08X9uc/HO6XrtDRWzCAm8fASHT3Kg4Z1g2lfv
o9EaZdc15YY8DWArW0HRpcz6a3M9csCfVa9z5Jy6KYQDisVRDFgtAFpfGaIL
WK5O94WpBp1nIjGTM1q3DQQrBZqMrM0YgeNWGakfzfc62p3VdP9iUTI+aRsP
ByAdNZ0Fg2dQBXlraTKPnyb0rJLx0ng9dJmoQkUxhupyjtesPt5P/I93d0GI
w1MEzn0dkf5vOiOC6Cgyx9kp3gNUX9LBxAiZVYqZkjviwR2veGrjXtNIWG3U
091SNABp1IIQPQOLTDGhGUOePphKoEL5s3KeaRwOLFR6zfAucbw4VuYrqlIa
iU4xa8YeuWLHVDvpG4IBfuxpBqfjX/FsMIeaBy6GexJGpteCbYUkLWw+wyMa
kc+wXnvjbwWHfPoZPLaPhVip+Fas9tLn62wmq3nBzlSZxYc17Kh51P1ir43X
AS8X3eZimhIVpiHJ4hVaiLdra483GDeNlQXsSeQEP/ON0BpJX51yH69yqfMK
no0CBi/0F8tTpQvYAvnvab6Xz5kzIiIK3uJbi7rcxU3pFkceN39giAn1f0XC
iteA8u74TNmi6pS/5gkLG2xUZawB6Is6P8dZTd7AqzZS4NQJqsdKTcYxAdin
95uWCEDaYV/RcnKHMryPRfnPbMf3TcumwJY5ssrIOkM34yfN95dALaKxHZio
PJ7XtPVfpR3R1DrqMH247ZaawBlUBEymDAaYIMLZOWPTZKA0BEUPdY5ZvRJ2
Fw6lPj46RfQbUCWniLA9dGblyKa81aLCc1uKYPH/BT/HFl9h5O//l8gJdarE
YJp5oRYE39mefFR+BdjS+MaXzOFmhj7fN/b/GPqFiXLb7eUtlhMztnZKFYim
yEzKb7rufqeKkFj1gtr7xGv6i7l9GK6OCcTF631CP/ZiBNznmlUL8DSXSXyO
MtL+5Z++gB2NNES6NNkV1hsESoLBwz/FgyPZx/fG9Cmg9I8lv5N5fumS3yq6
s1ubxKymeNHf3JAqnFvqNf/QHaVhq89kxpANA/8a9hPXkv4lfTZstN8Riewv
0gVMSFf/oFD7VB74LFsrMWOj7MZKzNkQIynr+eK6L/qWjUiA8L6/KGywOGtV
dSh2UCoAY62hAOIaUgHw7ARgjVlEHXJmNIm5IatWwIxgPfWP3b7bALs+QQOQ
mGvAe5leOEZ6rZAl9QvtmCc01Mpk4mgBxEyk8XAfGLJES5YtbFN08seU0SNS
hnZHylL4yyFrbprfqf1CwftLIIz9NyqBNrdPBPcA35cFElZ/WuEwPmUwc3+f
2cdQCauDZg5QMxJF9jB9ji4HqzzWciyPvmMUs8DhnPYoF/qWv7KjrPZRKRro
ekd7EAETqk4A7fAoa+5RxxouFFQH0zApriA7AK4M8a1n5zFRM/JtRdw5GXAS
y9P6XejT5jBlqTPup+VOqJmjWGKUcuF7FRdsLY8Dh4X+3xDWgQ7D2Fzan1Pc
vE66JDZyupl26E6C9NeNTdKUXoXN+jkY+kL8ejTEZCb1cI6CCwHXmif39iuu
YxRgFO51UwdgUTO4T+/RWXAGBo/AATgb0hDX2tHLiPPM3pHVaYLLbHigNeN8
qHzCBMG29u1cXijsSfh6Zjms42t3kV4UCxR/YuAW+NH+1a+Kz1C6V79eNNaF
P+YCFWU+DgL9W+lX1Fw2UMz+F6Ab7LMbE2CjBH9ywg95FwGd7/gHFvWELUlq
CMPEppc39U8w8r4fzehg7+DaV9OT++erwj/OIaDJ90HJKmjt21Cvl1yOtwqy
eCvxqEVFT4TV8xC4EINyINuXShoVOzEUqIPQxRZmU2J86Hn+XdyOwhDn8ako
JU24j3r4DXa/Y7rL6fdbf9TZakNUO7opqTR4IzuNLySBAFO/GvdLU3kqWz8C
8zBCQyiKLXngm3JWLBURHTcbnZ06QYOrbn5WbNznLfCyhhYUgRiqcS6WesmV
u8FMs8dvLDGyurDsQ6AuXgacqnHYDFtpRdJ31J9iwWt9vksEzevA1GGSInFI
RscpyqpajSIvyrWQbjg/7B2mHlvgvHVkC4CpJ3zWzcrtZGUEKnkgOp969DXI
5gqqHrQejr2gPr2rVhmTfihwEvJlK0CS5ceneE2eeyLW5gtJiDutGBFmpLWq
kUy2U/Oc5uPkVKWB7z1Oo1PINFuW9gQbWC9aeamM8OT9UegGSgZ6pOaPDyti
iO6mj1GF3wMZRO7q8pRyFo+eZDatoUp0TG/8J2klGtkITbkhSHxtLEiyzXqQ
sfhupOO5FnWT2Nf8seX4rQxudMPGSLh81K2dfSbVWX0amt3LewqWipnsOu9d
a3msivm/P35qw3H9jK4FDDGR/JlIEkVA0wJf2AL7Q9dUVtBFH5kbPZux1962
CoNAQhrAUao3/Os5qybJ1jvC9LgBaoNQF2kN9zShF9AM2wOqyYGmFXF1hpjK
I66/ZuzVzNJJClZnYb/M/EfQEJgxf8NOxW0L5acCQEGE4ywZDPV/5Fn25m1i
2YZqd8DQSUBjaFrhBW5/49ni9LATDZhCKwhcoiVDILE+dFbxtBcAXsOPWsp6
yg3hK6hmhgVEEhtQhc48+KJ4HU+KgQpuJtp3TWzedmwxmGSb5ewerJQKufzP
rUw/Ms8LKOKvWtsucVq70oPlNfOaCovJv13rVAFALipmZRGpMFjuNXJMxVoD
bERCwQa6DoTHrb/LjZsZYgNF9FCVxw0FkjaEsRPJxPjx3X030TsnqjHXauqO
jSYQ3fUjEXjiBfKXA3PdZPKZUAyyyjv+ZcGOgyc19ls6RVYSbVne6KELTLRV
JUXgNoIGK5yhhz1Pfb+JSCGAp7suWDC7WFVMcuhE+0Mi8lvl2KU+WaWyobSB
ix+y93TYU8MEtjakR5e3/xhkSUhYbcyA3nqDnSjH/+lav+ogWgRI6fdXLY9d
A+S0m3duhANh4VHOasuM7bgeLgx6iY21U/zaqeh+npbPHmPG6HbglFgLJigg
mWS3Gr7AadpZKyi8RW9pG/bRrTVdiiFfz5ihR/QFzW7eM6j98vkIutj21uOS
daBKU34Rj058fu/+aHo52JU6Wd5K1vVV906fZ8d+XbkF7omLItmr4EEbDmvi
1+77B0s9hppJHtWg13cL5bSDzT5ldq40vpx7W9jgwu1umKdLBGPgyPK80XrN
MIKm/WjeHhWXA+YBXRPRxE4BOksegKCLH6uQD4sptkRUuv3nxJVwhLpxEnC0
QDSplwHcixwFzqiNC1FsAF2745gyhgrV8ajiChBpoOEHQu7SOcrkmFZPv+zB
Yih6kwQrj8D1iomVJU+gUrMc6tYaIdcWJIrTncHnxyG/m3KtHSo+AazXXIKX
c1iuORTqE929/fmMCvPp80phP5+aWRPVXxNVkEsC3PWhC0G09WyHGtRozNo3
iWTEV2YUr+xJNTk5TgNsOF1U420fhdTkvtcY3Wu6rWzuCd72KDnkFhXigt4L
a0J0DZx28U5/L8XcHBO4XndbgRinjnhtk10pxfTEWvpdHnCV/LLYCR+8hGmx
4CymLQSnGcnGcbwgwZkyRzpwKlGLk46jxCkRsdwFzRT7dARAoEGXEaczBLFj
I/4BI3aDSkOlypPLaCmX/jZTB5IfotBH6q73UXVOBpAuY1kCq7p6Fw90Dva5
+TNjnlCJMGVF7J2FeYLffcLNuPXcaGwnJFsycpB6m8MJHuH6rq3cyP51+e/S
MxgCTgllIaDjn8yQ4wSyvrRTlY/P2c49DeUnJnqIg82BxoQPIAN3suzHgVl7
8GLUYYQ9Vl6fKJ5XfjzIu0GRsoX8P2GLPaZio1Uxll6yo88QSQYGeqSnUbUT
4+eraevI0lYPr7MXflOQRzMY0M3D7AThAAGcMom4kQOtOn74F0WL0SpYeZkh
c5A4HIIfs/5JWXcn4ubTJU8TvhVatRfiW0Brcusf4bUSjmDfi0ez/NL1ANiv
0BelImOyBqrziEkgE3DU/KA8xeMWZ3hJS91/b4qIYOkkAtllVoiK97IiuuEM
o7wybHDLvwxp5eGJmjwtC7uFK8JGekSbR6tx1JZ2uxQYj22qnxidOIU/EVuN
tsMTGF62nwQZTnY6XTU/V8ruMRHF8WzwAGOVQKSqCCsqfKDoJm21rr3k5Q6n
zSQZ0c55/jTuhHSFHYke1SFvFmEJuXSz5Qs6LPZ2RiEEL1Ef7UvdzX+nzjc6
Bq09NzhG7ciozvuxMMasLc4ZbcC0x76r5t2E1holNLbnoBxuNPl7Q0QQ6mX9
T3OABSYWEd+UhPAd31CF40CqiaWlTq6esoQU9ZaqtS//RiEo5k2n1P+Jx+cz
djYPrOF1x3E7Dr1V21x1ALun4VKoyYZSC3EKNYhOqTI+s8dnsNvtrJXbdciH
1GOq4yAMe24s57Y60juKsRLxrXiCh4JMx7Aa/SnT4mqOMS2naaZLJ07GQXbQ
fmSvPyCIQ4pmtYkGOfPNF2WEPgVREXq/9LNZKIZSxFxx1iw/YMvDGtkDd4J6
cIq2HjBOx+xg+KmIs+dqD0u5naHx6cmucHN0PvRBVGa7taffpix29OyWUixm
O3NCH5oQOuUn+GHI4/VEZmBTkIhmZevamxbQizXo9ahxoNmssohEiU4spNMq
gPECg91exVyKVglt9S6MvQaBFPMTESXJ53ThXylSy7KisJUrMEomo72R7EE3
5TFHW55DLpuwZira7MQKQVBnKW8a0elzYMlc7dels97VSAUTh+szpkanLNnj
yYj4YIiwBvWPGybgi59BjG3+rVHespczkBAFYMvSqvyVx/SCEbff1hGQs3Qf
V9ocL6r3NtPhz2YyKlIXmNxiDkrJgKFWSwluQ2wLGhqQQg4x5wDHFnmE2KYg
2HK6/OkJiiTOcWWL7+wMtZIV7IoENvOQFB2Dkp9MdINiiSYxHdfBC72ClzdS
FGqXId+QUGQJcXdNpELyNvAFNoVia/qzysxVDvt3vc7Z/dXrruJ0sKgf/vgf
wvtq9Y1qRnWtraopXuRq2AVbU/dTiHUxdKVpPgLq5tSA26NPZS2rEGMeDGrB
f1dD7rcrPrWRZgKBRYKgn2jV3qqJHmzpP3eXSPbIjq/9gTjIP07myhpMOAeg
W+CNB2bcco0TWyzX6Rhdu3NDWufuDINurkyCG3utT6HEbzY+WRqEuLrZjpZK
o7SffDBl1CV2h6tkGIFrTd53Gc4Ci3AbCo4iMTysMle6LNb+k/N1+ILv/6zM
rjLRvNbqDJd7q25cYy/L8UW6s1Cc2hGbzgxcLLBTMK0j+4XoNxW4CBkBFkf0
Umt4P2RMHEPOB6qw7trUt5jV2RulRyhdNztT47NPg+2c9nmJ9bFmLYMZ2VYP
qU0YKyxI7aLPHbYCT4PLYwzKVryGy4IqWAc1HRXBWAHZatmtQDUNggt6PoZ7
/xxlWPJG5MLN6ZiEzBwpU07E2pQFWqFYvLX8rjTj7KdNQAXca2+BEuj+HSpi
hWqjo7zbeidI51DP71tsU0fxJQP734U65yGIQsTPKjaCRLBr1XlJIOTeiMnm
TXHpI+WKUUR1x0Bzpp5XMgawt9DfB4gz+agjMeEMgr8iDlNOTCtrm9yvETe4
KN91iR7hDZpLzcmjhnGhjAJKyVpymkW6yg2P9I9hA7NdSrxmx0zO0XJuHZ4P
IOnfrOv4CLkiGGZg5uR22+om48vVepzhPlSGJbyQmn6rXTvKaXwAqPQGK3b8
jPtwVJJ24ymZXrdNoD+f3byo4XaqVjgtH8B0AwOvcuz8R+GjU7FJhSYsLrDX
7nqZblOaMl68rLS8Q8uxeKyII2EijiCy2Ksei/JjT9qNN0YwqENUONcf9rvr
70reEGrdSjFr5R2AQsv6s/2zRn9Ds+Zk8/fM4BVVnTaO7TeRJUlOvMS+23BW
ywzxyfq2pmqwL0cEXWEK6rdsXQEfBDRqbqqiEqAi41y48Z1qMPb0nM5mVTw3
O/DGCBkIefdMbUYyk0fJjmnghReqd8MihZsjyBdE91CFa61vuUEH5YL/siU5
jhIUmFvoX56Yyt48RnFANM3i+fKVBFiAUECXh/vq46fuQjZI8UO6JOdvjKCZ
gZlhxQuBTX3ktPOqT1tETrdSJZCB9SzSbGy1lxxW5y7tgfJPPM8+o7dA7eo3
byH+ukSxwXuRv2fLjMFapANqWfdBXxyxbKBU9UO8rRGRJdRiQr9ArrHBgvFk
bStbQDEkUHrt+MthBgdJmmSPYCQQdFqhQdROh1ygTeqMV9Cgh1akiSxgS77Z
aNAA9CXw1vf7trUYWrhcqzJqjlRsPO6tdY09FXIdLkLhZ8NXOFWC37hI7o99
KDk2XDb8O2egP9k4VDDT98+pxMVafDejQS4z71RxwP+zSjWa989qmsWET1GH
pUU4f1YaIoKA2vsArjKNKObPtDK1PWJD/3RuHaEPJPh+zT+V2v0OteMPte4f
pupNHlRY2TB2KydGXXLi3Y8zbi9iZ+NKAjrLFzBBUUJgDTAdYreimA5PRtza
V+S4whKn7xLDaNkOEleap14tVfYBIQ+okIQECnWGwMP/Qv+6q5Hkit/K3mpD
VjNv+bokxcACsYEuxVhySJQVx8T2P+29o3hztGMJrI1jqftql5C30NydTuXl
iYkv36hq+FG+3St1w5iOtuWFkEkg2mEjMOfKR0XnQBYTuBqHS+eGTuE8+8fi
59wxBF3KbCCteUVY5dE99qamFMYwT2swjy0eoc0iDwYmAw7ecilQ3tSaHtzK
YG7QmN7OVDKf2X8P+SwgLuha/BcwzJ4O0Qn9Z4MB1f+D49RRvfMJvV/VHics
mkNKIBwJa37xSekbn1m3MI74XMGVKjmyrJ1rXhhBku2cbfLScHRbVIyNiEow
raBi2UAw3WLH57FHxe9PNDp39+WSxV9zXOK2D5XHWyjiJFOdkomeojApXtXX
RgSsBLjG+ZdZwdzY8HRvAbBKdLcnV0an2h+ZuuaPDr69wLjmGhwGXG5ZFB7g
wGKfJ8zAe/Wxa/+GMHHVAW9P60NuQbBEeP5bMTceS1ANS9Cmzcj9Jy+BfQ4S
mpBDLsMNAoqhRuEwu+AYVLP5h5nEhcnAOK0M0AIqgeCehmm2zibl1Jmh9KJT
Ck7T05SLhkDIPR8BSwJpfps/TiBWeaP6AnlWu+fiNy0x8ZdbNvkq4o8zx5l9
Aq6025obE/aZen36myj3pRpBzILs39CYxNje2uz1BhMNSdlZAxlnXGXWsUWC
llLpqR8xNGUmdL4sHi3w6oE38S5M9biZgF1+CG7EEkZl+9YP/WZ52ZjlANrN
j8LKyp6jJIVr1NevOCC3sKG0/jRHeam3UF3VhW5iEB4q6ynfT7scuB++z8/p
dDyxVg34Kx4lXMWdZCXBBu9KCN9DCw1u+AvrwpD4bKnz/qXZ6sctfDXcjh4t
sIZ8h9wbI31RWeCq8+eRSzqwg1MRkIZbnPQEhJE0je2/1bOPXL3RonEqjN4v
3Lb+KIo2EE0npyuv6Azju8NdVYQclST/yTnu4be9uD4XesahVXyLwo2ZO6Ym
3M4YafbqaUb0WPj0oiqbq3R13dCbREKQb/Dyp/jqI21nMYDi0uG7LWn+kCIP
TQn8rkvLGrxY+D8BrPsEHyCeg6aJ1lHUsvueYeuCJozlx0+e4jGVD5+EIAqs
01MVojRMj88ziQWuhRsxlSR/IkEBoeR7g8TYLYtDM1NCsAmGYkWMc+Jy+d1x
r6uHPzLwwo04X9u2FUW73h/N/Vr/LMr42K7a6pF9v1tuzDN4lhishxJdfKTR
ZyVVXLyIdYG6C/7qkUt9Dl7lIK87N39XT74mbOPW4U/RwaoMxu/bs/OriTnQ
XDhH8+ab+1YCJwIQblEZ8obBkFVO3LWS9h2IgFYm0o33hyGplqCWjKXneYoR
XYDY29eUH2EjkiE/aEjbgYUyZDxN2l6QES6UYbkxUuSMmzHPUfJ5rgJYf0/m
Y64MijReWNMl0jr+twTK63vO2oke6aZcE9d61KBJe2NayzXzdn8sH34TJ5Qp
ON4GhM7X2lRy5iscmXxcTr+Bpxz+MwNBlYQ8qgPgrtcu8ONP0a54uwBlTcEN
BoA3kCVXOxb4vRx/7DpJtSo4NyNnFGFJNW8lm1UmuTqFWXVoMsofyniZ9GAs
jyUWMQluEV0Gm06gcnbm8xpgkCwZmxvKiJ6dC8LeOkpwnM+cf2krkg13tVdV
d4dYS5kTzWucqBdPCysOL6fWJQfPi3JZqLlbqiXNxiqwCeJGpKm7GMUlP00Z
NIJ4yDqGsAjAFZSZWtaYCTOoizf31u7V3s2Z0Kwhr0ocI4Jkl6hONTUVFB1v
A1cpmW38ip09hUTPF5e4u/P0fQMiQhFrmgN6m3FPE4ifjQ9eSIvw2ioU+Fgd
Aq5F9vMgeIgx1IQ6Ak1EIMdVSdCU4knuFoZNw7GnSOxMqdzA8aMjwvF9fATH
xvnL+VEu8Byc8snGW3arYzhNNHyHPSVFq5y55ceZ0Ic62xAi4yEvIZgln5TE
9yhvxg/aoM/8KEefwYGDnV4kXkD/h/3OxdYVmqQGpPJaARJXaAzbFqZ9Vwyo
LH5L7cewKg3QgWBX47B7lP9/DXzqsnoCGzYsFm4DKtcG2FBone5gKEEr2G+i
kmHC+zOe0OMJS1bqQUDULxmtTa2hPJTVhcoTTYJx5WZgMoBSR8uff8GWGP43
ZrIfH/+O8UDXWy85HTziyWttfwc6FVzKqo9NM4KVgSd/hsqaNdXhmXQxWTcT
uji8nMQfbmq0RrT+bPLAwD33LPCqWOY/mA7ah6SN78/ljkOEbbzd8oZeFLWT
db2sqFeIq6f5Z6ZdU0TzwFCVtEt/DY6JVf4XX+Mb4tKxYiEEmIQ5uu5qKCNi
vi/7eN5cujk14RpXNlFYhd/vvAcYKe5sjkLIMhMX49f176ovXjjPwWVXRp8R
KGjRuOUr4J6DTGRC6Lg6as43bPjk8eFMjlAypD+te3h85K9OUuGds61hl1JI
kvEwGjD4k9xyNwz9IMMO0fap+dZ68/ztAlfjDz99xXbhmJexfigJhuGrcmjz
i40x2lkyOZugR6L2FCHJ+8I2Z38eBT1pAmGPRfs8kV5BXd1hOl0Etu9cy7mm
3aWz7LIPUOVYFlPMe3OeQkJ64fwEIxXv6I2ylkTZktelgx88IRahWuNka1sI
ZPZFi6ZCJxALNQGivfOP/nliTys4G20yk3Of6JnJAIFweXSKXREfptf8eW8P
WWSk9GRuMA2n4lKOJWsvpp4hlIxv1GVBC+pUz6GBDKdOxBeKWaJpMF+3j5pm
iGsqvh3KV1ybEVvfGwtZs+/Ure7gU1/+xJn1bdLEh2RTZaHDI9INTaq5rmsl
eEhlvKT5ck7qGhPTrq3s4GTX6Fpdafdzxl44YD994TvizjMW1Oc3Xg72tn7C
VjUofUdjfcF+jEU91SvHWlgTznYS9xQURLUwK4IEDOgIl77DLUXVyb+/lY3v
BZqr3D1Fv9qGZwJv3a/kNJ42CM6bnOCgsVMaIT3e0MAre4bxVR+z3SIyL6oN
9uX7DgCYlx84UYVB9ea+myRCsME2dMfWKMytgQjifKvRW66CL34Ous2w6LZi
2QrbsP/u8IMQWQry9n5ckzDbCxJYpppB+5w0ukMMjyVWQo+VTrBRLwXKR12l
9CWHcgT0BQmXM1Sd5a1cAR12dGeORaw0mkmWid5ZNZ/R8WsvmTXltTPtXaNH
J8LfnyVFT/qipezK3rA9wuWd8tlJ6gRzf4SEXUsIl6RQVqtBNVUxH9L+e7v5
tM+JQLiw34WgoRtF4ItW6irST4SSNStfh5UuWskP0197VzrwHch7A4q9EPMx
dvywxykNw+xErTVxaHYgO+4adiQsCoURlbwU7ISBpEW6S9moXkbeq34G/ALV
6tmbu91DHoZcR53WatwYAt8SeeUhkXdXS87sYXzg1tM1rmuMmUudPkAqASG5
YE95bFkvQqrBL1KbrM7RIZ6zN3WKaVVsef4Rrs8xLizINoBvNVTFOSLie0pq
VogH4AOb20qxwD4iYcFaGTl+ppyrbd/C7CQ8CUJXs+8kwZHc5iXszpwdeejA
FlI5hJVhbBc0J7+fG6v5CKDU64I6WNwzc0k+5gvVyoAghNVFY2jppp/m/by5
UaqiwMw64zyj+XBgeercubWvy5Mi2qujbrTX4aPHBgHVfoELd34MkzJ5/l0f
tt2QS0+MMXJJ2fA7VzZZMSLBZZdMYm3MA7VXMG0ODG3V0M08yWDvuO4k9LfZ
kCUP7/I/Vv41FeqF8ZPu2YpFPt2P+mPkzIsMCxsRMDpqsylzk0eZfPuQL/gu
i+YqjbCXRz6PiU3pVhJVPWS42cUM0VBhJmI5h3YrrnQLLv9RPzZ4ZEeNOG4/
pkEbjDA+Ob6VUwkE2bDD8/gcErDyRiC9+g/DPPCQbj8RSthopEtgHpT1mj0t
vSG2deYfPIBQqvzlywN/Amtm7Z5f9phOYN1XagyOpj+zc3o0YDqu2HiC3FyP
5s6vmZQ9xA30Ukh92mjsKH+Vd1EbxvsapEga8EzjPdgqQJ8+aDLE1Cmrntau
4qA0fPnLnn+zLPYYBx2rSlANgbMzKnP+WqlK1P1OyM8iFs1qDLTrSIm3ny3L
Bium2G8gbiq603X3pOfa+9dM7LSv4pOzYdu6qsbLmppynk0Cc0B/sG0cBrWd
baE4uXCsjxKPILu8zqflkAos6NPEkpmSxLp6+xJ0YIaPzKi8hihLmPV3zzWu
mmcSjLwaqp5bC251bkTkYhr3YuDknwAR6+lC3aBXzf3poS460eGhoeDO6fgc
H7geN4jbNXIH/RhVMXRJWu8SPr9DTTpbrDyABcNDosL+VGmBVo3GEKgFUwE4
zhB6Bf4j0oy80HKaKTThwvVgWZpp+sB3DJ9pwfqb48t9wDf/uB10AR5rjOLg
otUck2yh5jDsVWvTB+vBYEhg5n+XmIKy2fsjAxTY8RK4kJeFlDCTdO4c/7U6
PRr9mm27tTRwxASkLhSeazKM37vNtNjg/aaAENeOB7jFAQK64+l+uJWkqQaK
8F//G/O+3/D8+2nrx/OxMB2KRmCiRFU3PcM/xcCDcHyN8oPZc+iBLn9N+xxF
jbyz+YBtWJ9WmBunosbSBL2vTqHt/P5Vqgh/38S1CVspfQvpfePWC6XVrY0m
rjyLWLWBqnCjVDCTSgL+CcJHUl4JPuoyoaHHPJrfYNSFpFA0rNpxIkTiaZyK
YM0EM3wndbOS7b46eR+f4fZ26e8ppnov7XEDRITRbpSmeoG6HEJBqKLIVa+c
lkfXkNTeRCqvRy7qAjGqJ664RF4I95GMC6RHophGrst9sIOj32We24096pGM
WH/kFG860ALJJVnoJFyFMsXLsOi15IE7wNB2OOWOoX0vgCN5FH0Cec0nO+84
mXo6AVdJb+msWngJWR419YBa4pRRcRoLqwpbot9ufZPNJGJ5Al+nPp5U52zC
EGPfBucig+9gGxC7El2mSuJ8HFzeMZtNeYPn0wPiI87H5scQFHQv/Rb6FzD/
/0PPy3/4X4r1yDJUGD65v1uo3q0V32XexVvZ7N2Y+0ggF1tB0xOB76wJPTZt
6obmysZH2++cXq1cMIf9M0ECATIy9jQwO0gTHZakk2eKyopCTNHGVq0xo/l/
RQm65uRpytN7xKcoruWQ94Qr5Pd10R9gW/lheuTyX1H2k85jrHF/pPSXpxda
nMPocwpqpFGMO+FaaxkkaWOMyKxdM+BoF1WPn1RTCpQ2tGieGm3Rz3PnfVT2
NqsR5oZgSyHjHVPqQv9ua06TQJn+BpPMLA6G7iVPj8Rvv3jGMnlpnOlCltsL
FKWF0hC2E5V8gs3LF3U8eaGQOaUEfwbpvy37p8k0dQAILM7XjcHByyg8EEyK
7Y2LCRbDtRxJU1fAemI+wMCE6jtOaMxwdfNiy/sfuqFGR3oSi8QhtOYLNDjP
xIrS45Ri+4ilkyHw4aOJAZiLxNhNojnOmpzqV2TINIfcEZ6UQJGwO5Ub93ZO
ADRHhCR06BFjFBWW1Gw79H6s6dhhq3sY3WcpMuT4QKxNTKF5GDeCtcFDQ5Jl
fzGIbPpaSWDd6R8OGpnfsMtp5muzApZ5TbWXY65p97KXCNOXjkE1WC1s3Y4W
1bqYXi6p3HAQOVSUqhgvCXYfD7WYbikho5/lXX7Hi6S0foypks5pCmlnG4pi
tfpfJo+eHYjX0yWngHn8VJCENoOlnYHzmk3KUVeK8f0aKapYvNfBLYlOyCjf
R730272EOnhnv7gf3FVDPQUrHVoRjTuOjPxJdaCfY8brkKJuzVXof2FkhDVo
O0KB31diVj/coCfZqT/TKhJ80YG0B7fIN4MEIJRqx2o9drOfId9rgkjuQzK0
4JWQK9ceZ2UnvBXOX1ZrahGDnEvXTcm6Mt2VKhScowiV+y7Q7fOKa3mnM37e
HnZtEEkq/qZvl729CwtI+Gz0FaIIMDzUugwNgtVfYvoqer6tcWTsExO2Edw5
xe/E+amNpDNOQpJ+e0iUH1COhfWhPojSG28LUjvex3bDiWbrTdJl1m8NQOBV
I7wUgri2u4gtOrU0CQEoeFYIHret3Od+C27HOdGiXMluj6+eVHHEiBI4tPAv
l3h9Gc18Rs92BOrmDHe0YgG9TB5L+l4joLb8IMPM75K3AJGrWmIT2tFGjaAG
qSGMuWUJ6oWK3P8tj/T4eStmsbhRJIv6IZzBsTFiYqyiXm6QFPMyQOVlWR24
8bhAEB0jDZpMBK7dTo1DhZKfp/WEAGue2tSu2S+BOkeuFiZeTPYsA8ahoAXp
f/ntwGXrhBelOM1s2A+tHReFhEIkEM2nb5sC3PfmfQLrCymQEwiiajteLe8J
7ZFhMyZlMs3ro05W1o9AEl3rUX2XTNJfjAlftlZwWxI1r47GIw+OW/ZkYIzu
1vgvvY3I04F5H3YbEatxdxVrAxVxRB1t56X6pvsQJAZTZJ/3jHOKZGUJFXTm
pqhK0yAwn3ySG1m9bUGqRCrOgpMlKiTsxz0LkJAr61g9TeZDX0TTLvjIzG4R
m0Bk+c9/kPr/Ypo1Xc3me/T2ynWUtIVyyaNgrdBNRz8IM4YcY5auDR2y2U3e
i/4NYIJi4t4v2z/iUJMa0qRAtqHTW6kz2TN3w6TQV6T1boOVbElmQO7ytqi+
bakT+08roPvt5Nt/2aPUhW/ovBy87dS+FJlYi5Djy1G9dXaIFzAZzJ8YdfRH
W+oHh/zeQZGZyrKOgl0t8TflZhjQZ+sE/k7E+mFmrW/ttk7NUkh7NJNmW4HV
Pr4G1QT48T1RE2xVrDPT2s0HiPxpEXCG0/7yX7bNlTKcfxPFYqDL0rfy0pNX
L2xXaQbKik2+/B6F2Pctiz3sanDRDSusw1ctvHaOpz/qm+DwRwE/fU+xbaXA
Rx16BEBUO2Rm2q46tAoAnkg0BYHmMllU/lEqh9sk9uL7b/F52otkDAJaoZFc
aT7aESRV8KFTwEZj1FOvjNBlliRvFmR4CnJI/J032QGIKqydgFrCj2Iyqu55
J03h1fGfe0y9al3KUtVlo70pN8tVHbk3nOvHolHLBO2ThFRSD40bPoljvbHd
/uBhzyDmFy9yXcNrcDijnio3KrKRbgAsQNVnonFXkjUTnMlkqQEVNBu7fGri
9Q9edFuGf2N7b6crJpzLWAoALZt+tGM0CDuh6iG6yBDsjcrVV/TWBS55qEYg
efmJKRL2xtEQ21UJa/uzakfzcVpnkvDPJ0/XG2xABLD9QYNQ6fkLvksLgIt2
sPoIeP0cSZZmqhcRJ72BF8MRNdu5fy2ZQhE3jxsoQmdg0Q8y+fnkRR0DwhZ0
RZ1Fu34lQ2zRMld9W57KtersX1X/4/pTOkFzV56k6ZELnNHugWXR580Pr+qr
atAbD/tctOy6Ca6VgJmGfUCxopsZC3PZJJNTkuOq3IBp+5NwDNT2SNHgzreV
svRHlRs5/elol9qPpsbSEKa13cnY3QdMidZ9nCcplIyiiu9V5cmLstJlPBzX
US+ivga2wpJPBSM3E2XPiDimqQVgT8CV9H3qguIdWaiuFlwFFxLIBk4W3Y/x
ZlHwhBWnJ63jOPXHoNVSYIp07gRJVCbUz/h0AcpbIN/Sj9NjH9RQmP5ilf8z
8lXAzhw5eB3wJVq18ur1ee74aAgn8K0YvmOu2dPTPhJSHRd9qPTdyP0OA3x5
U3BgG71QiBU2CD5AM/E45c1ROLqlQ6Z2Dv+7cLPNOt012nXqr/sjjTDATMxS
9ZSFfoQewoE17ogT4ihvLMY1dGFcXRCm/L2IgjNkutKlsg3lp4SAYESWT0Mx
m9MQ8550PPBNcB/HF5sX2E9uKn2G4OLWWzqoBDES+3MjQiOBCIUEbUMwHs6d
wZcYarr7I8qWIbexQ/LSF/tl+O7sm4iuslVTgef/NFj/xEbiUgdNOFLfnuEA
GK3iIQc5hpxYXcxRJIGvAxvwg+ep80kKfy9INEbqR7LohtyWNbasbvl+z8ES
PdsXvt54GHEAurtCJHLkKbE+KXCeh9dvMQWc/PUEQ41HHgz2WC1FKB259Os1
T7xEnq7oj3D5ejvHxd/zrY5cDJ90RMy60SWHPQ8CsKMZ9mYj4HeI1zPt/y4u
XSiE9JNx+bYwa5+DYwMr4bF3HBgs5aiEUBAH67EdsdA4DLFpIezuUB6307mY
1dvPQSSMef/e5NABrzbtwy0sfGtkhL4DshidQonSrgxlYA26b40WOK63HdYv
VUJ98Q4XYsgcEBDANLDE45A1sVOAl/AwaBRa1I8HdwPookgl1sRFGudkw0Dr
DVRNbzII0lMW8ZJx7RqvY5Uk2u607On5bf0YCLNQvkPiNa90b4zrU5OXdY4k
SCcFrfp89YIgoIYQCOA9Zl1Hy71uMWa/bgSDTmHPQiief1QxS/0LkQOCRJE9
gubXwwthtMAgdiSoMFakVmeOVFuqveqMULESjDYeeOTWJyiRK5moUHYosKrG
WDQ8e7O0VB+CQgYSMdiZJ4E3X2cSklvkBiMoM4aUtKy0FtUAZ+vg17ktp1oN
IYIHbwsHGDqz6/s4urZJ+XOwPBaIeV24e87AzLA94mbUi/Lgj0A40JSuWowx
a5RXPLBvG4xsqhqYiE5MWLIBNYte57rSzsUHYHHTSOrLX+4iJ7aX6hm9T0XW
xvJGWI/BmljSDx47ylb33pNzDEHGDmwxVP+/ZiFaUkDGvfmlIv9F8Iqp3qWo
sxcz+1w3NFMTN6V3ERQy/iU8psn/c993qF4Xny+QErw0AsQfnx5lJXjPJOOh
5oYNDrHNmLndyeTJL5BnK+2JLgEifCfA4MiEQHv0imuMnZGhOW+d2Nzs0F0w
agEPc4ZmFj62evNTd3hXJlU30Ga1iNSLFpZULIusq6rVyAviG44b3Hft5UNd
BXocI/sqLl/7BizT7vv/1m3fCA91y9XdA9R4I2J3kBtLgbNFK+BV4HRCPion
zzB3Nd4Htbqci8xuBzL3hpGSrHQ3U1u1Ix6K/ZP9Wk81yd3ly7wSFuSSIv45
YeoG8IUXJQJKKR/An1X9WTbHktMoXuQ4mN+5MsWyO0lzbPqo0Fak3qGVKoVu
wqf3qNw6bbF+Opn+UCuX9YmGg/faIc3jikfs8ar/UEVgmavYSpd3k/7JxmHV
5GGCcOpyimjd16tpIZ5vro6Oio5EPsWs2oUQGf1ApXrGlDXopRn1bwtYaK/e
Yt6jfLYbbB8WVzum1wcA6UWovq7cpmpkeK8Y8qy3H603JIs1zbshNXhaOwwr
EI0AuLk3j6Kc3h6AIZl70VnEXxZbcFrOJXNbG9yPgXTRkAc50OfLMaGD6dMA
4iCpOB3aD/BhRs+3LIQk5IiRDersDD3Nu0nK91ubyUxzUe0hN2AYqJenglZY
V8ObDrDACWSbxQNyooucNVXetwa/LsblrFsc0AEgLLFvfO94vkqIZFcAVJB3
MlaUlzPy5mFV2iEmnU17VjXW/p7bVyOgUxvLSg5pKLTeex8lGreNVgMpGVTx
Qdl46sDZdYLZ5nt630fYlbFJwyv3/mZqxPzf9UBUs8Mdtj2cwKwNZtx//xj0
ZfrlfXObxG7cGvEPmGmAKIHzDiW1KLezVGyEm4eDO1nttjF53PoYnLOe7MXO
z7wQRQm+At5kdfVvzophitQNaVhG5llsbbvslKCf7GJ1/7/UyrCWb8qycVTC
v4vk543OT2OlSrLviHMUSKOGXayYZUj41ExkNvLYNtWzquA2uA/a3gQD0htW
xaCfOwj956esyi7z5R5JngNyU2SMQPKDgSheQK4nANDlhUIMQCLG28n9Ldu9
Q2Z7huULSIkF/+w/nWBihkmYeGddCgzDPbeKWcSWpRtdDt7e+ruIMW/ZKJJ3
5wG4yzuV6SmmU8nQyQ9VJEIQps/k65euHDqXMR1hUpYa5nLTQKzuCGxOqSYp
2TXUscvnEo9/CiFdqRpK/cnRymGWJtSxNOyg3nIq2R8I0UDOah4437l+gdq+
aVOAacn+WXI3bq44DifXhNr4snK26OBua2vFjaYgWvWw1UdyX/BEgYvmdn+b
HToLDOQJb8rAFOKf9YrnPiS6moRYBYS/81v3MpvIWC5f6W3XUYDZH4IRbiDv
RPh+liRWcrpRdORCwTMMjiYxjun2X38kSWGqvKIl0KXW3cY3UDIinZTVigCc
HPzx3ENoz0awQaN9/v6iaGXIY2WSpO2bt00j5vOe0nXVCYyvkFmS9/DwsHHl
uUadVZxrIHBozf/oiwTPDbMhHkPoLYoAb7XMn1UH6cEsnGrWnDfuaoZUZ4XQ
0pyYHvQiGJzuhuiqQ8SfHjCOnSNV9TCowtTgpPrG+g/lyC/RvkIToAZ9zQOr
z9a3nypNPJrmiqXQ2sAZDX1UFgnJTXruEgDUpopo/bZOJG6KqlcB1ZMD/SeU
2l4LZTE5+pZfEygrzdlbfQvxfroIMdvRf9NyPkiGoy5eIJ/P0ZrZ1yMGySJp
ccsds372Dzb6rvRScBs98EBy24mklgnl12iErO1lvtkpGt4NXOC5rYCNDavn
MZjAa5G0i/J2awUTpvle54QDelovrACAKq3Qu0581/x2v+pytIeWVsHVjJ2O
gnZ/f5akOWWoh9inbUiW/ReNdx4kqpRfSxr3U8Awg8ld9CmVlDXJf8r/G8XJ
AvGwu2fyJvAzq7boLrr1FacEbutsvolnr0qrMTR8CdHGKm6NUMT7ynCEQJYS
M4DaqwT+atnobBOOJNjAsN/pdB+DI6JJ4K9Bor8RFaS83eY1jaGpHTRw77st
Zw5iUJ87YYwchqs/4tmemStU0wSr2QIEOdyLxFlxIf7jsfBANNgS/kuVp1md
R+Tb8aS/u48avZcEYZ2fGAI3A7ynylFsWe/5Q43vCcvrcNBU7qcwWqnTTWDA
o3GMmQ3ujddRAg5JUJPMIhcCF+Q0amNIX6poDT48W4UBLminq42q9cvG1wyu
/dB/7NGwmu9mz2Fl2oo4dc7iPo4kc9PQ/j8BeqrC9kst0gaEN8u9EQ1avytv
run9DH4pkm2r3n6UUFpxtcH7PC7aGu5ATBeWo+rXW65PI3CdShqr3xKEuSG6
FojdeQmV0wj/yz8mR/eG1If7feqIoQOUVBJO1HE9fu62SVkVnZ6iy3hokzEv
+So0AZIt2O4sVg2akSQbO2Kxm8+OzSYDzznx9fRtx7p7wrorlvuO6F1IHGjX
M7sVpuygIgEeFtSOkJJuSvBZz23GP7KUu+t4EYVPK/XmhMnuyxSfjOVfZ7IG
jythzd5WkbpYxTHltfm2xuh32TA009PL9Dr1//Zn3ocrMRKoDI7/D7hl8tON
KFTG/6+JQcWDwQdjuZElB0h6uffE2Aa4pV51dudLbQUM/EXU6CD05oGDroEf
WWXB8rQz5vfvsk7JjyXlB74WorzBFMS4e+qLSN54Fl10vWD/Q26+rTewNvDV
xbyN44/d8lAbf7QLM/4Ntn173UWuKtK2oZF8fDneD2//QelVsNPpZ57J2k6I
4yyYYiuiqSn2mXL+Rz94Vl1Ouk3LCYa79lyntMyGLmCDf2G2bm5n6YbkJ4Fn
cwTUz/uJGCC+yjlD/KRluUP89PMhevaTBkSg3RkqdHXKN2qGM1XRe5MegW6U
BNmCTbM59+j4Fc7Qndd89YHye3UNLRFuBFXXEDejRSzmRHd/j/q2Zkei2fNb
y27y/t4cSTuOAUYs/g4MMJnygzDwFAkERqbeTWEepDLqLQK+YNJhRTdjq0cy
yRVWMQrRN05J+4yNvaZ08MKO7SYjpiHqRM/jlec6/xwIvvOZIIumpCMxM9jc
jhNpZRDLVSRB8OpnWGX9TEE5BHHj1F/hIUQumgU9FArhHs8BflDHZbXW7sAx
ytNPCBAIFg7+N/ROQhpX5EZN8E3hoJV9nYwwaOrIB8rv3WkpmTnAMRzjZlRj
VoBtv+0OXwmxv3YX071frXWCJTGZSNywdct1JxD6QQ0ZKhu1C7iVrH9fX1IB
rA8+Gf3hOh5xWZPlJjketSWa3djAvqRRuKeRd06fAkfT/v2H6iK7drgG4sDL
kqfyQgbJicqCB8SFJG3O8UBbwA6HKjNu4SqVSdLFcqcrCai6vQCJe58E53D+
TXx2VS0nlFnjNL7ecTqRWxKq9gxUHZK1vlSc99zLjeZd6polC12TUPjl46xc
lC5CoomD6AX+EZfX+mac4Mv/JjShnVl3YyyVEqGGm8IpJVDwKy3LU1rTrOa+
zRQHdf+cTl6L/xzPLepYHgmLwPlm0PNZqzO7GjyqoQmNXIGBFGRMjun6UjVM
Bvocp1g35hW0lLkilXA/Si5hqMwUNGzVtWStSL/0LXJYvkddg/OHBvMemmGt
XTf3wnt0jtdI3wTtOTOH7q+LVdoJX0cXHX/UlCNGbR0eUP5mGnErZEI9nTQw
BkuCWK6Tkz6ionwV5UZfBt2gpYxpkhAAZA8YZfqG1Db8Yp3kd+X55LWWvjSh
3BgEl47074Y1T4QSOi9bV/yntaRlxxnk6gCWuEtlHlsCYFO3Ga621IGALYY6
KbGX5PBP7NCH+fX9mf0MTSxSt2vvScc9JHjVPSvh2qEMElAUeuEyAKb52l2+
/YovY5E5/FpoiMZ/Px/mSnULqWaKgY0gcpk71ILVeTYCYoq8qKwfw63a4ioz
x6Wb34IUtKp2YvL7nBa9L4bGiwTD+gcRK6CTY7y4ndD1z6z/8gdCggpuRu1C
EGvPXB1JHTqW0PNaFFWy0RX1vNc6V+jykCOjz+5g/KdmIb5rJ/RFuj2BFYtU
9e+EdZC6p5cFn4d5bnp+ml3kHGLRqJHXg9wSmRkTmnsj6FiULgHsgmw1Tnes
yW5QO8QBAzyir2QKL9euUbC9u+MtTcAEiGztkpXhCgbc2u7ZKBoxm9Torb7w
zlHvbigfunQpbrngD+8SRmkhS0TCEDYkywymanOaVwHN6Vh6NGwaadzV1JPx
wr9whzlrNb1xzKvz6RpGn44rCIUBMucBMstVQfqnAb1xO0bVjvhSigIgn92l
lc0yJg3N2B89y2UllL+PoSN3tSCU/qbEzDDluYX0jyf/2cy/XmT0vObpRFTz
Jyz3F0SFpu6KhaGYWOy+CUcTAl2wi1JllZA8KkLyARYU5JmMvYUQ8+5QLuw8
S+OwFjyNx9AYu6vXWlRxdMDXdu+2QSN+qjq2ag2qTd3mWBJ5xD40ok9xRcHZ
CTWEXh1rDdBPLq6NmC5eG4y+DNxjApNowfIch1JVT8xPyyhy4jwvqE4LfTQk
0FkVdDjHmPN/4rtTYaZMDrfddfyQjwwB2W9cGN3qPI+MWb9XqaWMrgoDDNPQ
ww1/Xa/m8wqLHK+9pxCXMg559FWI9XAEvC7JT7xdsy/D1p0URt921vCvR3jd
dWP8aeiXNUahskvt8IcihPKLNos4QnE7g9todGSv4kTTzc3OCzWybpxYi9+u
A8U4oD4u6lm/7H6nATrqnePTJ5L8Tay3TVWKKnmsdfnVf/TkLcrrZkIgBpbP
EZAxa1WyxWMwGFOP8VI6GRI+3k+U8YxknHvqdNktAbAdPsP06ks7cR9dxhlq
DNLIuLBgufTfZh52e34e7GKnlHW84Ziyk35FW/eZ4DOm5QDcrXIi1f3hd1tG
dTUyG4RGZDd6Vl0Yi0iOijQSTrg8cN7nYljpbVtwLmGDUOtXdPZvfvLKnmwf
K/UocQadqOVhEthALYXeAtoR/YYXsyrSNxQLPVMrFELxF4dS0bm7/JP7pSQw
kcMTNbdtm26G8T+PKtZRkRXLVjOZ+mRiZ+MGUDLnZeGBhUCQPs3K2hocfsnM
PAiukMMihtxWmTTv3wnDXmNx/3lb9cj72sb2cyteqz2czEVC/aS5kMHBwpgw
vVjIsA6CeUHXEZVJsuvuWBbLRhbAaoiAOlb8GuTg175AnEG/szXIoc8seuAC
1jrgF73Ur1QecIsbQzVl689Kx70Ua/Ip3FpqHRxU1GfGKsBz0DzRWmOwpZ+/
8L8GPBv42Bh8zhe6w3+R3MuQpPS6Ie/aBAaXUgTm/wmSR9INRKV3h8VxZ4ft
xf2KX9pxMLeTcdDZE/XgJrE9K6EFxOWC8fw81ZzwgqkL4CHXKruvUU+PMGm0
X1f3ut4rlCW22GcoRC3UrgJhfOF9u64AM1O2/nIwhC3rF2r4eyu9tp/n8qPU
wRG+hJt0iQSpmwRFuyK5B1D5bKJPfn9s81eOxtVxN11jje/WgwljujmAxrBN
15IulAmcAFvEv2u46id3QfLFC4mVZ6w2tAJN2nCowu5askoiBqnhQ+K4ibFH
+qYcRBmXOSQ6BbK4CHdpYr0OBeWM5Od+hOKYJsGMc7+VsWtJ6xWJGmx0CuqZ
hB5Aeq/OJXox0Fr/UI65zQco2NGM/rS0uoOW5BpnsJlw6q3UXUL8Oq0ipX92
iUbUg+2OCHl0ToV/w9nHhsARZASBogfdaYJYMqWGsiBdHoN/LQ6JAxVRT6qY
z+eDUl/lBS23faSFRIoMGwLXuqGQPKxPVE434CW6Wkd5VRT7xwGafzSMsZ38
b3MNMXstwWTbjfeZVBJWzk/NYubJzzKWAWcNyEkzAdO01JYNf5ko4P4apsGp
hJeQEl0d1NVakBPdkK5dmuq99h8UbRRQW8suQO8u1qS3ZgFwY/rXzXpXT8vQ
cw4r54ASt2+32kNgLBs2al4KalVC3mdhZ2kOu5xyAWvAgH3QVvQ4Ef3qms9t
dsmPJWheiD1bKEenpMa/fsr//lfya3oItr4rGa+SUh3uFgT+blk77ZahGIry
mTL8ucWMxfzD2nU6xhsjIRIE6Dgu9XkyxQiiKDDp5spmJaYAFqdmGCRDzgdf
gb3nVgTWGAxAUM/P1fDbQs5J3/c1ClranHsnczrpgpymPytnGtqVBakwkuMw
ieCOBnTQCGyxgJBk/ZQAW976V2ZQa1yCXjuL2JOma+MCrTB1oMDQXNNeI+as
MVAEnQhP7Os3fRfJPlvvv+xv3ly/MVUoDZ+b4ASHezGg+znYiQUdAK4pUyX2
E+jYYw/TiqT4BOEaJ+RBoXz2weK0RBK9gwyTeIUGP8ejNd4Xw4AjL5r6CQTl
LmxdtOja6TvNqLvMWI+gVMMY+FLVAa/pPOvJzpcIm2zCXG0GHQVnYilyvwtZ
+ulWUf/zc2N/u6MciMU48RkVDWO9hcP8PW2Js+c9l315j9SyB7vgt+xnH6mS
Nbqn0TIy6rrzptu9yo0eYD3e1sgQejUWeEievaTWZdUHYuMhkm97639R2qMm
ynLm6pNR33VglKcaVPx0EBfEdo+Rass+MVhKi8Y2CQrRU+uJ5Hy39I1xp6qT
xxmUfHaBfUPCjlKhwUUe+dz9yLAQc9d1QIXIqQuKLO60cCDlvLnCebJqsGa6
pfXcmxzQZnJXLrAqNfEf5KTwzotz5UMSpURiTYHePuMCWTNNOmxoOhUSlMIf
6ixM0UKIrjz+ZEGgw/ATp6/rgXjhF2QaKtq0e+hAJAbRZwzGvJgqCnOrQ+72
ab7VOTxo6fWaCsO3SOsRuokKcecNYehkp9tRw4PXNXCcYNEJRUa+la3QLbYA
7bmO/zVlnR8ZDM2/1QuZNBU4aK3YYWaigClFHBzVXPo8O1iYhX4ho/i3Jfuq
jSCWbBK2ZlXbwvK/9b4VJbfr03ldiL0vt1wahb7aw4fefwo9aB2xUu3IjxfY
SO9kp1yrsyjSFbDCGHWzl2MSikltU/EOLlpVUdW5+A37yoPyaTwHd3YOxmih
A3iZZRID6aXoZl3kl5bGGgTtH8gM8zOgpKOED5YXdPhyy7ux9AGP8ukUfmPq
W4VipVJp2eV2u783VxyWssLUrJTniyMppf5spc11p+DgUwbqqWPZ/3GEvEfj
jdD5cvWhWK0r0k8GylqyAxIRLSUgkwBkjNzMYYJhnM/jRZcIjNJkr2bLi1+b
e5Mc7ucgl7elGslri4TB0Hz4Lx8wlsSeUhaHdGfLAaeKQfKpv5Hj55UvAz+R
mnZlThUa90JjGi7toENYFpNFcb86a+HUdXpI5IUeHDTKD4pfjOm0zN6SDYnT
z5DUrhztpo7mR7MORqSFFStV4qJwWwlvzhanYC9RO/512ZCNST0Wj1uAzOVG
mrFjXegNf0/cDlKDRRrISpC7dVL0h3cZ/BOZU5CDqsg42CUemXWdO3XLZ3zs
zHN1p5QSARn80ytPOgfQOa554EI/xI9/wWxZpAeO3vjGwdFPA0y5HcZ6vN4C
1SVMzfQihltna1/TdrhUgyLPMCneE6fPoc5PSmIKg6D3KAzHoW02nqFDULD3
xmG71Z7kS/n1+x0nXiElvobVh/zmnKN45O4Q0ws3OMhjWn4A8U9eYPf+P1LY
zzx+WbP2qgH3kIEuPnFDFQs7wl3xIvkTjjisjn9Yg47o06VWP9FAhXHxI4sM
NitG95wwNgL7vFKBQUK/aXzxWubjlS637QB/bA7oHmAb1+mRAJCjgsaCfAOZ
RxRUxwS8BKnCuCpw9GPA/IWBvvmFQBhOx38JRYs+3Ac68I/N4/mCpVTYuwKZ
f9fGjqP4vxyX24akLDVuZVn+HBbXoGvsBXKefLPfhmCalRnrJhygonCg/Xmh
vFW191g7+l5oPpzXmZ99IytWVDGr2/fHAn7oMiD0pk06Oa6aiDy64B2Mp6J2
Q0CFysQfmujySvuE8oXOkBUhflp1apyYffhjw797eLXZeJ5jwJf4rQ9uiigP
o63wq3NcrRnOocwwwHspknUn69kEiZDPijyRCy4T0f3V5439TOf+Sj5c6RBV
/X8IwFD7VpuZeMLT99iNZUKY1gui3vVxDnYkM6/B3ENDAYC5pdRFKIuCs1lB
TzmeLqLrICbx17EkPyUh5wsvFjujwpqrQk75MQEG8vwaSJG0WABpUUEq2WJr
7CLEYi49/ViaOepzh9xs4eMdRy1872luFiXAW4lGiafBglc106jOtyBgqZdp
tcd4JSD3TxHLH+CsbjLs4jpmD91yhl+5WQDvJf9cPS6oru/IQgANfe/Oxpx5
I/CW8wLlxxk13NZZQ/oZzpQ6ykomJD2iumL1ZhzuzSzVUWc0XZ8sjBA+obBC
wFlyK8OsvmTqztwwF1uZ8EclutpS2F0KxazAE+E+R1UzxIPM9HER1OPmxJM8
UFKGFNHYZXF7OH+fGsms6lUnoMX20+WoPbvAh0PfBs9XWxjw1fyzhxOrqnSm
itVZHdjpleJ+/iIdqdQktkcwMzVCh7FLYTjQt8ZYG1TES0uWsMUXFdHW7EWP
jxDjrfQKeJPdzs4motLaabVYtvrSCCcisICgZvGtBuIXZkJnB75bCw5KW442
aOHRct0y8udk79DY6xi7Brm9KyBrXGKGLo6QLQqEzFiao2hO+DSjAHhH073Z
0Rgbr/8oEbk08UmIsrD+Ck4QMGXZdiEGgWYW2fmXkNZLj57i9z+mr6xlDMxk
GdGjRAdhGevk4KOAWEn4Ip8kxvGQKt4pQn4PCXt/CFju4iNnd+cR1yNmvVEt
OzztYtCyquVcwt0zqymckPCQWda4qZGYb34j7mrNVh6aGnHbX/QkIRWR6Xm1
5V8PTNClKHoRERsHpbaMhSQAQsN9wKCvaQd/kc0++F6Y6FbOFB2lUz9w9Aku
eZztyLayn+QGgLdiIAdlwunQ0fbxO/JNovoQzevImWG4UR6XYoEfwaaDpddU
97fHLFYcghoUaIhX0+cbSoSt0ljLDpc6abXyUZ93UZcIr/YBFzBHzyUUkHgZ
zlmPeVzlglTo+5x04y2XVMoH2KVc5ZL4BLWpfEQuc1yFaAUTm2jWRLd93VUq
EO0ZDgvb6H1wqWL2+pyufHXJKO0N2H7SOD1Qfx7CMLP0xwH3jwnPlu8gHXX6
a7mVKGG6SDwE6f7uSnVXxcATHy+5A/aqMiWxM2WC50VnOfa/zofqqSRiBxUs
9UhcWZCyP5sC5ck/yGGnfyOxXUqOAv/+Wau9t05IyiP1Ho5/U7uf0fWNp6L+
D9TTN1c5UsewJ6dcwSv5e0X7HCoO9mPqCT/6IPqn+thURyU3m19BEm4m5JKy
BEHNE5N+MNDo6Y6Itylvtd+kN5A8gtETwZAIpRnqlN0LGikgnd1LiQyvkS5R
l1XWRQshgQUY3lYmgEudnZ4TdIraotijyV6RwItnrAYdKl4/wJZopFiPh5Lc
A6Psr5jcg8aG5YnvqGeLpwXaT4D11ycl9o9/imKXqIqWZCw1o3yp3QDr6q17
3EUonnfvqJn0wckmdchc3LHHVOFIsGp3Mg7Am/bsuhZpM1K5IiTr9nHoVLqn
uHhSaitH8ZVSeWQX5XXLKyccc8AnOyYDis8GR2SlWDIIT4wnNrMS7TLu8Z+/
3ac4TamnigjAiLZZklqyQAhYWhrq+3o1lj7eSyVNG28dQV07qjXc9LN779dH
mcf3XARe1rESeLLgLSZ3UAX7TqHd1yoX70R2xo8nyat7j5xQFVbNLn2QTsl9
MCPSu4rkQVg74mhbZfOda165Dx1wsa1sA71HiHMliuukNrNkePk/R6FJRMGM
gLkIckgGzDjo3Zfh4XCzNbhqo2S7mqlUDIMu9YSoJGKcDuJ+p8dfPNZOrIKj
6Kuzsi1F6XQRlIBCNIJ4UO8rV6TzOpg3Mo0nkUYOSIWQlEldvL5/TUDjrriH
dgV2x6CFD6XXxM8Mt68LstoA4D0P5wulQuiNunywgwLFPH2UsKswopAD4Xsu
meHdE6ZvEyAsGrILTZ1rhoZ+jqgXLwlhpLIbr/t2UTBJOcRqDAXUa/SJ0bSb
kup78M14d/pmUmtzTpttpr1c+p5pfchwHxS++2dykJO4NIQAPME6Augee4Lr
SZLw32VAbLBxYJnivtuAkr+beVTp2svCUayjS6gtdNAuzOfTfDpQpK0jtVb4
RhWpVr39yny3eSsvIvVti+N4ucmYPKHoYv6IlaB9XM0bRIpn5A//K9xjw74e
22LBTgDVWe7v8vmNqu/WmweECkR4a4/CmXkvKDnFDTeJ4OucbxWDoxr9jNtk
+UqhEDofrU/ZX/mK9zLxlyw9NI+83HWaJwjknRwxH5LgSdPZnO6ImlWhIYSb
Jt7igZkJAVAMYKH+Tvhhabmqzd37b3wqeR6Wyira3fjMBnvre5WRhfSGq1xL
sYsQaMo+Usox/UZ/gtueQFCef70BXIs3OXPpIKKg4Af2vi7mW9Ol7OsZygRP
uLqaAcHeJL6GPDqzh0sFYABsDeqFI1RlVFgc5zDgMLejJjkyQ5vtPd3y+zWr
j3ZS67kWGu4nXOfTRn0jN41zKsq5Ht3gqD5ViTMK89eSIZ1GOTM/egyUpgL8
wILwjnG9sSigkNA7p0armV0PFqrvz5vB2tyScfXgWv6CarhKXfOSpkvLj24W
B53noxgGuDpABsHJzSbRGmN0eGp4jgLFGc/qV9+/PDUGy2qYMx5CBM7pmsQY
DfhJBEO5XWPskUKjPkZ3yXW9o3fNHpVa35/raH7CYt2SUk67npGJMOY+9oci
32tWMNeIDyQBB0lI1d4XJKyZQTOmxxNlAJMgFP9SigeXO0k/H+l80Qa5fpPI
jtM7/ot6/2tFqxGUsTvFWZUXsUEY8v7t86GApRL6gGB6MjJhMMeo+51+598m
sIqxkx5wJFOOjxYb0o7hnTuWm9bVLFjQmItQlupIvl15NEzTk8upop0Qn9s/
vr7pRMCKNZCksZ6LzfWTKXXAvJ8O3oREJr2zu9/gpDanIzz36emQULpQQCBM
cx8sjxFZDZt5bQf6IvE4RyMq+y+Dz7UiEmHPZ3ihjwKHcx6+lNDcr+9ar/iB
LCcUfaHh6nI5nhcsps9EEB2fLIZBi9RuN67eCDEMC7s0M9sQleV6Ipzln9ux
N9k9QmzZJ5LUSVDT0bHuWkgxmziklAWd5xu2pLQSEAJ01xNIXX0hA1FM74Xd
DPcSMzRDb8pdpTmsHO6MW1+mctn4/l3MfNgR5shqei9SaGXUKDMpyv5I6OIC
2F0UCXXlnJuv6tudc/gOjr8aVJZBo/Oun/B1ivmZs4fqeRl3CVLOsuAJik7D
fJFwsFreVzo9CoPch7nJqHgHveC7PzlA/j4h39vTSGN7QsGt7jtEnQVmUJky
hhCieob+ZuX2pcsiJPWw0CXeQxz/FnUcVx2SD9ZS88LdiSKt8sjV1YblxN5R
dmh04YOj6OwaHSGJK9Ey6bqUXhxcnPanCJut7XGYrgzafBpnXlkRKyBOTYtg
DFrkxNp6MlNR1XJ4f2L0exu9FiAcGe7kSrOW2f2luS46OWjnWcc0HIcDU+nI
fWVL/oelylURrbkOocyvI0I/XJNQt5uv159Xm2yfKfDOYnox2bDrPeF6Ci20
Vcip1FJHo1ugfmQvWOMM3lIM1nVHR8AEGFNNNB/ryOuAG4pNieLiZn/qI4lN
mY96g4jx6PbkrHW6K2HLgb/x2jJeRfWSuXsQBSvm6kllbLnh+7AHEQ4/UOsl
GR8jJ0xCpyaJbrWK7+8sY4Brl60HCNscIQB5JdGSbncLEMAnhev9nCfEKqPY
gZV1EylxHWVGi5uQ4b9BC+B8gcYqe6yCiu4OL0zjvnQqfdRTk/iBESbjnNRo
9JjA2/jAkGYVstxzTpbakJPeHEkfi+Am0O8qtFXimQGWdOuczyS0/NTBK6w6
pdtyh5yagfO7UAcWr0YtROgJI6HNSpAFskDSKq28/zRDg+oOOfqAd6wAo2ma
2B4rrI65y+o8GwU1mcfm6vPdmne/SleChbihklGygzVev+t4ss36aTO0IYUu
EnAU+hLUP5BTU6SurtEC2XPhP7y8Rh39QhJeJsR9MRmOSC3qUoL07LUhgYKI
jH+ges5TcQMBKMJwr8drfRyE0zwVuoDYMCdmP7cAmnNlKYKKpnVjRnt6BDK3
h3Fivny2oq82jwcPCqG2lYsF4i63ZOarnixz41osyPBcg8ZhGAxXBoUdAC46
rpi5JqXHxLDxv1SAbXP43dPKKKMxlXHsCWnAajxIEiqv9gaHx8tctX/Ry5f/
/maSz5lOw+mPbZ+2CGdmefUvXOtcRbsuA3Md/OZTDSXwR+cDlzezoo05+Ohn
jtoigZKdOQ8W9N9QSWNkk+SVqIpojQB/GVdWsEGsgGOXFnuHgB0d3IpsF0RP
wzlPRpxMonCylh0jqH1Y3FpDHbdBMVuHBnXyIN38+iwMVtBPX9zlkub2zaNO
yxETDZIieX47o11NSq5hUeK154ezdDV1XLLK1KdXz4PM2FTS7MKgDpiDjKV8
qJm/AZ2HlWwQln+dDr87uM+k44vFkhYdK6x9SKkuGdyoMLaX/BjUc2B2TG6d
DisLu7tmfKJmMoobsuh7gN0UYvsRouu12HMd86y+RQaPNkJ8sV9FunyeA805
dgU3ZS33NW0vRwXdn0/8Mal4lx+r695/Rw+pP6Y/uYFVi2zStybCUNaaNKpX
ezTlKvzkDzqUoXSNKHHnkS/818w3whS6sIbbXZtM74QMvxHDikilz/m/SaUr
bcR8diUFogZzSfmxw0b/2/FoqPCg6rKFlFP5O7yYiEQB3nOBGsosHFxRuvdN
ao+fifFVCu7IyGWICTgv/Rf072W8s+EfRS7i7h+ac4ZbSQ9itbLYXvdfI3qZ
2XYQuMKwudBMWbaw93/BvA8KkQxch/k/3AyQx3/X/mGesCFylvmh+gDeVbUe
XH0wXgYm1gOqMmI6/J1vm4WtxgC5GJSH8DqspXVgUB85dvANMVSSzj9/U03e
euXkIHHhMJWg1AEEI9Pm+leFioRghZsnArA4DbtofEC2K+AjfPSlJVAc6s/v
W01i/Y5Xa8LvLKyQjToWZ4Ei283u2Y+QGxqv1RoLf6aX8LHOw+06ETCQ5Lyr
m1znwmURLrF8PbO/mIyPdekLlPXR8OwFhpuVu0g8EJnBCJuWbnTbdq4L4JP3
pGw2UciJVAyeniiJqOCcVoSJaK8yQURI6op4WPePRJiNpRB1352OWGx6r01Q
nn750+VLzBhfxZagTYxKh4vjxc3DTO1kRydOpg+4ZZzgs2JcZK6kXX2dXlvj
IXth3fPU6sBq3QdA2dWOcqkzGnAhPbtc9ZVrOplQ6wTSNYW4pLHgSllYtMhF
LQqMoiGDPV5LmXPZsCDXe1IZFviOuMR3oeqOeKJ3j4RwAseAPQGnnrCmPqS8
3BZdkbF2+IdKgD8buObmlXkvr5ndyi45cjQPeT6+bkIw2x5YqpfUr3LS+sWn
nI+kzzakrOZpXcvsn4FVKq4edVZfa1Q4LkHI/nQx9p7NXXU/pqswMUFmdO91
RbGE5/OYnBl6+POClgCD+PIH50L9W/jkXZ2Ka87PvBlDEqLA0YxL2Lx2fZxM
GUjOX95/lv8sex8y4ZJuUTDSQlthwWgZHnfGySpleTEDK2qNTujgfkQxYN9r
fOdUX4j7IVth2AbP2/8pk4gwB3CQLNQJgH+45QwlZ9YLVw3SvzLP9Gf8VaLT
ajJkA2PIaZK0FEki6uHw4q84VMl78lXLmjEs5DF9Uz/Z28ukB+es37Iyix4u
TPkLOJu2AuC6wIIi9YTXWBUkJZBrosrw/4LbnB3nBRQtGwh2NffovX8MDViY
y8kvhvu2BBKSNdstg2V3GqBZ2WBVW/nmSKhNpQVpSdeWxB6ZCeCVwd2NBGf5
URidVMxZgvhDnByreXhiFhTxc5bjdZCuRrPF8X1gQEE44uuYRzzDkNR/NDHg
bvkwCQPGZHRGziZrakpLU/B78OaeGMh3UaB82uXFJMr1xl7RJw0fNoSOI2cC
nanmdOI9d8pxmNCRq2NJasAE9sK0N0R0wZnaNyFMpuNAo7sTuytzVn7/Zobv
MYAoCwDoZOVakbJdl1V0gDl0coQ3bPlpFZLfE9ipCy5d+fmxcJbvXG7X90xZ
o74GPiOwfr5ATpzDCw5qle/hiNpPZDeSNeECxfAc5ZaWUcQT3mOceIVPBmwX
plWz63pKNQ/9SQdiX3AA8FVTw19N7C2POFKpGrM/3kCmlcRUgpuWFsLqcEqc
U73CnHX7TMtjBO1LPRcFzF4FpplCFRos7BRGHJhitl/wdObBijuVuVsHdahJ
Hub+CrSPhuc9sbHACZmkfzjbKbaZ3wXY2zkwtuMwlfQHrW8g5dcyc4V3DaEQ
EALQ/cap2mJK/YJHGSa7WGPVoRFpLG+P8qLUEaIcPKiQS9jXTF0c6JuB80g7
etH/VORFwv8ZvEmpr0aGbNlA6Rez94bIdGCx78R+iqh9nWEdZYW0bh+C2sjQ
YNMtpzdG/4QbGdsDvlYsN0UyH8RB5wlN2JCsJP7WOmu9tyJnk2Ix/uYMVwbk
xZnRSQIXkMW28DwYvq0no0uw4TozgNJdkdDlUO/eGvSu7+RxwRbKdnNd5KMX
VJ6Fv+1+0XiJ53hydb4cCsDZX5bQkTKflKGPHqdDxABo22y4IekNm8DbvH58
z7cbBwHln2ctWXWZPzKy+pcRWux7s/lT5Z6GILbmUxaclOgBM+81NCELfyI9
9N4rgr3IGRPqubcCjJzjbMQqoaCIDvgAkKFv02Pf64xmBK4JyDMbunPRSkh5
AvIaOo1PRjYPno1NXumUz3MmLhspp752T4TgEnA/qZRqsKNfK1CtOD/5S4ge
DOancF7ytG6z6p+zoMzsuz1oR40rtcZiZT9HhhFZ3ztYGKqQiSbN8myY2/5R
5kBROVyFkd8KDq20BSpmg7Nj2wMjpgp/E2bV35jTN5mloElztugGTYnAJNn7
ozixkWzH8EDXfrDxNGW+FW7o9kPWCFhu16Rj5vNX4xxRjfmJF1LRSUsLY1Mf
/OIV1SfmSDSvPx5oduk1L/KRofRJzCnb1PWxOnQua7M0z1Ma3rvl6XiEKeUM
AR9jEtQjmwcM8hjRQ9nAt55ix5koVcahsEiVKxnxYmXtfuGCwAobwzoiycUp
DhpBseWV6jDCLRFi1NUK426TomwbdO0Xy15zmUiysQ8/LFz7oHBcTxyJJpyb
kb6TGhE9yzwImAvraTaubF690UFMBNesR6tPUgEibU1oQnQEg9OR9vfoDqKx
t1EaX9P4gnNMs3DQhyHnOsv2qTTtkBFC0vt6tPJGO4lcGknRHqaX05JeZTp/
5KCcjbXDZo5Zp3QnBZD1qkqIXhJnqVp0ph38bgisfH08szTCO/pHpmDaoFDP
ZxnxiNAsuo756La1CZq3TNi71k44G2y3IkErQa+j0fAJvh6em8qOMBO5EtEQ
73/8keqxIhQKD81rKcuBD19kl27MC+VWbsSdy9rllEVLL+Yep/xAkatAN/hQ
Dw1/oAUTBn5w4hV0dm/ImitRdiLvWj4IESoohrdXs+jWSHlc2lIlHEnQzXSC
f/Y8/lMDIiFCP2FJnAWcqc4oDyLhyeuYogsTNAze7OCX1CbzFi1J+uhF3ZAa
YoJQxli4SX/mT5PrtQ30NDNSLH+8VtlWC3KfSV+wozLMAp1Cfw7KQbZqWPlS
dihvBu7S15hwQ/8ZJ4fZEdIABrBq+U/z2VcFxiVk1TGjH6E29p59pWcB7NWN
go/Wa3qbzt73CWdg7p35PumeISUINTEPL2mQA0KHJBVXr0d5eJdm4IMat1WO
sZPlNZHzGsqZll1jo1FgxmjRGvsBsAckbIozFxvzmSlVQhLyv8PW89wwca9H
/KTchVUpSyqFMZ4muUh28s+8yu/f8RL/jnR41vKWrH+SHhRidErcUEa0huTt
npbsmB5i4ubOmPEcgpiguAezr8P0Mrk9WoeMeR2FjyEz4utTdVrltpQ8m7eX
zfqfnjmHhdUw4mNW/Rbe0XaJLLUlDoaHqdGA1yeO2ROjPHKnPjILQB1e0Jnv
Uaw5Udt7618oRZvfDSZ45467M+HgN65kW4VcNaukV2ALKAKmHJY9nZ88tRuS
q0goWa4hZikGACuujOCKbTxA+hDagzUoen2239pYe/6AwwhpkNdvax63hXqt
SFUXn/ii7giaFUkd75dFJYSK2nUY+7F/4Em43rThxUy8fLsRz/GPTpxln5cP
lioAjkXgrKuqLKD6tcSrbt63O+aJ8/daoyTSZkRVVH7jLT2yf5wq2F7oQNZ2
M3P4KM+dRFT9nAsBLF4WNsGAyNqa6QijR1IoApfGUvHe0QMvXQ5SuPTdcQY/
6f8GyLkUiu1eIvTdZOVVYyfq9mlBEbslIXVVX67zYtaynYJ0jWUaeNSeMUZH
e3rxw8bCTcZx/dnL/kmzOaZcRHldfx54E+JMS2rLy7lroRsRqpDMfU4Asj7Z
VS/YZxMtE6GM1i/KiyMId9eRjkzlhVZa/JKgu1DfxXlRwrnfJso5uuk/Ym0h
bmsu/NwjImCo1fbVdOWpXPU63R/tF2FwLur3iUkGvpudaTKsS3o2yyOeTWlz
pzc8ItjZmOpVR9cIi9i5CNMzxX5k20FZVRTbgtgCGC4IfdpH+FE+eAX1xMKU
0B2l1+u4ERrpO3hrShN72vikvWe60sDllLphAzvhM1M7tpvv11yPD3rjIfWb
N77TjRIYw/Z8TPZXMaVcPzldyuZYu94i8SnzwYZe9qPX4u2/eO4qVSQCJVn7
jBzfiH1l7Fboxa/RIRQOi2HpkI7Wmu4tsRtQOIdVt8NIGYENTQDU6GcZtwpl
Lq4I77Xd13X5cI07Ri9m7gYSXu3nvZxiQ61KetUp0nTQxOXnPmPfGFmwOHul
lQ8R/xRsKjcGNmSmjj1HrAYTKwyUTOGy2DezAAggCj+mFDtGhjnQkz9qEfSu
u7m9Mm3/BZnEWNDD1QU7zfi7sHBHReQ7B4yKy3dSKRWf5a8iRJgm/5O/gMZ8
0SLGuWvFGsqgIM3z0SyDeTDJS8RPyE3Cn4Yv4EBXSYq2Jrs7RLqmA/3oA6Iz
vmeEbXkKr+lf6wONW2ZJCOQuqECOd98eUYQ9ubmCJbfXjKXRt0yULZSJpFPi
fEdWZYwzZO1EqAyvKp4bCTA2kL9Xg9pH0/beb1HrUQgeQ8Z6yPvJ3gZmj5x/
+gqZlJ0GhbEugIsrGC2qsvjPBiN1Nrsf8YjBIGcLqKHvxwmbmPqgn9IXQfcb
MreDXwsgUbKIXDqlH46Js5PvQKvvlOCKlxghfQ3aukLpg8bTGQs/s/RJ3SLh
JiQfXBC4wotTXgbNWcTqMirFfht3kpPslAT3oTMubrfYCMhN/LsYVFRMIQGE
GRkbjpU+PgY576X+99eGwcTnC9JTp55btKskT7Gjd8jCJp9TWkZ0I8NQFhme
bBPIs1iJbpN0IWg9pB3ZKEiHP4fpPmmCWgaB2z2+wsxx5J0RrSiPG8xIuxlh
AQsADM6qVDLTb7ydDr137S/c4Ha26FysRRaJiI1thq+wnk8gca/pU+Sam8yu
WIdlRpGugud0S3Ral06Z85r9FY1dPTC7GlRqdzNhbMxopCjW7cZvj+XbI1gB
o+0QeNVBNh5B/O6nOaoWJVO7OHGZxCXPDPNMCo/3Nl5MUkdb3CXajU3fcFoa
nt1t89El3yNpgaqzJCWM1U84zKZwPyxdzGrscMwGjCFvtq/pjthbg/fJE3LV
paCG58qG7cfqEs3VPAbd54wnWXY8Ih6Vsb5OetKVm+pS99lm6s7xViRSJzMZ
59qJvWzokDaYEb7bF3J3E0RpWF8kmiMgOax3/x7xOfnt/x2JLbocEEbcgY/q
ziZg0220D4F7GPQpr8/IlCS6r/YggnFsv4vXqWzJguFs0IJj3HAoMw7OlobV
yqZfp4oYC40jFvopHkAOFd3achlmI2DWtCbnZDTx31zALFVfBBWzylK9nDMu
s4UhtmQAybYaKo2YWkulj8ZM+oLAdMc830lQ9kGNpAkLof+eugpp1C2y6Fn8
Fd6+LMtCh4Uzh5SWN704TwjYqlI0kM+6kptNnnCMVpTqjIuQ7OfZbg5kDqui
tuncBO8L+jvxrQgFtpSkCJLuCUYK5IHW7astm3zS9JLBZVieL+JnnTuDtdq3
mkOAmDcE5NeVhP9hewVy1CR+hJoTe+2NjEWM/Gz2yXh8uDgck8VDwgsomPqJ
BzUvHRCvT8tz45Ta5t/Rx7pYP6pekOcr1IIx7FIvoB0gi6g7P9txhK0uyIp9
gtTpcaPv3X83gaSE3yRTILHsL06RkU0qvHUfTMCh5m3EJ1hY4HpWrtAhqkua
FueVOyxRJO57ySpCiTk7ZIV/HluLL2dAksn8GM3ROdeWgJu9pCFzrvPuWuja
aKbFdte1bnFEXJ6QvcFeF6dmXmgYFqj16BC0CKSldSMt2FwyYNscj3W86jOc
qeWA3fVT/CR+8W7sDCQ8eSjMC3Q9wmhQx9uOfe1JBImTchSQIfdum7rUfADl
DRWc/CrSN91DnMiRPwoc3d4BvcR2f7e1hxlp8aMj7626wQh3Agne1ODTr1lp
ZV2OhZRjZ+/Nl/U632Nppb3ZkwKSXODOY/m7BXXHe8ooCThoAcZCfj1BpgJB
mhDPdZ6esCMqM7lm5myLaiqRRH8ZTwXifVxF8FYDX4DWaeIaaVMfjmX8PFd9
GavmNT5h1ojem3JTu7dIJmEk39Pjs0TzsLWb3qI/zgVJZwuBFf439+JafSXk
ydLiXskLBPlUEoruloY8gUGQFUhX9bKeMXRiFEF97jpAE//4DlMDs6IVU0HZ
iWS7MDY/MzWnuZsxY6yJ7k0qPRdaK4EynK5mnY+Z3+gCY8wQ7457DdeV2Hgf
L1UpdZ3LkKaJAYKXtjDwIKAWeYYc/h13fTW1O2wY/bSr7dyxytndRx0Irn0J
bh3OcGC6yPQ5LQ79JFcLHdAD2hoEaQB4+4ikgqrJjGUOrRvU21hyuTxdXmZd
+s1vuKzayBWUq5tFK8oacT96l8lDIh4s2HCpbTTSbJJmWMBwpwVSuf/FzXBQ
f5DcFiQyE+MfuPSS+LQ4Bsy0d0PTFEHaJGxIf833ge81ROCzpFwrV5+QW0Gb
fr0KRoVVCG3Y7kOcE9PFPISJ9X9sCqi0rNHzbKboTbOevX1QElBFbKL4Zndu
7pOdAJb44LuDh0LWQnIdLQxGz3r8modp0mgH81F44abmJFuQAkQ9m8FS7Lhi
/aQ8UjdGXnflpPckrQNxq3IyR1zCK3G1b4kbxmxJAengSikrCimEmHyZvu+l
bt14Owuy7jGe7Z0Pf4mR1F52ZltPyUn41DMwUI74Ys3mgBHhBJULkZySXl6y
GPmXokwBeWNbAEkRk3WjIdS4O6qPkCIOG0Gu8cbbG8Gxy94TaXxkYKRMabCx
1c7pFFkdLwoD1bx/SWf8zt4Yt4E81egAVgWzazjUryMh9eAojb46TKMZJVn0
/Ji+cKopTF5TWMNU02lkYQvkw7nHjjqWdlrMdpWeA6wQViTaNGigepX36Ent
Qwyp6wymrmnaATgGNBZnTcntILTZyPCUOWkM5C0JZjFkNnFl9f/PNqNVmxW8
cdQkZY3mCWUjDr+gUfvm25+kZP9dwZPBhbp3YA1+qf6ZoZXKZzQO7YDYJdrc
bErKlS5DlrBu50QHaL5yjxCDrdPN/PBXwCyuI7PRTKqKY0p1JygfHozV++0W
fUbSd6MPqmvQ4wwK26ho5p5Kbp9sEDLd5hSAqCyirzJ9gcgEHIUlSeTt6ZZK
CjtYCdIsszm/XtdesyxhlxL+ei5YUiGOjYa7pzgbuGIkBRVrGfGPKMaykd9J
ykqnZVXjwRGaAjhLM7XQf+PRpr6b14JzcUhVrzrzRLcEukIWwKJKmo11rSy/
CuSFgQGtKfcihFWnVb7MmIDLJHBOHoFruBDuZYnAIUxqGmFoD6RB3/cQFJhB
8sx3fpWBm/dKnOKVFmbtx1yi/DFXFznOAtZXHZX+rKEC7pf1cASvxRn+Cz36
t/kIiAjPLm/PujeaoZFgmKZ0VMcspgN0KI6nkZR8v0d4hz+uARauWbM2pHLj
XRtAyjoH0BCpZgSFmIqsnNElsBIkVMQfP7jaL9mQ1fuR7C6s98+bFbju000m
Qhho4NfS7Ml2huANpbThw3pUKo7x9PsLSsR8RO+wMVKYtwu1Ij3Kjt10ww2i
WXtOUpZCLEVOKo4LF4E90DMUDTg/t7jDLU2pD/fqvrlykVzLOGOac6pZUP9l
zHmQejTuJqrvFi1NPEwjpQlQsN2SPLUuecmGRaq2oeOT0x0JWW3sEPFPVK8B
YT4wIoI2SZi5HRTIU2VB1Vq/0h840HYnGX3zVjuZaihUt3JivfVgd5LmFU3+
FdQlo4JMBDwAHlDCiCQaZOBtM//trnAY4sdi+N32msdNTJfMv4H+kAppVmtS
2UfIYvD4Z+ONWyzYLNjsjkrIUnnFG1FBPHSGHI+Og5baITdn/e8XyC5Fbdvn
1fFvBB5Lp//w5jZh5vDA1lP38GFNQOfR5DhDAfIDCW+0U4BohxrjBGiEEXDG
nBbkT6Kz3bw1s2cmNsCe3yNbjl5fd1SzBQVIfi6xZVP2Tp4Rmsq2+tIPeXpt
aRPnQBChTJ+8GQV7VqryH5S/KYP7bxJNANKzonczeYzK4fP98MAtf0qNTcHt
1BPNBtqWzKatNS7iILdJkUFsUmqisUvwDA8DGfpO8Srwe+RIWKgF3M5E79zr
eGj8Gi2OOTePbrdygj28w4HGcZdiKJvoEafa718E99PmTZlYNlFH4YVkNmsJ
UooPfNiyjX4mBfCKiysFwsL+4pEWevk2LqypLBLl6LUT/GGS6jGaJDLdb5vY
QmhL+U+/vocmdMeKQvUDAkjU7hID9T/GCvVAgO3Ah85D5loemc80/y+HIErC
S8tJK1B9fqrMm5G0jy0PSLvd2K3T+ATlkY7c9U41DAeyyJ2QUCsvRGB1Chf7
6NSl4xyH7IBRK4mcVyXD+42VbfKHlgGfkdfeh2osZ98FT5GH5h8aX8GTRkCG
w/lMLIHbdG0b9mb/6Ot0eJR2d51EduOuKvaQxzhKefPI103b0kc2UeHGoI5J
q5KaD3CqhlNNAK9mxU7Qyw+22vw6i3IBOxJhQsYEInsgU2wACGrC0yJUr/sp
e3veZQIZXb+oCgvkLI9CzfRENuU06hAo0qWwQSnjr/bMv8y/e+Mq5l6Q2IaH
U8PsnTcPShHDGGfbV13YjLuBTOlc5ckJD0foorTlQbVVDySnw6qK1X7iDaUt
9BgeZHrFXtuECOtzSwsLbleZuy4BpS3i+DAJmdIg6DOmTqd1JsQ4d/O8+CeK
4gA1KpLIukv/4n0YhPK04jqxRhYWek/QdactNXR9Kekb3YXLDn7dR3+tMkRN
4NK/KIsjrojZhVfFD80nwk+3QcsoL6K7Aq1rnw0KeqmrYzHpEk/7lmD23STk
xsG3BfNSWoss5mJ5CCc87YbbNAVO486dKF/FGhbxuGWQ4J8PaIzGA791wOM6
YVb968rhL3qqjMV9o6kqW2u6YI+N3cuik9lmdXZFAYd5x5NzFlNFEpv9Q/zd
aSQoK3O3Amgphbruh3SKj3oixF9GbXqg2bliV2mLtJ1pdNBOPTQ616Nlq0Fb
6usQFBa8TeOq5BjIhs0fP6ypJAsUo0M+aZi9iCZW3dYWqCamNeYHPSlTMZpE
VqI6Rf6olwfWMvSyG1Y7ggJtfndhXtbV93o1lWlZZbnm504Q11C+EKT6p+15
i0WpwmI4K7uK6J2wbcxvc+5B569KgckfbLRPAt79YMhdj2HaapUpXO9y/dfx
jW1mAm3jt2OYR5yE3j+9/cXUaJMJrQgCj/BfUvla1+EfMMKEu3xLLy1THHfX
CE5xj+j8xy624pkcYgoqOVSPrYMMWZT4qrwH2wQKF3QflmgtebtdJHr9cP5w
Ux+XlVXXUiq/YBbJl1bimWR9rdUzM9sNH0A5kO8JEq2LNbqiNHNlFpR7W7FG
5lqPn/4zOlFdorNUghWUcylP0aCQ4JejNtbjozABeyEVM+utdeBZLqixEuV6
+NNjP3d7PVyI2bznmObhxhMBHzbHq1xfiRMXeyRisrAs7Ds+/hSiRkE9AuOI
LTUFDxvUsTl6tGvX+dsP9wqAKyfXs0ikhDtg3mVa4y0pWM3mn40c7jDvILbd
bMJj/xABww9Q9LlDUBMB+b1oX8+7t5+bTDw/L+OvV9U1LzuNOoG2Rc6FyvnW
rmliE5N/Pj0uJH5GQEI/mDxQ0cEB/Den/nVQ4AkG02AJNP8Uah5gqg3rccEp
vbpPf+PaLvGhCQQeoutbN1fXtkUsOMsXOabX5dR1laxXM9bSK5zZuv8r+Gee
ISUUI+xqQQbMh/QdeMRtoiBW+AVk4T2Morvz93aMf0EZYD7xQlWwktdwnceV
diDgzSOt6VgcdC0SU7wu9SilyrkEkGw+KllV4bRQCN5NgOY+o0lmH35DHFV9
GTIzswGpHQhHivopwMfftOBGZRMx4h+BZkX/eA9Vkq24wiur43foyUIxv/eP
c0MgGOi6GFku9RzK2mcwlqY5xfBqUIA+toPrlHqm/FkOBugai8CNmQxBdJrN
NURk8vbdTJFiaFGCBtlcVz00BONks1z2jiMiSXt2DbEJ5h+3U4qgnqNDPgpb
EBUOVZ6BrJf/74BKeqW4COVlaojDun0YwW3yMQW0DGjdc2Ij0KF2B1XT6sjO
mMvjfFjL1c2RtmkBfv6TJfGL1Cer03QA+PD10ZS4YYgem/BnpZNSyD050lgP
fAqa5cj908RFJoHk+7Yl6Qz/roM/6P/huEd+ZWznWODJ4X51p1nt0bn4jAVu
Dimza208OEiP26P6tg8AuCh0T6zm4eSvGkgVnDyIlteTCRL2XdjWpydkwpjp
n3oxdf9qPuh9bspvZ42tikAjRHmph94r37tE34yTg6XtLZKdf8mfkDV3fDJ+
zdkfNY209eP52LB3PcvQGV8ugKrywao0Stg4M4xpTRd3zF6TSegcuLSqOY72
oAkIiNYxxDjuv7HtfylkrneIl2OCEQOLJUd1DHzuS4qeL0KFqlSNMxJZNqNS
fmo5ZlxdoRbKkibSipqE32gGWnmnzM6cYKpjH+NkrawmQFErOMjx9u7JNiZ7
twYXDZy89vw3Y4JhH6PsAnwFXDCi+6JFdjzSXnxUSBTL4GB4Q2wRPaHquTuL
9Zm3/d7mM+c9qYh4WLXseNMYXFVjHetISIuo9JzvqRbsQE8+IrI1vJjlyimS
s64py3Pdx1vIVNgChybmMDa5jVPlBNQ5tPNntKpEKBTdlKQB3Utdvo6z41MT
Stt7j7a30rO6dKUB952jIX0AIOFexxi+ER64b+zxl+dL+2rUnY4HeUXja5NV
cUBuPTNgOUhqNlqBVK2suEGT0iA9jLEG5rHSI2mXtXUkSfe+jJQmQPGfEOlD
DMW2sKd6zBx/SY1QtqcUsUW1qJRTFSKOJNN5nnPqwHNBsQMg509MjyfaYD2+
/0K2LfIZY5bh8VbgzHutMYwvMD4WXQew63asTeHwCzPG43zro90dghQdkT23
VMrkdNcKWtXROAFvNDYkbJoQTdPfMZrc0fMsoJlIOAJpZWHYA3HKvJ4nFkHb
SLNNKZKTbIihwUl8AIIVFtkUJ8vUYYTzpdVhF7KthHfLHB+hP/m9cdB7J+M2
jUL1sClgs+3Y4GOgX7S8n6cOKX2me7O2vG416IJ9Q16oB9lFwEypUVcqBdr2
2NCZfIBIZnYanwA/kcTXtzkQQEFbJTRLslZdj1pHfPYw4CiT6FFyk1HYuC70
8LQHFMgwSoPA0Q4zCyngvasP+5OS2MruwiU5KCfSqYaPrasmpLWaB6rKbOde
8x3q0ALMvjjrn1gH9XsLDh/HKjF5np+3mrlM8FLPVgDf+tYv9N+YhmfG8lNS
fvkPKiXgaS6WaWbl64m/zvNES82R73X0O+nIpqjFo+fXqwOdACgz5dYiBXki
0ItPz6UQppM9xKkxgYcjwWmu9fYdyW8BOgtSR/r8YC5PtQKdENQMoDQZGLiz
RwFqTTbsXjPrv0p1EMIsO1IaU6bQYFcWMIgMwYjqU+4gI6448/6PUZZZ/8kR
jmiTjrGOuzod9jRNrMwR2RgPhUo3Ki11trtGGBCy8C0osD46CA7AvbRvyFrY
608TdszJCpMaBbi8ofSThEIZBB6HCWX1yR5Ughkscdr2dhcK0JlQJgkL0T2f
oarEBjwqJWDCOXuInX8NIU7fTrNoEEVNt9PGKwy7VnlLDmuWxQ0aEux+DnP0
FzIzQ7LxdcERfKpP0d1hTqoDdRK6H9Noj0t8KIF5SHGa0tH756lxtiDB705Y
rHT4T2Bl3ZL4Rt5F6Ty4PlrGt3rFv4BqohhtbDt6YeG2hlRolR0VxoEqcapS
l1UC3NGZl1/Bf4QRisucPH6YuYRZPLrBuWQf30iAXDH8+7Dr1U8P4W/n25Y/
Ql+VGDE90G5FjXo3EGBjfCm+LcpXGjw3wOQLDCEmemaX3oWxwDM3h24vnEBL
PR6SaNB4bLF++ZDq5S4OxxOlGG8ll7R8DoRFdVXX/tMVKOD83cI4g/0sOaRO
KbccVMQUZK4+FrNxHIOk78MmF7c6QIXzWl3Dx5o3esA4TD5sljleI0hXPZ8L
cJWFhy62uePWgmlsJLIlAsknn1RIqfs8RYE6QknJVZFTEcMYJyvYf99qrxSi
Dca04NgyElyncfca15Wp0cFoGP8Q1pHvfUOQPQl6skLZQnLZw74ZWJGZ7ucX
8DgYrCOcbjeOx61eGf9cgeTmmct0yVBRUijXH91MFtHDjRGaPArId3aCpSV/
1hUXyGlntRd+tb9mFkJ+6Jh/rwwGfK8Dmdbo5yMBOLocT6V0wvvWQJVDM4Qw
KkUhsPmF0L/zszmZ2NI1cdu7yIJ6IL/Y36oYGtyTtEDZC/YBu3kiK5Z/sr9W
40iU5iUVBAIZu+mFWYXVoIZQyINeTwp6kOvQCr3SYdycc6xeVeHaFhPqtYLO
WnOBUqcqKEx3KN08OQVavw6FMbBERzpm7YvEetgC81m/1dixFC0dfAU0bVYa
2H6jocWKyl0DETStKnbWavc4CBDW6kxR1RSe6l6VyiqvOEt8tDfQNCLZkzvA
usbWYcVUEqt15Y06ANgOGZuwwOyp+PRZpeCEQ1I3uFWwaKh4ToArgkAhvb3m
kuCPTM3eF6xvcoFsOoRSIO1hJCOxM+2qc2RJTlfp/iOYfn1TDakjfCZIJlJ7
P+BIvlaTFLhNBzQssBTDtTFFRu1w1PZ/PFqQbksf78Sx3IPTIJ47KyUuVq83
dyBHfCApsyE9/+YyKe1h7s1XxzLOoM0bSxrxB9E6nAoEQ0OyjQA6yU4oirU6
3uYvyxUYNJ/ZZE8i1/Uy4kuTJNcUH/yFk1XoQpu+ioRu3tLs84f8OfHR8NIw
l6EKN2iPELe7eakEJVNUVlLVcY6FgsS/cx/+gcn40+fB6qhcZNQdeQFEzA6Z
dUcUU5XkLYZM7jbGMlHJ9NP9WhosSo6PY4c1H1ySiSpZeqqfLJoZkQSk0V48
/NXZZH0BzzMz1KlBchXSAVCPDbLmDJ5mTpJwC3VrA/WiKUiLNHZxRjFg3C/T
rDKpzEUOESUk4L1daauXgPOkW5hDvvjJfb9lmp3YEgrzq5+vuoWEKpwpqY5h
ka4CUEWzAX93LLVVrhuvAPQ32P3nOJj2HGbOaauI5YS0ietnDI2HEOMomP+u
9NkJeU2+IA8NWYEDME992+a9DauPkssvVD4pgKJQ4SVyeRuqtOzrje7nIG61
zahIAgkZFrDnWqqTkm8UgmDTpwIMmcB0+fzkXdQ2TekaKsfPR9XBb9zvrQEz
5Qv66AzEAL2sVG/k9VtN1Y/Sv0onsGquiwtYqdK3Iyp4zBh9FjRgyb8ESap+
9XQXdUxo2yI8ZA9bwYx0s2RwcW/cmO8pXxWDN1/3b9exUtCsTXdeP5HnuYyI
eJtTxGsfm3CquxyenDOgYNMnZrYe39DMXne77QAdEwW8td+30xMp9qJ//iZj
TtbEwrUxRAPEIy4IKkiYhGa7DbHXoo7SoOFZ++DWdvikXzWEBRycIwh4UL3j
4uk1JYn99Z7EvwlrKS0ig3pMIhLlaCrVgVycdXSjcs+sc/md22kAfj8QVKza
+0SdWxhbDbu7DT1d1LIDm+2VEmYfPQ4KlOXcxcu6ter2L4f1C+pMRBS3X6hz
RrG2WOIKTiXYOG8TX0NI04OkUIURTzwNrPCbNQ+GO0gPVgmHLIYcbID3zpui
1faMzxmulUk1ZKjU8LC/ZfXI7IqE+cAugKdZMzPRcTU8D6GfWo+8zYXdUZz5
eB7VWNkIqhufZLv2MISuAFUkICritMTvicpoWMmqPAn1BDvPaVMFJRPvDZsF
6QhEmPfn0Huh5gPrEr0fNFlRO+SIEd6+tzCywMp7vHwj8aNu785FUeVEAbEE
3b2xQhCrqIjUJ5cO+LOkSBI6zpTSI4bchdU1r9IA6NPIQ0jXgfLAzhk8yDuP
u1ipf3cM0pU1JaaZ4XE6CXLNWWAQYBFKEeqqB9QZ+5L6+9shHEPTsv2ERpmZ
6QRnuVdXbuyfNGvY7QPh6te1C6CbZPxkwd6YNGF7XWgAx/10CvZSc5NyMCEC
JtXnRFckmepkYk7EZ2ogcFH14TT4wN+41GzxJbcQ2H/pGbjOhFa135YsN/1k
aDeBF0MRKoEkBMpxc56R6T24lT64ed+oKPQA708wJ4duIEayaQ4sNid5bnhh
fsLLdU1RFkfJ6Icu8bhh7Oqa2j7zLWvNU+I1FCULhBpohXv3Nu+mxh6DTD76
O0PxkQcpy5lr1KfgOu9oNMuIDt+T12rtJiGfVIq053wKyTbpcocFBiNw9o4J
Q67/0fkfguEjZPwa2hf5lo5QYmU9/V9rCvSkdBDN5h92Kkld1ezrJkdjnDuQ
qQeTedPQiqDNrXqhBLUxonLZq4pRD93K0VsEX+E2yt6wiC58DXe7Oh6/ZYaP
iPcIT/EOMLoAni90UgBepWG79Ryh7xSTZHZ3GkSmZ7Nh3NVMsYcd6+rHsYGN
l59BHi3BEJgyDKODBLXv/yGIqNvEOz/kOCJLw0x/bbfP4WSKh//L3U4oKm4l
iixlF4fnEUwctZ/gAJ8pb8Nu1egDGSNN56mmtE8nfj4Das7Optn5o6NKXidO
4uSZnX1zSmHH7JnkcvYj/YAPbIXfLFJujdTi7HmZ5RehHVFpPIx9u3tiM3Eo
zJdbKrxztA/x5h42GavSd14p/zRZwkq7D7OUBReMorwfVfYTpwM5AXs58Xbh
73TL1ApPp9tts2c+sTnToxG1etcTkngP52h72T5qD3I50KWKAWoiWfhQNnqq
gjfcaB9DvnxisSiMIGz9pkKvDFIIbND9ztrQ0Az135uMvDCFXKs1JeIoLZtz
FN2Hpm8mViRPJb88pvzC7+pbCVuXF2+1pqsp2yJaX/Mlx15E1BVwB+Tflkua
1oe5g4NCS7XeOVrvdB9AfhfsmpAKX4neEbLgKv7Ho9pwyhg6LgIJv8yXs2GL
Y89BROJ+uRawg+pXV4Ci3Ws3ionVDVI7RUW18bYxakJkdpO2+Cnt2hHotZnL
tdCuP3ofHczPBgs+D4+QvGIbguM1C0uTaPchlRQSS6LF3MG5zFSIxbu80iJ7
yTiIPrsUTBHqiVSYYdvqS/PjxkMrsHoLARZbuMOxZxOjMbZcEXLZ8pGZPepg
uybzZdpFrXtBI2cDGsAm2YfD9/G97sHKbge9R6QgsMvQwdJgIpkfHS3/LAXx
UWdDqhjA8GjAjW9SYvGsRW0IsjmUG3yCWLOkzRohfpaBwMNJq//PP4ywdKs1
1BouIjrpDHGhETe+PrjSE39/jl264VscWln4jMK6dIPNS22Tacqac0Dyun+C
OQuaSqadf6wvVVAhHCZcS5NB0vCaNE8pJ+9nl3bTHriEKFNzG+5KMQIm1bjk
Gu6Wvn3ZY1m+Pg2jZC9fj5cSjvfX8QjubcfLyatSe5/gOe90h57iLIeiwDp/
LIXBYyKTH0c4+xYIsDMwaZaqtFItzhTicE3DM6dY4wUOMTmGcpiX3vEQ2jY/
xUqpA/gRB0k1lEZ86NxI4BiccFHVfNxBqu3sEwyU0cgD+J6BTINSObnvNl91
ffxDWxHVXZVom3/xkBGan+zreQdXxKOQPH2hWwjZmnLPhup6Q3twVDJpuKIx
r9ieuoKQoj9l1oE4f3ixCDgn6KWsfNYMr47nlGwWqzcdFZ5mcRUWxRtPL5gF
QQQvJzNXH55EYuJREcYXXoujmEwcw1kZ+s2tgWwEsCyu3fv236AJTbIfxdHw
W4lvOZ8e2ad7RI9j6mRC13fXhHiYpW2VOGHz77/6iIC9RgCZ/jMljyazTsqA
4zyGtWVXgxzqHntbTWo9vLsM731k8eGMqlC0RXcL0DEsIxh/wRhhYXgJthAq
cMTFZoY0lX9y4uPwFXj0inDM220Dwab5lQXrgZphTKGGZwcXtTDygtIdkdFX
OKWdoCtqpBeo79xf3l0jL81+CSRaESBnC1gMnjPzoIyVwzeCPjgZwNjrno4J
ZlMovQNVQdoKNy+cwPvGuKv2WkFYYHnV2F2WAs4PPFTlcUIartF3VHosFBHK
sON42Zr3kLt4rbAkSn13WA3/cKl4GEuD5AtkQfbwo5HOQln5hwwoLAXCRl8k
7AQjouC0Fjp6pSZD2f5H+D1Eia6kdPAdR2M4WbiE6f2uZaBgWayrMXVdhh+z
56YKFpEMqhD0A+d/m9fhYE5VHO+h72WWEEblImweQVk5ZryvbOkQHEckzqzH
A1HQ0q95h8koJmZX3YcBM8Mgt97FpY2uKe4wehQzN7nw9I63akNpYjYlZp65
ximx0Uu2ZFPe/x1rgErM/xVGS2ZejJc1bjyNrRH9CFNx7+BW81OXPBw/dFKn
klyAGNuhWSsW0tinY82fJGFyUoyvgttQFHH3z1z83fZm0pUg4arMGKv4LrQr
d3zESDhJ6I4aekbhYXaOcGOOzN3bfoQDugRXVjK+PPhq+jl9bczC8Z3AxgXu
FNlw7rZ+CdESUZQ1oPHlk3Ij6hGmm+S0jwph7v9ksSGy2RgGcxZqaU4OaEMQ
EcJf6wkRi9kVyjc1GTRrpUE6hVvOX9EOIES1AMd+L8oI0QaQLygcOB9KkPR+
OOEEtOauZGVSNPlZJwFCBMXaEbKP7ok1DrHvsmpIWKbYTN+Oz8W32QpM03GD
7tRuXPKkFJTXtXUAo9LycSQ4ohfJHizgo/z5vonTQDdrdaT30TFFdMMbPXWU
XD5hxsfdPlN7+DDceBtA9KwVtjLYjKKXROxOU1UB/lrdR7TRsOFH3HHdq/Y/
8H3Jc0Fql4KBGyoNEobUgOD6b7R7PrZ2N63mbOvI6LJX8G4kgfR8S55n4WnK
9C1OBoK4QjDOvPFUfqqid/xWwM8xU7sGTjk0SmsvLh2Ql0BsQ0J7AImLGY76
vfhYYqqW3+xTW1bPYhYDJ3Cu9R4y6aD6FW7T9tP94Kt2pgnlD3b6iFubHV3S
V6Fx9WNI+M7XUW66phfkXKkt58usf7uCWDZdSB31EnzdAWufCKg7eL06sk8K
7PE2aTgwL34G/TauwjRJrXW8HmTdx9A4YVc1FAxKL5xpNIbLc4lA6AJL9fao
PO0h4KoHxACLe4IV1OQo9iPtYPruQg6iOkJ89xeOrvTrIMJgiUWE6AD6CXf3
ReqAuAUDhxemtCFTKVtuzC4VQfkQkrzuA1r52R4yYg3Ae+i9JU4TwZRan41T
4ykaBpji1CaviO2a9ApA/oqDtZG/IHLf2rQ5ZUZd9k82PujgtoJbIpt4O3Qr
nHNEJPUIhbo8bZC1VwSS1IG0Hp4jlYcF7OHyO20WpsmXzfk+CWSwVlxQBq2Q
SeG2bCakFMxIfPvaNVTidps989dvAK4t9UnbQKyaVDqBt0Z7KX5q43wCDN/R
xKgasAyd3tpDaEDhzHFSfwKc8gPNWbOcab8Zj9FWgFFZ46LEqc0GKPL3XUQo
qDWLlvM1/kNKx4NdC5OZt4VE2cdY2N4Z5DmAQWQmU5uEXK206XSwfPOxM/jd
SNGcQhb95zecZ5zZURbeF7jzTVPwLBvZ6+t6YkbPnVG53bcj0ZRJ7m3ikHOs
eBq3cEoUhhXrW4+BOj66Ls/RDnfV2DOSWzxk+jwPSnWO9j4xgs4tFuiKq3oD
qZfpGxor2HM5uJ28SqbklVOTjtPIrshHBRphHEgBtN9t6EkVHcSQ9+A+9sHr
wUPqX7gPhFqAQHbHumvXcXaJY5uZhmbv9s5mFMQbvsACP0P1uxzkCCQDUH5p
KXW5Ly/Fa5hZSe0o+aC7oMNpy6uHB2dfDVm7rmej0wythmW6PPO5Q7dtXmSE
kRXulrEEQmEl+y52SST2mIjb3JTEljgo9z/n7tBlYbO6hBGe4phQ4ylV3nxF
yPfQJke1ZwIgbpFBztPzB+KcFTWq4fITpev7PQFZyZsg57FCkQ/fg6BYKnXD
uyzcGy2o9XAmwgRVF4KGiGbRsfMeITp2vi8vbnBOyRM94QShgE9lHNy+UGKb
L6nH7sPZwonvt/J6hMFV9bwIM+T/GtjzBmQFnzulbesum+QJ+ovsKH6yQ9aP
k9IdImX2PN6C4tT5LV7jYCueqtYkXb8sDYDY83EGXJ3wno7ZCKRMclnKR+SL
XlT6QzUTGrPEUJIq+wXiLbgXuoFD1kDK7PuCWDFKL+cqQllOF+35klIRmunl
AWUmMECr3oHK/LasDgvhKFzSrz0dS2Z9ACFQse/xukO7IK2RmTgC/s0J4f+O
cEyYCIsrp60dYHE08NEJQeooaYv1buerS4GTgnl+fIQuXts5Fs9MAoyE9apD
exQB4HET4CuYAv2kMUvqH3/aSjmBIQxxNjVZeqUwCvpiFCmLOrC1+Be6/Wwr
7HPYgTOgFqw9tMREGtiy+3YuPHbsq1Un+tWoYrlVBXqbAGqAea+ykFhpqjs4
8Mt/bC4WYo1X7BSVYvqzyPuW07vwpi/XhWEZNQUYBqEdp+ROI+hReQbNI48a
bsZPMV2Sn/YDznJz188mBufKO52/g29wKr9+PGDwfyYyKD5VDQVw2HlGUvt6
/b8PV4C3EZda7UcqE9FENJVjMQ0/BP9x4h0ZqZwKtlAycg/rLKUPcbuSOtao
/qdCHQ/hp0cnhxZilQLzkDXxQb5JMa7V3nIA2+7sRkRvyjdgVhzUmpK89+tw
9fUgXw0yGxDM+BJQwOXnDA08l7lg7Rws+57dZ8W5sz9X31B7bGkGN2lZK5Ow
aemgIOa+K20nTsF1tfA+qtgI+t0Cz378UtS4coKRVdH30e8RyHC0qs2DRuVR
UCiI+6WwXwYFJGKaIMzi+RK+iCNbS1DWXsC6BTS/SUwvFqoMwS05/UCQ0LtZ
4gwMVvMpz6S39jVm5TtMZY7lXStLS2QeCwdE9L0pPvg88sFgFWqh1/KjZuz6
KXKPegNslZg3Q56aA95P6XVDiAOWsmMP+kn7UhoyYB0wzZwMoHddwBDiWxzJ
3OdOMelwIgCUHS5x9ZPUIStt6AAlQL6r9bndIX0j2qaJY/EfIUyWwyFVkrOo
/aO4Hok2x2MxOpkN8ykj6QczqoAdtzaXjbNCjIPslVj86yBszc+rYFsEg9py
jOslxwmWyu36otpouRfJSVp+QgVx3v6M06+UQcbtp3ELD0p7Xckeirz2SQaG
GdnRjtJkPptOOJS5DWhtwfmG9lStw0YUoAvylrv9gwrY53mbF241/FNgbtae
x4vABGy1ZhXPwFEllwCniPyM9CyPsk3ZOT92SvsOWQ10WcEqYnzWi/QugHKa
fQA+sQQGhnPX6sgxxuFzdlTroa08AaQ7PnbTTIJHq+BmJu8fGNziHNGmRhiX
3AfAgxWe1NqzPGoup/eYN4uRWyEwCJyI9DL+faROWDa1Lgyai1QI1IgW7wTc
d9evXnLFOYvaubCb0glbvzsOvZfB6CgvXMu5cx2jqby2YNccLILzb8pekWKs
4krYYsLzdnUF95VEGQuYjmvnq5uwL87wLf3yO9WO/tPdg5ZZ/fFu6GfruQGz
7Kcn6oxoV+avqKO6xi1fTcgQ9Aw0javD0SSRI0qidIOOuhEm4gEy+JVKN7P1
8FU4i3FnTBAbakWG2LJfupRrFLZjyrqJPmZQ/YtqdzGeT/W4ZAb1XyGLCqI5
SuJgVVWVewwOwWSrkEdbtZ/Qg0l8kRf3quSxXXlJZV301OOzX/MpYR3j2LLq
MAKfliY8bzQk84JfE4kNjdCbKJJhMGHfKTVYjUArvE+E8cye8HSQdlZwV0Ez
j9Z/crIdeQyevhlZYMh88626Cq1g4eNeHGLcjpaVIi0UXZ+POrgWb2CvjBB5
Z5N+LQx5UXHlw0GjXuy37lYI4nW88S+FbRE3KVudtHjWd1jCSo1BPd8bS78D
2QOAc+yACMCzHG/cUT8OX31wsN2q/7r7BnhVtMK1oqx0zzD1uCOfziUXRjSA
fP7Z3utJOdgo58j1OnDNwjitZLNVhKiteq/p/p+uGC5MqqOAmp2qllyMBxg1
84ZnedZxn/8vDf3ZXUncf4ztaF3G2oXLufk11P6hRnsl5Dz0UaGOy1aIVJNv
A/IjYLhBl5EvPBIDZ+Ntg6IE6WWajryESt8TcGbPnO17UQhhMe8wOwDXqQ/G
aokYaaveMOWlJdCm0fdTeVA2NGZK6P5ScHbwxRdiYhFDeTsjV3F9ecDzHJJA
N4y3GaZA5UfrJOi2XH6ctXfVLEYmrXFmM/yO3zvx0/73jX1n9FxWaEDoQ07U
0NxOJndSi2J/F5fY9A3lSBZchBdrh6cZ9SJ7KdzK4PMZSK631AcVxviy5/p5
1ZUNr/gO8t18UEsnGeHAGteOlCySxXztf2WAJ+R0z1HxHQD0vuE4Z8kQTw7V
9mxfawXcEctbdUMM1w9wdzp5tm4vPcAdEsHmUDsvG8h49pqRjvnHSoMS9Iwq
zM0kbdZ9ukFGasxhB1XI14SSMzamA4/tr5nI+UZOzVPiOG1KawiuxVdyO1HD
AKZB7KwYrK8Z/fYi93NX+T1bOgGO0PMjGfsw2nHTWd3StCYBjSBZbAMVtWkw
PvNEcnvhNcgWsFCLW/hA1TGQsULmat712aSiBusMy1yS/q5gD9PQZh5xGoM5
2/pkq7bwdg8+T9eZRS1sjV/0t2w9r3V0Zrd5B/0Zl+SlugBWiw/wmbZcm2ND
t1br7+yrzsCekHThTK1kfk/8Fcoo5IGWVtEMP/53rpbh7OGQy4JFak96T22U
I+PatHxy5pPmuLGznMFtn1U4el4UXx04Cv/5Iz6rohhs3lBWbLKAn5ECO2CP
QKXMc5f5oN/6TJHUV6LpGgj0KcacpWCQi0HI4k+JSNvk6xlSvGrNw+EwJMJt
V143cmBgijRyOykSFRdou6F7MMBIg5zNhw6JiodBh/ssKUUWj5qBIZCV6eGP
pE9aiN4MWJJ+HS6lJRMu0cpslWMs2X79jmNAI+JRrVqHaWfsSEuoC2iY/f2J
XC+uHE4U1iYTaTe3jozkjaZ7AiuW00nH56nrVNOuPTJyINwvE8rcf49IV/wb
I7nBtDLtfucF8xQVOM0wOR6U9v7G74NTwqlLd10dq2x5vuURudpNVdWMQ292
Ow796JduZq6kaVZaTPfobIdHPEE+bg0huoVR35g6TxMdY4RHz2De3rYQ8q08
18Oyg3FY35Le04iA2R7Qp1QnFe/YZTE08qEKvgEUswZ8WjXshgDfg8pqgvxH
bn/X2Bdz+CBFJhAVCgzTrJCmO80c5wOgsCpmj1PDhbzKydjZ6v+Ru5ftEP5N
y2Zj74PusJjlnMSQBnP8hwSeGyrbQePB1sJsowJTz4ppwn9U8of9t4zNCMgQ
irauWAfalbOT2emvfpq0ub2cgT40UjCLLoxAF5cpv6xknQIimDHa7LF1XNyg
AQoE6ehjGWgHat+pdW2KaYfxRJXPPRgiQnFzlDEfjZOm5yGxkQmtzkzrWNQn
MKPL9mEIUGueoSLGZci3raJyr2ljgW2ai8Y1bMjb7bR0hCd/EhG/A3SdN7xQ
Km+AyQOOLRBqtlCottasH25ldMtbz3h/3wzemJns3CjJU2gMiQN5/Jr6Vvxg
H4DdvCPWafqS3QT+BYuj+Q2CG6MzkiNLsmIYKyUuHH0YXCc2HLWkFj6dNw8V
peSwh5KIj7NjtQ1/z38N4DnlwuiueCS7M8DyYZa072ONG8RMIX1xOpiOHD7f
1TBDckLqXogDf3NArILZWYelY5Ub0M0R8EjKGWYEsKpp+Xa3qZcvTvQXrWaM
bPzTMY6Dvaox/HH4O2+lo1E8KhKeZ8lRg6OqT1FRmEqwQps1Uaro+xTNBB5b
NX8SxNEz2OVBIr4GNczKs+gxLZpHYwKTnhtisl5ij/JgCocpx8yI16umtsyN
3Hm2ST051nrhgVR9DiqUlbRW3pfkc903cosEFLgz0oP2QtWkNdO5F/YMH25u
ZXkVUtTWj9OMjnUPoNuwS4SuSfKIKfdgPrFCG+X2CXhJnT1aHxaoK7I6Ajc9
0Znc2aUR/mX2M9+YxsNdi6bHycu3e5pXKrauZbN724rtBYriWKUxB15ekT7R
QMEhykgNHrh1HANUqrpa+TG4yDmZ/fIv2scRNKxSiuuGA250WNZeLljCTmrH
3WCajFa1WgDvT7hKEcfJCwQdnufH11J/5sqol1Hwg9wjxw+6bAVsS+qDOHnP
ojhss6zIpYLCignEyJTg6KXjmB4eTQAGFJJf9ViaQEN8RUlagpBcEClVMy/F
7MtXBeWZwEemUrZPy4T8pSRSsrLu0DESz+rTYUkTo9w6EgTFJSwhuaDXr/IL
n0UyZBmqRbQjheB3UuLYGc2bi2bchPxwyr7u44eZXsTTCg/sM77ZPQeFVOXD
ebGN6GxF9vERPtuZzcK55VF5tulGZjxvMpvptvAjTlMLG+vS6qd5Msw60Mad
bSb0/7ULpjqMk0/adLBRtVVMmhM0sXvOK8xlsCDV9R92vaqtJ0IZdz6GfglP
CoIFpPbMypTC7x0lpVUKvg0s/ichblIQn/KUNOonwVpgb3BQusjyrsD9KtBB
50yHGW3w7QcDGPmJ83iXJ5q6/7KSAXvH9pSIpNGlXhOoJMFWgCNWLwbMlEJw
Fep+ePy22ekeGYwEodnrNEygQGW64lylR/fBjWfSwaYb3RlLFoFsojDy3Bf+
kJrjYGP3QrpcvyyLcgOxSOKV1CBUScb5PyvnpdKQAd2afomj8dRVRsZiHk6Z
x3BK8LwAwRoSUkmJdn7xf0aU35DXZe662fBT1euuiUltfHmMFllnc+itXicK
ctX04AfUoNSck9gpRvAvzjttP4Vu9TFyr2xsIMuYu68EZmdEteFQpSB5tIWf
JJA7u95HPx2f8awj/2He3NOy6jir7fMC0PTObraAaboHIuOWZRBbNEDlvEsc
KMtZXKoTTEiuQ6oyLLKx9KdT91jbYKEazAda90tzSAOUrUWZ4P7I5eTInEek
AcF/WMFqsI5vg1CmGY+rtJepK2ECmdmyH/9yOoTJ9xh9Rzja39MtpI3vgE56
ApEDdSd7yxF9ZwF0RXMgaPTHoFlTGHQOKplhtjQ8nRu/Bbhxfi4mnqZK/JgA
FyhJC1D4qVgWML7d5fsqkqLrvRiJmpeKi+6c7jUZpeX8WfRmXYqEVfUx6XzY
IBf2jIFhkJ8g3EA40+PIaz2Cs/re/g91B8I5QBB0DwJcUl4YikN6IMJwl2Du
tpfwWp97+iDNtjEP5GTpQe/1Yprh7w8gIoYPTw8TPAOhfRyNbed2pyf8d9E+
AHY4McMJMQT8tThJqt0M6S3D4qzOVuRdbBd4Jst5TxmFsPj3Ws8TsW/Yc5A0
VLTJQvyOI9564LQtmdxC2Mt5vFlVVQEYStMMReC1o0tBeoWBy72qBxY+C5bs
ePm1S6oBrLT4m394Kp4lfhkrRWbm1oR4tau/Se3f1+9tpajhEDGHZ5hSlLG6
NFmF+hgXeaBdeD0t71z28DtJRaVrsebQIstFMgaHRB81jQeSvN/aBpI30feb
Y2PH1wnJmCiD3QKAe9YSsDFHQdjRI1R/BoxHv/wrdMgMiRWPqg5BWupBUMuN
DtrVvLFjMhPKigQ2PRzeTFeLExp6WmGGNG0fC//tt0iXZT61CrqcOK8I6y6S
112Z01d7QH2jtHXzWIJHpFe4LgUt9XXztKT6ZU/bi8vaL14f2RQGkNAMF5uc
DjFKDS6zISyHlwRB1WgbtWgLGUiMZPMxpSjrqJfZpzMY7vywB0eiUjTbX+ha
M/NruRrOUIfodw7dJ+4oNu+VWa74G9mHgFPiHY9ZkEL8mmeTkuOpL47fMQgJ
cAp+R5yhLP0jo5wIRTH3zfTPc1EzuVfr65seMmgFKtNwWNIzhhQ2TjH7a+cW
eGRJoe4nHy1Q7fG7EL5Lmx34h/EoPvphtA5rewrhLR2w4W+dVCcEl30OKxhg
aPVqdnKo4AW2X8b2nGw8m8yQlKEhwuWeiZIyRdNUqzNMUr4d8wrB0DPLuHxY
TtJUqURzbwD83MkLL4iVNNNYh1ellYIGk568rsG2fo7t0OJuUWN/HMz/zSTj
Tbw27oxtAVmTaQTjxHA1Qys+ecVNDC4EPYLp3iz495QbLVBH15GQrhjb4Gsu
x/timgIuEc//xDLDyACxZaaXG3xafvNhKD+YCi6MCvn/3Yh7B2PmBL16Zebw
jI6arLRzl1UzAb5cu+uajW7kRv4liPad816Z0chnl7reF7gBkg76mE/A29g9
EBJR1XvTXcxFXT3eOUEziIXSwVRow2quZeREgMtXZcxnyxMNgNEri8W6wjHg
9bNyjY8bI/aWxbgH9p+7B6VfYstvyHDc3+p5pwFkL701lvISyFcqDw6MT+k1
fNvlDHqkZV3QZbOrLsf9eyAsiTahCR2JKI94IkS7gzhdBDUfXHCHlNwYbnq3
g/elFUpzgFbnkK3HnqhRNDWV/jTi6UE0/LsGiumBhJ05bSyA3H9mewYHqY7G
kMJ6K0Wb3lA8rldK+zER7iq6iJsWS3Irr2xrKRQGhHGIwCZBORprHTvbReQ/
MsEYsUnoxjW3F6Ym+240XQHfWoTSbkilK0cDgC6weoFkWH+kcqAjw8pi6QSl
Md+qftX5naoaGQNscrGPW2s0b7/ju/A788PQHmjWzlJ2OgaZnivL/KL9s6Ig
90UOG9WnK3+GsJkM30mrhjyWYI2ZAjo3ZXM7TvQvFRdk8m41am6F33pcepDo
sWnx89QdRFJKf6E3J+nLefbyBeEZuildLHpae8wshR+weY5milJBQBxl623Y
vjyy6JHy+vgcBW06mCR+aj7QEDePWMvAY5amSBAl3nEaqVAxmg/OCbvHSyVH
CJtxQceMpjN49qTP5vcDBL0Cqa0zbZSkF5aocXOgtE0JEdmzBZM5+o5130sS
YZN70ZxFBgM+LERzTI/4JWxl5QxxxEsmSaIb0LYG6ASF8Y1gLh9GIQLhnALS
Htj0/vgnzA5wYjnrv4WlFLbJN04HmFPTuPyNtJynqDKo+gptDLfnKMYL2J5r
nlWntfcpGkOX58LL05DWLHMGd0Mhz/Xot6on0lcANS5R7snsB5+onSudAT0j
ofD17Nzet8XK6u4hXkm4MqambA+Uy4bmU8MdVyU0Yf4QOP9DOv7sE+TE+KPq
gF++LMhF4bFxxgC9tZD59sC+G1JpHZJAF55G6LC40xfoBuEj7mKkew1R2FIf
wmUdAFgHjVi1PzratV2iq/JnDwtF+Y4WMXqVTqFmdvkmzyWe1bY13PW0tyJS
enxTM1cXf/jhd+f1aX6aWLt+cuY2qP0KNT4Vf1sAe5neHPugL4IB1+TsREDf
NNxUfhRkj3D6VbMzEA4y/KYYn2BvZJWm54ZTMwrZPRznLfR7pV/dA6GxW73s
/mYUQ7pvTNNilmdaN33ZR0Wn+cT3tdHEOdW+j0MomD5blphxpvxLBQQlnXkt
hzmdDAS9JNCSmkXYewQEYV59wgIHKR035B4sQ8Hy+6FgNG16TMaSX91uU8qf
ntrnI+hW75dWj0iZDXiMfS7TX+aAg4szGCJbdIsA5SqTmiBS2AALxTvS5Gsz
bvTzBHzCd2vv0D6yACzWvexRjdNzzlxQ9ABqO6csCaQDTFGMKW0+VRI2dLaR
kmgYq7YyNAlLIMsu1hw4nlZOgAH76sZsH66M5/nKeAEFt2W2G+VHk4igLYEd
/awxPWvDe83ZS4nGj2LxfngDZtsO/MTL69WB+IaygdMYY6rd/c/1mFk2pXjK
s6e4jI02q/iAz1VB5wAFQRkScbmlH/39ma66ZuP1LhkGW53y/M86ZMOu/8H2
8ZQbaXpk8jsXV3Awq8J2zKQ0dwk8c15xuOvMAJGgwS/av9gQYJvo3CVeQEs5
gYMCm+lUz4NpyKDjl3ygKqP0wf0OzhFiw03lzJKCknlLS9EMip3ihYIAL27w
j6EdguUzTOv965rGF/1TZn2qwLmXXOO1oOSECVfGDtNnIb/vl3gENQ1df/Mo
d+USXDuA/fq9kyJtrBZmd2CRpg6m98m55GY7cb9TBUiXuXikDmSk86I5+wcc
4njvOteX548i3btiFE8ANXyf7oW49/0mHerrApqeuHXYlt1NkyXY7AhiP6eJ
6A0mgH/NRTWOKC9x+qYYq/+xhYhxr7elEnaChXysu4q/V+Un5u8C1tVMGwUp
oJfuJNS5aeXjZp/nKHWNAgPDOl2RrDbtUbL9uc0GAOHj+Lnp+SsbVo0ZxL6J
yXl9l1HOE2bikAl1XI/SMnWyG/EjgBl7QvdplFLRnCO78bAZptcdnnOxIz25
2uaTtR4L8TAUBJmNwVUn1l2scuce0m09Ywvb6ZpzUNvZ4EOLa8XDIogoLtXH
3LVZ9mvKuqL0bJQxQOtbikLscBoeHCp5DcRmM9+DJUe7gHhK3BfVJNKfLOig
TkYcCa/tuYkWiSP3RzJVxA3I5hwbROyLjuCKsq5yc2kfYbCF0sBq/+kWxUrl
z1rsTrp3thKKBBLvdS5OV7iOfAWyvdyy2KQh28+0z9JNSEcgxpDilY46Fg7T
7yqZx8LLNfcDkd0+Hhr5nZARoA2MiKpOc4+/UBnOEaNqi+T7rZZ9yJLXpqVh
Pdp0nbZINuXWxNgrL2AyZXqeTGDuR1PIMx0VkZPcbPsGyK5VBUsXBFYFz+GU
6KeRPxv1NMyxcgokXqO0c4fIKHcqGEdJ3bH5K1k9bRB9XMyhyxhBPgCoJQz+
i+JEkn+HvP2/0W0lSAT+bCsS+ur6B/L26tj/UQgyO0RSrMF8iPttWC3a9T98
BEZH7ptKWnhbuT241S5iUaGwNMr888gwxPp/kt+uaWYFLMzCqqEVsukDVuTW
H3A75RnERPx+Kb9k8d6E17gj3HmgBvPXa4AYoFCnD/X2wdK4P1ny/4M2/QtE
Gq2yYrXDJ8T49pMxWopCctYp7BkZMVB7xJA+YAmwKHjjd3cRAK/gFhcyq7d3
hnvbghzgJNVcyhavyoTBWxjgL3Xuy94rEYHtvoWB7OkRglv+evraQH6lCmMZ
lpLyrepWdHmAN7V/PrY0412sceIVihhSy3la/MMH0auyVBhD7LErwK+/ygh0
aL8N1FPh4cIy9dAtDXg+5+Y3Y1gB6Y59YSfpojoo2sfDoX+HCm9Y1AeugG+2
UlndgULVHbFQ2lyYshXID7PEKfRsYEmojD32D6ZnzPhfLDGuFWl6T81CLmLT
O3xYwhbSXVFXXHiKoQLcLsdKg6eJ5YBTbK3PqD2g92IaEVVYOk2uoTlyiKqo
nYIQ8KTlQLFWji/i8pD5TMioreX+J4TzEv8qJJYLd+GNVoc6w96pRSaBq8ml
4sZEYOFnpA8WnTcQUIDBL41nXGqX7KaipbjbJUaQaD+xl8tapT8HzyaSTnAw
IVubzytNk2EpbDwl/nLMMU6HoQv+0WyEAzUUysxeKimumIUoiBSwF+Ya+71T
4OtZJQZl7zs7u9NWwf0TJUbrkyWRRdc0zTDEqf1IkgENshSB7ecRrufIBrFd
yfiKhrbw/IEX3z2jQbJ4p0P8dinpRQTzP6uDiN86b0lLYaKh+j/N8Nbvdzg1
hGDfPs1mH2ShV9w9O675sDdjtQQjF7CQnMLEP3f1pxCWi9bTzIC+xUORDVba
F7/ig7Bjd7ciS8sWIRPKMO/9/wY8HYFLAHq14sh9VXZIBNyv6lXsdlxHONIi
HI0iPmj/EQ9AobP2NFaQImTuuwXsOhMfgFSM9Va8tWZscbYf458tvSSJZMfL
SU/eeRVI1VHBmT+QpcpWssqj7GJWK6OHhRITOxtuFe1ZFkuh5KIyw+Du8Y7a
NkwGB1bQRQyQRvfFx97jM8Vj76rykh+K+wE16wrL/7bznfjfqHJUMZf//w+S
Iq/bqFfTvARROsVgjWcbN5gzrSvkPUH+iAvW02gIwVA1varh7JKvlGTYuOM0
Cyt6SNqDZ8wLGTMubFAPkXlt2XzSvg+Q1cLO63l0LY8evx/KpWpH8mbvHDOQ
B9+HV50E7x892uq+5IZtkPVfBr+hXHo7Bh4kfH9RnolIT1KYxDH+XB2XQr4c
Oq+xX3gsk5OHhH+VXhqvWS9n6UHd59aUhvZDmDCktslvxa5vcAZug6iWbK2L
dMYsgR8NbsOWp8oevZ7CYh6OkpH+EgBlwBPvbSrYZMwz8M06YBROH9g+7qdL
zfBCTK42YeezizME9OTizXU3jB2pjsYfROyhYysqbxJNK8UD4UW+/x29X1DJ
AWzCGBfj02KwSaNQ3rrQQ8mah1t1UXDK9Zds+lCSkXM1KlCjbw81I0PA4UfW
uPd2oYk/1VtEmSqL3pHG/IpcpteNwF0NDUisOzlN3StIjEY6FwHf+BzB6HwP
2SHhBjXfXB8qRpZm7f3bA1By44WHSM9ypTi+Yg1m9CjNJ5wXdDCf1a3GAgrl
iSOFaYQynlu+cRP8115RrVSQH2XHCQRzUacQdSdTZLUaDeus4hi5Rx6+T77W
P2/yiXStjCB9cYsT96irBXKG1OPLXain/1Pj2GUjf/8zbjVT4c4g/nlBXt6g
/1cP9K+vtaVRGhZsU0aQlObAlfYBgtqdwfqAYrfIEwYrpDqaLMw8SsVfxRrT
6O6X1CAj+cT9QmTglOspl34QtPt1m72/mLjKq6yC0ktMMx9y5rxtoi/H/Aem
Spst2LRZn9hpZPWnOYW7zvByBPqX5EkRHAxESkbU9HF0QElyUvsS5gAJEjyY
CkW1Cn5U7Nj0WWU84xt1l7Hh7XNEVCx1NgMaXW/nlZv6S65cRYyR4pq+5qKo
E2JCzJlT9hnv4+HFIJszvSqcDnGDWInX1zupaJbe6xoNpVJxpyT/tCqnwGhu
BNOdw7rQBnyJ4oGTttLnMGym9Uab5w35twbgriXp7Btes5wLXNxoMiuDEElX
x5My6qL8tAWhoGi4XHzXb3NlTFrY/GYsxiSHt+2Zs0ika2zBYmF81DW4Vyym
/5y9qlKzT8YDeuR74FOZF0uTJRwZ7UAT8HpeY096AuWccyWj+WJCvvmLWwGw
5ZNCL5wswGF1Lf9wqXVEyYekrCTMqOTiJ7MTLBEh7Dlg/yUn6jy1d0XtNIqf
1fN4uCNPwT5Dz4Iok1dryUGeKatl4ScNJH0Pv1cFdaiwTJZuao82TPrckiBW
B5sMZTKGVrI9miyaVFN1d/bWx7InV/xRh2NjIUkWwfjpZ17yqF0tsl99iiLU
WvbYUotAhJMDsb26y2iVyUqObpi8RkmdvOqRgB/zlvUj2uiSPKRRbDI3mE8b
ENkb327/4R9FM8YpwodyGZZxHDqodV+guRiCVLVdLeJcCw6tJfrRi1lxjNFh
LtB+9PxbPD01x9loAe0bk8VTr6mKhnRqqzmS/DQRt97n9OpTVHhIttUGRSFs
E7UVeSDkk32Fg2TflXPk+gxa7tP4Cp+nmrWlLsj8iCaXBMxJQaxRbPxHcUX7
Wd+4rqUYb0qfWShaKKr8GoT8nRXTeNKYqPoj1oqSrROdSBZRCIaXzzxcHhsg
SLMOedkvNCnp3XKDAQsVSR7W6sdrFTRSHz3HQjj67kHP3W1VMVqMcCV775FN
2ztgYMsPiZUDmzoG3AeEQI89vXsv6n6k6pF254Mipz+VLlcDbbVXKrNNd+Ee
2f52MLgAPe+zbIWJRDSnpN+osOZ73l3eZ4QPCjYwW4Mdklpk+2sF/wFwozzv
K/MC6psOpj66KvWfMdAO2PWJfzEl5qrmB1TMbY35dme5gqsG2Ss6LMayfOMh
4bx6gRrTke1KFWZip307RHKd3eHIWAwUVrZ81tBcstBd2DFnbzNitozEsDUX
6I031EB3R5b83z/8Sk4zgB7TtQ7B6PsBbNw2q6/NOY3hqk449GDNFFGWlj4B
4t93Pzqc4P01sXiTyIclYYNrjVtO6zcKVLUGl7znu0FC4YMJV6RDWxc8hcUs
cr5NLVFp5WVXcBnUhmla48h6M89FHa0g9fKdmitpWKc8aolzwPbtPv8t3HzD
rJMZdfpBLzqAk/aoMO17LP/ABS37qKSZPgxmBHW7rVaVV2vceePsvNwAjEdT
mGi/hj1+pUpoGHmY1lmw09ekZ1TOpU1kfvstpDGzmlb9BQeq/1snVZTGLMQW
BAq3da5R4wPHaAJEqsayRlEnOdCm6uZAMz4VCcPj9/81W0EviNoR93la/rUE
P6iJtZRqnFMW0EOx0kpnwiWNxrtuNcdIjeDGvsd3x3taSoLjemjnuGxprCbr
js79rGjSlkA4MyswxN1AEA5D7az8NsrD83O2pYQVr8LrDwgJtRls3gk05c/i
8fTON4efjt6HYrK3QfHaZK/R7jtf4nEAPKFwalg1c1TOj5rLEgR+I9UAO3jZ
I4Hqke1Whh11zZNGn0SEQxeuDecrBQmSTkpT8pD+wPpV1fWn43h8ahw4XjCU
UnzKRe8amGno25/yqzWjPHR5rW+Onk3i715tO/c0Pc0WLl7uh3wL/fxtIOcH
1Aqb6db7rQkTFA9psgDYpArHf4S4XGJ8oXVUzqRnwLnLuGk4mUCFwd9WRDbe
5k7rzxizY6jgVh+xvbHdoZIf29OPJymOMseV1OMiWaUhVozSCF2r4qp/SoXN
38069YmYOYMdGOH9XoMqZWGgWgpOv93ltN5U7uhC+dlIA7b5EaA7XwXqGv2p
4EJWWw/zTmXGK4AY3v1p106vVGi5AKx1SXWMBWuXDt5NAhBMapA6djpjOPDz
YSFcqFM6BA0bV2UIzxqri1B2n+PfcdL3Z7b7YYUXEokPX0wu4VKfFDA6N9zB
CuLamOw8WIUB6w0yhQNvl6X9mvQK8/tY+EUd4rmTmEcGcG9N4bCx/rYVQh75
xjJJlfJVfFP1sJPvTHDVc8sRcYKpYgP+B64eWmE0EFZom2oNcTcFB4p1tzdY
uWk30A27pKodpgUUiNjzb3XIg1x9AGWhvHH6BU6O2i3bkh3X9Y8wzsvVTUkn
UfBU9jocL2FdtH/GeFaueNZVgDLseaYyS0PDx+KbVFPIzRRFoR8DzdsmHEye
BW4q9FWsI2vFGKuYQTJiLxBZypHLfj+CGOjm8uglfwqgieUtMbsApJcILBcf
qONu9PB/2w4brnAD2qMJlHQJx0sDW3V6tlBZQxoYzGlrB77yM/mzAqIjkYS3
qTFQp59POzbD0ogQUr1xYIIgjqsSIXy1qJpuGJA6hq8KaNKdB45oUU/GWVNC
zdRAlMUZrwX5q0HSjOCCcS1zmIGGgalUZYlBM1M1fjwJ5GYWxn9p4B5iRYWD
e6bVgoAj40uhToohAw9aQmf+i28jcezOPpX5ui10MbWNYTa7sZej/g6JrzpK
bG52K3IWkAY8X4/xwwL20s2z/SUsre9JoH1FHnI1uv06vTPMA0s6bqIr8Kki
TS4a/Sqe9hKfAVlHKSTCExh/jJTp0HucZ6HB36W/AxgATIwHWM3T0NKDmFDG
Sk+y8vJ3fs8j5jlX3ybpWd3t2vobLj4XqpC2ugfAmNxbqY1K5APDzMIAxjIm
d2IcD5x0VftYf2zuht9Zj9wbwI62ZfvA6DQND6B/Nm+10za13icnMf27B9gH
o8Rn2KuQEwvAwRpE31zIfkG3JqaD3rImJgKtYPi90jWFSXhQVoV81kFd1p4R
HMqtmBAhGZvFaQkurR4GK7idM8onzQlSXSK1Ne+pkmwvT25cqVrqYzhfbnYU
MW7VbzHypS67u6x2VwtYAOQ3f27J+kd9yMi1/5WlcvEeEKZvHou12FYm+CnB
9RxnpUYBhvgp7atr2FYn8bbIPDAI7EH6uJN7nNJtCH0O3DExJPpOwDoeyAsa
odOP14h6kjLTmNKRRTCyfYMv2PC0F5blQvosCGOUZC/TqyJzxFKZjC0HZja3
Bx2bWE0S3UFk7q7/rrfRC/MiZSHHB458mWmNpfq2JziVJCvobBcz13P7+OMA
DlAmWOTeXZ8MtpujWdpgjGSgha5JmvXDMl/4F+Js5pzUrZ4Q/xDXUbySbU08
DeY08mHDbW+t5vkf38O5wUd57sSP+beP/MuYh5aiZwAkEjVHHgdr6TNq1INY
9xo3XeDRUrRuiK0xaO/vc1eboWOjPtrJSKDCt1vwQQR6g0MVraLxDeOxbp8y
Qb65RgQTxOtFsnKwgHWcH6yz9epjUjczII+XAwDbYQO2hj0lwYC4C7mGjNWK
EaAtY6cy6CSIoEeei4Oz497JFNWo/QDeROwCEqWmfSwQ5GcUA1Zv5KCBc+VT
PNYi7+wO7vRpbRfn+SJLBVNAnTdScmtOwkzSmLDmoZqe0tl6k1P0jT8wv0UA
4jrECyQrmUyxtoU+A95ISM6oRAbFCduXJyhJUGUnuC3AOePj65SB61DtGkgu
AuRF6eQNeS/SVRk8wM2ghdn8yWfORgQIbchjscwwcGmqKUfwFoVCAiVLrgO1
Fhnf+orwt0q3v5PYNhjqFr3bNgcDV2aGj0NEo9Sh/jsnt/51YlEOgbnw3Qhy
dYTIN78ZVQXhImunn/Y5hJRfNTVQ20dg28uif/XhEAGHRj8d/n31VEtvemW8
gx+fnOajyp33cH2fwz3wnwIixgaQV0sk/oUut9FQixwyXDlmYYpcNeLMs58r
NB+ohKfhAyagHaYw7UzrMjKBH/WMiZvcJO3+gzE+9Y0mMMW5fx605AeIm2qv
4G+mqxOPJ0KuLtpXwgbMUi2R5Eypwiz9y0PQv4MQjP5G8z2kl5q4eWuNZDB0
m4UbrTLsZHPp2lptmsGG4+u3enIAftyRWdRx0CzJOVuszC2SvJN21EkH1uUh
egmf/zPOwndluWRuivkceWdrM1yORn3JZ5VfHyFwOJhsUVrOy/RF4Km3a8Hd
NUG27gZZHbojWD3cZPTqDUjXhzeJ514d6JG9vn4V0v5X3jgQSWAM7ohRQBv8
QonSaSgMMkUJEKCHhL8bn8QR7ldhZITFVLxJqi08WgPrC2xs1K04pH6onOsJ
WTo6O7gCfn8SUETnrf9+/TyOb9qiFBIC8IU/IygQF9STngC+TwyDz7grNkqI
N5wb+j2+hisA+yx709pbqBBzAgpsDNT/08mgII6zd9pJF/c5w2pSbiupv08y
vsLPhYXO6BVEw7MspikV0RdXA8zhvfasx1tuo62A3GM2WtQiF7e6N49MPR9b
RGqqtoPuz0nQmnvGyajuSIceNVt78ZPpgNMp1Tc3MeLz+78bMy5kMUKT//Ks
42VL2KTEwFze/W3CUZQcKnEPRqSeZhitGAtf4o6gra068Ed1nCP0PB2w6Kof
dhJQFcUo77ZpDIzcWGNjaiA9BknfSYk2uahPu+obfmecHPmt43uVb/MCvTTN
TS3PaXWrBQrKR1sQnxMnCxT1PqASl1iTJ4NYMl7yOgtMr5YMg36X3PKIYy60
/cFU2BNo1OwJtltoPeYt/9YtjJjyEONWTkfhQPAcHjh2TPCdRvy+TXpAPEAU
u3uW0FAn0KFnXOqhISK9DcCuY/A5NJhYZQAKTTOaITh0G0AP67k6rNeJG9Lv
cABLV/Ho3aiRUxCUIwI/ka2CTdSW5XKApsY/+LVzcZsYEDRmX9bb3oyh+q51
706pd7aP8MbeKDeJPpEYE/lCICR2U3bj2Qomc3IzoAjrYgjFUyhrmKFpJmJG
+IdV4uP2Tc3BiPlgtTdEA3P/BTeF+6mGJSIAdETGn+smh3+y4eLDUbNX/ia+
VvGawC6c5R3nUo2kTVbuLS8cSfZeDJEmzqg+NpDpYDKrN+Ezdula4GB9vXsh
fohEYb5/L4p/Bzpt7m7oMzaC3qrSeJCc/YQ7WD6fdHvvDFB1RadUHvbqv+N2
LpyGVTRD9cHZ/Gv/7Ee7S6c67EtySe/Ulr5TXckKcF1S+IEyRrzZB8yWLdG7
RbxJ8K8aWMXii49ugmy3M94X0gRxXba/4At3sPOOo8BVmkYy60sGS4NqKGv/
/ZalemXfvG90nRP/i8TR1OtdOXRKtCtjmYQUiXM0CvFxBqcJ+iUF5BdOePPm
mRnvDSsNzrjAaWlfPF7PNkl13BMFJpJR6I08WOCwJpLSuxw4Mbu1Xm3c5Jzo
W/6e4vzVfnLPhtyrH5PSplYPxMjUqFdH4Z+bwmbT7Uc/U8QWcrJs3WARM8Ha
E78koOWeT47dmuAsISASjO08rtU+snpqJk5UAl83x7SpbOXJTZA3TZ6ZH2RU
Of0ze0YqHOeja/Xi7w+NVri3bzoO3cA4LD6TXxmSlt+y2Hv/65sGErAW5Zu0
+sL5ncfqxAHzHsozfTLSgMlhj2nWz6cOVYhlVTXmvpglsjmKwMFjjO1FjQ8p
c8LRJhcq0bhd96ZSv8kSKshv4ekhE75L4Pc3vNHzImSpIKQiGpSJZUBv5e3N
8oMep+m4ZWQZSBzJx3T1nvWRjESMC4kwKXWQ1uB1cxkw2E5z0UtcYwHPbdmq
i9/iMB5wPYPqsMhsaKSB2FBnCs1ttxkZ4IuZfcqGSlb+4Olf+AtCr5Sn1hgv
QplQ0VoJigPfGU615Yi+G1p735ay78WzSDZNkWk8hcV5pnxfTR4yhz7hkcAp
cKFDDnZ69mASiUxO5k9JWizjgvSb4rv126zbEb3+NsXpx1uHiXL8eEgJriqC
A0XZOQg1no6k4Ozc/5MqoJUfPjIW+eHYKJmU9RF02/SmJrXPTQLj24vqASOc
8mcWhGFsC8IbHX2XIbO2+QE8gFnCIL/aQcD2dNRumcOIIAosiYzUgvxl48gn
o+1seROmeutqXAmYmNwzPIPX65IaoYgYoUaaNe+kt/AyotSfWi+qTJpvZEvu
dkWs+Wli5vgfBruCzXt0Za0jJ1qaSkBLnH4vtAg/M4kmjG+VVQyiYJ+OxWKK
lKd8+FkO7vV8TkuL9GCUKow8P+cE5lcd5vXGyRhyyf8TBUEQz/NhQsa+O1Wb
S4VK05q24LisqDhbEMFwaIaZ54FBNjsfgTLgNf4qgqWjCU7nBdlcJIPm2bfQ
pwf/J7FrkXLDkH7iA9iqT59QmrTyQ0Z3qdRmml3kBzoruhmY5wHXJhTwMhGn
tltD52HJ5NSlNPsgfDaH3jF+8MN+dPYmnG71Ai3F9iXOh62ZOsx76HOI5Xvi
NHAdcyXujmwMGJuaPCI/DxNxlR+BhWpkdqY2GXgMFtPUNDFOOdPkEXNg4UUV
H++Wqkzx5LXpajH6vJ/dTL91NAEbZlKZx/qk6ZUMiWYvIXoybqOFCZDdKuGe
Kofkq+1Wgfun4e39brhzKgjbzkb3aOmNav8R9jLftieoqOwOMScrnQbDfSRD
5BRD44qxGpjm5uoYr4Hio26ETynnAkosaci2jNO0gaSdO6ck3VSZi64H3g0l
dQyIx09mVEgOqAy+E4D0IcE1YnKkUF5sMpkV8ts+MTJv3BoUw25Uk2B92Rpq
d12ViebSlO3xNEfsD7tccFzT75sKUx2QlpKLcNfrEZ/ktQi72mDLpodhrNxQ
IDgP+cuSb5Z61ZMdahVj5r6U9Gfr0GgZh5nAn0CaMAZJr1tU7Ygiv9u9MqOj
rSCh+sZ4J830OrPbWwOpLZZjnQQ9IHzq/FArGEIOIAF2F7iZ0XtIDa4CDEls
ZnYRJSj5hACZS5wllBLHbBS467VQZMLktcNkdsg1T/XqHZiXnEoObgOi368l
ZayntxrsiNw58gMJM98EznnpgeYwpOQSyrJJ5uILSE4TwyEBZvpUVCQ4pb6l
rZ13eZ/JnUtT7I0kFnOYzwijcYbn/lVBLWxCPU3i3PhHKthMCRoT8nR7N5zD
HBrO1L46RJLaU6WRLlTSymHWCYCxodGnT6h3vfLNRLGhC8Q9fEsFKmkQRPtP
s/5ud6boD2918T0XeQB41GWX+j+8jFiphh+caZKOwfR8iEjnFAErwUa41dJW
tn8zYc8dz4UKle1T7bhqNY+TtpHjDWr9zEYqfH1qCJWPN+tIY3O0uYjBqN9B
x2XxO4xAaWhsAY2T2j/T2qhoJxjt61o6sS6YHwkm5lIJ8B535ikE/rCG6wXd
T16lLpJo/5U3LpFMqZzxEDG5s3R8s21DZYjgxHnQZ/Vzxq0kOIyM/Qit7R2Q
M+CAzDkp9THQNEn/cq2EvJbm9nFWg6rno93cTL53JGlu3VwivMQlYgfKQwz+
elTtvyWqKFf11xd1Fb9LMx+Rx4OfRwbCp+7zKrQykRU4JvHzxT6PMCh2Jbor
C8PWN1JhelmFNTaeZJ/B8i3csuTFIaN3Ow76EaD+ZjqV5YxT+q5rPLtsdAGQ
WpY4S0Ys422HkkC/L534OD5AEqEtniM7oWvQRJR7uomEw+04p7c1pABrO2Im
ctnj+1QHAQqZyRrPf120MediBzwSVS6hZB9HHFlW45OY8kd4KtAKM4uAQGoS
Tz9ZhQiJPfgjCyTe9Dfs9Id9YPcRsR+IPm8d19O/H3kp9ezYjBhWQ0yGVHSa
7jBsaWMeQyvf/4PROqmwkWndwekCYWIitNsHFoq0P7+mA5rIgQr/Sdw7wEw5
xAmMdtMAXLYiWyNtaopU8oPYaNXpLh6BOwenrUJsPdT4xskfEpJJ78+za9cI
3cGbmzmTWgXXlrGsx2hkl5xtt7R1O8IsGo8HpfZKAKSK9EWblaz4uiPzb7of
qXVA8pvRZyj1vMSKstde0NzDCN6wE08q2J3BD5CroyrnSS9LsXIqoiRAn84T
nVuXOl7wJiuks8EAdMwDOr0aA1tPNYY9Yy6CymezRysxhVVv99AyfkFpvLYi
wqde9+bTBgF/nj+jH4dCxHPTSLh4HD70N0gVnIJuAI3KtpsYUbmDmdu5b0l8
wXmYLiRx0w58FFq5TJJMSFVABprmUPlBm0Fr3FAgWCwNijTsFcnxkeCkn9zM
BQTqN3s2/LJmID2N/Tq8gm5LS7FTjedkSZHO5OW2zw5JVRaA98vipPCvk1mX
2+7txXFDY8YpUwi653ZUlpInr5GCaA9EL793tmR/IWc9TPhqBvNVbcmdFpko
Q6r/buwJEyZ3OtJ8qgQTfY68dDZOuYboVEWN9mlccN4wcP9kku3UZ2+juVaH
ADExHcUChHa+h0lc8dsm4x71Gh2nl5DUf/vM1LVbfdkpoN8nXtDIEAszTAtC
nL+9mF4ie5Rhing9jXhmjnIMu94AHHAOl9g5xDJtKq7BM2S938FT8DAxhjId
PkYDmRVxwI88Fjdg9XukqLUeeRt2I8KH6tFHj9xQGy4jIJBRyVkKZYOB9Ydp
x1IQ5fBMRyVbKr6dI9RGHmTYDr7s7/o2m04YSiZM5og9ysUXaeVpU4Yb5A+3
YKqjInRu1bCtC7OLwycrUlnK14/vjXpUsb/1F1qT0+LJlNm5ALmjdd2mAjXk
E0Y9hP8h+v2PlV3DEtrsv87lACTtBFJDcyf39M9qB3W+co+pgmB5pV/huMw0
ttG/1NR3Rp4MT/vFvXAzp0yTIQYwJsYiXuTF/kMhySTS6+l9rRPOh7DWLaIX
NP44v7kvLAoHT23L1reMq8K7pXH97SrJSFsLF5fS+nhWNOpfKGSVENud5stW
G5fwdb9wduhZqIKvu0Z+7gSYaz4+BrKXEe1bcPCt6bUttrHLinS2iluBG4QC
+Bp6gVAp/pTU5fM93ETtMmZB//EsYf3TI763D2/LCJGzk0EqynkswUZXjPdT
2Eut+5xj7kba+7xR3Lan0gBPqDwL+hGgtwG4cXpQZ9MhzuztS2vHiNOiZqYB
WU4pfGYkzOo6Pzjdc/ah/dMaqHQznU4w3G5dYhfpTgJ3bbnDJwOpEnRnTKFM
C/eYe0pyrvHIfFTHfz1A6B899kn9omIVe8OKzPhc8yvZmqRcaAZIr5nTo0qv
pAvKq2J3XcZCFx26BZUmWOw0rmqnj8nwxvVnKAqgfrG2s5EcFnzvPOx2oXwb
i1FhpYddi9HB0WnfnDXgSc31M2jBiRUMO35lKBHMI4WjD/Iy1cSy4DM4qh8Y
VZyklFOOiOpxfLdof1vlfWtj0YoYpWo7gml7bOoOggU5vvjgBxf9HXHGRT9L
x4sjE9GLdjLd55TDV6iEwPixHM2lJ9/Lfut3zD26qYgtIClAyWTEYc93K5Da
jQUv/DOZ6MHdm0nuK7OtPVp83Z6CtROjqVWsYn2wnf1O3ig0P9xmizJEXciK
eGt5q9nHxG2U908c9f0EdDUGnWjpnH/L21AzD+5ZHAJMSnvnRQW2T4cTcA0E
CePLOj7GZkfYef5G7DpIs9aITLkouJKR9l6NRsTG5osuTc8DedwOoNskEXSq
GeDMb/0EwV7McG5xAhqTydwpfSUQIqHB/uvlFQfWbU3WrpjviojlpV16iR5Z
nakZjYHh7OYPugFzbFBo2fnwBnzX0Z6lT6tYOEffy1S0AP2oxHd1auPyINQU
FfdqaIoQj07Cr+dLrO5Qu+BN93u6T9etkMQm/5+nfLrXdntrsrgbUCv4q4Ar
6jtMoypCAv1W8aBH9OFyTeZoAGunYZZoUugwJPjJHhtyPw7+XHlD5Jn2299L
7lBgoTzHBIky3mf4FFd3BAFLCsRnpW7pqtNRlazHyUVfh7C8iEgRVkVrcfBa
v+crXrYU8+RCNqGx7AbdTX97UClfTxsm1Q8go+aXydLGkfA0NRcqhUJBJLJW
kEwOpamMfyamczKiZ1vwS4PPJiiRvGV9pEGZByVSGxGjxALRN8SYJdGOF/Nn
a4dYfYE3KSRD7VJm+dYL2l98qYXRDf1VRm1avfiePT1jrtnIie3+WYpwjnDZ
oFL8yp1G9OofkVuoWNOBpNodv4e1G+eR9HsDY5+xKnBegMG/CH3JeiFu5ksK
hCGXBe9ilISSfTVRi76zPtXEmxJF0RjdsNrZ5xvU4pQohSTMgvGpInfmY70j
/JGCAHR3/18cPYDRcVp3aF2VH1bihG1iXSuIsjuxDX4YMljhj5nvWfmxwQT8
HoLIwpzo3jcsns61qfPLswglYT2nXhiMCqQSCMBBZKT2AqmhJ5Cro6OySPdz
hxC7eyttpx9fU5x++FGNqc39mLwYLPVqob+W+8LZmdBUZLgSrAT6fPh1YvS1
ZMotlXAMuyfkBUiY6khSt8PtvdU4E9/EZXpmKJdGKSk6vnXl6tKGxP7bnLD7
p85C++m0833l5vYRp5DP1+a+22vcmuBixA1x6y8evEEIDbZtVnNDdMERot1G
bTDcsKDj5yNIQnxMkFKSxRSTKh3T6rzF/r6HHzjorK+xmQt11LvSalB2Mkbh
w/Gfx44/M3DxVk3Gs2LLYvdkPtO72a56Ol7VJUli3t5V9inCgqJmauvzJRyz
FQ2PL1ExbbAl0zFJ6pPmvNj1MHHxmUxX+nwfMeiq7watfT5vk2ePvhpiIzCq
qwVGXGmgVgPPCNxlfh/hGA+Vqt2kDRiWJr+72MwjjU4NvGC325put1iJea7b
2Wt8J4ftK4TLuSWWFCSOTfEdXoRLFES31e47l/dpfebvc9IxcmIWPL8dRfqq
PP/sAtT7yDZlBcFuD0D95FMrT2Dc3EebJdlfEIzQV8Sz2nL+a56521IqIGrz
jJFhIR2TZGf04DXce935SwpsZ5xUwPoZS3L1RhSUhQXnQlT7lLWSy0akeKOj
8Tj1IAg5wl7drm0Oy6ArHhXxmiplMb7n2fWrjDkL5eksWXMA0cBi5htTnwhi
uULU+Yffa/cnsqqQI422zbMeIxwGyY7Gh/7z2l7Gny0PGWxgAmG1DJPoJ4ps
wbyqxJrhARKz0vseLyRBKuxxIpImb1F6aUvpNtPJVIwTh8C9PNRAAFnOApbT
Rqm4gm2G9rSB5DofKx4RXZxbMN0WgZdX0II1KDwYLZqJ8KVPgEFTwZBTCr53
mVZDwdso3u+L4NTufjGskCULo2o6oG3uszogk3+lav284tWGU+G9cTJp4HC9
TPvE2V29f1OUGe1HON7nvM8la9eRjmLdJLkWvLQA4ntmTv0XKqVbVw/HxgNT
yQJLRabarwO0mJTKbfJaHKqdlTo9zMW2RC9PztHKlzo4A9jLdq5lJu4/GjwS
/ZJqlanU9Tda85ANEDx83J5R+tuEzqsNnRCAKPYl51EQvFmlMfh6KJswts3e
mqCvZkIQALD/qc2HKUlpb7uUQ1acOnZ9J/RpM7V+on4saa3LLwbmEZ7R5UUe
0tHfAp+xeKdGuWFI5gUTdb5Z2Mts1jmyfZ7MYtP0Zs6TAl9lvDoL5xIr6FXx
3JLV3Fm3xLIHpC/AmV24QAkWC/DX03WbVvNiO/zXEvZvHfKTm2EKU/hUBVOX
8Sz1HpXpcKPVCrTNa3AyKmZTmWMCBkhgP6/6oqsGo6Vs/Idi66KYteIcDzis
lKfj3IqrOEy0nLGz31OEb9TjsCvz+dstPzt5NQa/BS1gL3f8EL570KVHlJ8o
Pf86g96ZKoIDEFnHoEBWQ8h9hhvql2D095hGlNpHBKxEcxUca3nOzjaJEH7j
KsPo14on4qn48uMbHNzw/HGnJZ9Ze6FPNMJ+snLXq4xBdVoBjTW5n1rLmDv0
eNoUMgHO+uLJpkwu2H6kPYsaHTZQfDFmRsFP7Dc0jnHgAZOybX6wRv25AXMd
qUShg8Almqis5E51qf+10FWqD0yF26jKePSFJrQnfUSSfym/erKNf8duMkAG
u5La0ozKnFFDhTBfG/wQxDSqZRqwsuzGQcCRDBY6RQtbNJ5Cuk9xih8I/0Ek
njFpBDB1kZMSIVHZfBQNwcIP0WF142brfTKEJrw9SaG7LAL3vuMS3bbjQLoW
su5gRKGBawl+KRlzPWRftf6AKeV0Q4z3BJi8WQmji9HMp9LHpFKtXEh5ov21
W9T27ApwsL8W1FK7NN1yuVU5POjSrx9Lc0P3jflPhIQtAIb2O0swht7IuUFy
SD3dlohtZ3q85vSWK/jC8wrsEB+e8pFIS2z19SMeQkq1DHmKi7zJLvHLUkci
rZWTXzth/pssvgBf/CTS2jUhKSQLjV6UuAfEHVHLDMG08QBbqsJcWbunPLXj
3O7pZd9w63mknyIQZFKKlLHY51VfzUZutJo8Hc5ZQDGXb8yHsEZaGdl5UdeO
dZPXOc5y5npZRTjZZTCR7tA8gK8Gu4Uzoa36ckPO+1VYqF3Di4cuRvbk/ToY
tpyc9IvxSrDyJ3HoWRin4T4rjQ+IApbykNxFESEI7mUGE9Vg6FfKYcHNqX4L
vFSz/mjJ2gx21ehhuGgiEW33+FmAEynE+s91bdQQZEdQBb5WF7Na/cVkLG+k
Wc6tgBwp+PtXxjclr7Emcfe3sO0JBPnFy6kpTni1g17QSUj91qpTOtqNdN2t
CcrcC29aoB4GWnMjcq29HXTuatWKH7mQbThw69J5XP7es2tHGqGQmBFaxe29
uGXGmz3XITTbp+/jeX71g5nO7J6vxyQJwpV5+kKPL1RmGLvKCzu53J0jIPry
2Wye6KtlJ4I5wHcJdmgWj8XaFIK2xm95a6HqiFXpJcqYf1AywbQupmbsbiLP
+9g+6gqGH/1bgV4y1QhpFAmHZItgsYn1mrNj70Yt1gKQIVM1pisP3pQybnDK
VKnMoaNAl6HDsL3ZBGyxxT3Hq875n14deqCfbY4KLMAXSUldKYnFhslukXTI
JrtFkYNhjynLgr4iZYAaLKNLEjRNjv/L8FG27kTNfKy0iEMA4Hr0y6N495A0
vADdt7O77eJDWoC0by72Yj7TRUbsBbc2TR98x4GCpVcM0yoSCBALWki+NfZp
q+Tp+SyrJUk9ZiG5bEG89TMvT7+CRyhGacZiCWwR4CaCoUEp7CIEavCEqidi
3y3/AZDhCee0GAw9l4Zkb/ETeDlJ4SKInth4uAKZzPnx/vXaaphtz2+SWuq5
wWT1tW5qMZaam7BTGdpqgpRt58KDjWC2J/E4HlYZptumE7r6Fi1Z/9fVNWWO
m4Jp2neLwAWsTvzVebR4g9dsLetino9Idmzb88XqbM0258qVm1wIcywK9Gk5
X9RJc6u4lwAXPS7eEMmo2dxTbtX6NWOF/1Nqfk8IbETKQ8FSDEsU+u6gzzcS
Cm9BUTap9qdZqxgsKIWQgp7iJLbnDlVUN1bBuE3Srq8icUyDPH8GPVVe4ru5
ekqwYf0ckxgxsUrBCihjNvlE38FbmBmeNl2YqjN2XIkGPuJbdSCr7TB+rvEY
UW/2yasXFxP9OBAtcc80JBu1AN7n7iT1dbyNS635cvjfmiKXixS4PxFVTds+
jql+C4ZGAXurbW6evlVbXhMsY0JD3SJnVkJdh2T6k/TXp8uvL1KmCaQI6xxU
jf5Z/wsRhFApvp35cU+w5YuS/lpJ/Gxz17eQM0kZzWPmM5ICpoKGjc2oWWv5
5VCup1A6gr5pUh50Z1X4rwF6uy0uJCu7lfhI7Mhl2lAgZznJUH7GTTN004oO
MRWyKHT+0pm/5Z1ON45nn5fcsz5SmocowkqH/rnXa/zrncM81p5x1Nqo1gCv
B2k+dIcfezC+GDQnTmKEnx+S6gojr7HOS2R+HXl+rlyR5fdQ0OHrwEI60/fR
1aqOJwutJ28HmhpoSs5nUbxSSThJ7f24aJxbFmfPZNLjXAIXawMf9FiGKmYn
A2iRp7L/GHzTiPcJKEBHgrU4jmbKyo/83gZQD6VQ2MBEgnFqmw2tHj2ARJW1
GDwVw8NlPckdCvUJ+CPG7A8kCKAVSYSQus4Jn0k7I5+yueZZtJZDoG0Aky6z
0i5r92j6N5FJO00TbxxYyqKF2KOCGpo55MQwQjibBX0iWSiCW7MuH9utYwdc
MEOrUL2JYX7FGT4wbIf5W2Y906qYIw7ykex6Djx2zWTL+95zcCEKDzEnGh+7
SAAuStdgApvdXYHwqHto5lSUoRBFrcvljw74+cPXKrBJrr2pThPyxSJw+lhv
oTSqky8Ug/seLEUe6Q3JC6ic/t9BqMawIvAjiKGHwymENHk068BQV4GvDzOf
jEyPX+rsL5pZIbO+rlsiyMyD3ZS3cGGD84ndyguxpXvIrFUFBr9VIleg6ahq
4/cdHFKxj11DHCvedyOw676shK6XKLrCy8srvv8hXdsD66WRYrUJKd8vgdXx
im/0y0r2rAwYCTSWC+9W5YBgxP4eGdmCTyXcunQsiiqXDXPqYO+pjbdzLGut
3/glzkQpNngX1JUhkDkuDcpU+vzDlMLVsH3tbu2WS4e9HeZtd3I9ycD+oLNQ
P4nphFe6Pfb0Z4fvFbOHwRNSGhmt7OhHDEuVA2NFBCSJbvEIxtu/C7Z6n2nV
JsQCMlr6gmPQ6IL6IBSEVSK2WsDpzqrScuX7PbT+jQsP46tmsnNYz72VY5ls
fVkYkYYlBlCJcyuKcrGuAuS9X6rdbz0HkOFSyn1foLM9jYsM1ai5plvCyZ7/
F4xOavK5LR8f08mJNjW4JqfxzOsUO4IIxVGuAVjgHGWggjKtfhwOxZ6Ah1Ql
CatsDuQeTwyRtwGDhMAG40rocgU1NR0laF+neH3KQaFpjYaF72xnQC35Mp/8
NaMpz/zkWkKadI2jdNqmwWLRP28RgvDakCPJvGVc+R2QFj29booag0YhDy/H
zAC1lYlXsdRYqnp9EWbFwQelFrQ0KMV8tndWCHXYJ4aHZXXOwDWLDVoTTo1n
VZ3fgHlIe+LORCyKDYbSuuGhn8icjdzN6zgFzxmvOfK7k2dZSFlJbTaRIMei
jFaVHin/235MzkzGtjmDN+RQqQQfhbrN7wpOwp9XzMrA39KwUC/5ZG5F/3j6
6r+dxBAfnqTDteBtFQkYNMpBVim9tOm2UbSUlHLGdkkFBAKOYBGoECPkmoOS
KAUUcFbk9rK0y7iwduc2aIM7gNsmX044ekFWNAMW11zAD6HPzl+lMiFeTZs9
RADtiJlo/Ov3O2z/0SiMSHjkErv3xaQDDmSNANYpoHBOteObE6e0TwKtUVVO
lHfrJuZ1QBrze/c27d1n/96i8NXVsn51Hp94RdBgQ78cbQgiPXLkzTnLh/Wh
Q+Dcpmj7qt2KM5tZd3qfC8awI6pLZ9LDSbrtCuf7wGaZZEkBth7P+C1jkEpM
O2dYxY0sXy6dVB8UfuCBdfncKn2NhorYdhPr+lYOtkmAi7SkJZ7Oxt0kV5tO
hVlEIYfpnzPjgZsgOsynp9ODqBCA1PDO5OJoUV4tjLJZ6sR5vOhNzj22WCMG
YmwWDCMaYgCWo11MPHwcdb+iGamUxa8T+j4nYVySAuyeaYylCz9Ct1qnfqBf
rbdh3+SP1tZ1RRmQ+cOAc8atXCDlfmd1tJvTMLCAOldxU3itMSM4cUGbUjJt
Om8ZerMIMdG4aj5YHDX1HIzUvYGi36TO0V6qH4BnenIZpklAoypGpgYKl4oY
QxGXlaouxbUmwCCxoABFSz/P9TRZ++eNgqTXgG3S7gQ//ci3jNOI33jdXX/d
gx5c/avYT80WNMqX9ElJFPIywsuklbgGjW5QWVdc7szzVWaM4pmOGnmAXIyD
Lo8nl+ciJc9vSy7F1cpxJ5dkyt+VnYr5rNegIgDa/7tde0one2WoEDL9caWW
bMyTrt9OJH7LK9Nv476dMNlyuKVm3vonnR1enIo5AZfBYpZlaUfM26jXz8w/
0n9WsI6ApUQaLGaFC21V28zr28ESZFpSRiPO4blunXrsFFJ//YbWtIs20UFo
B77XDSwLURgdkAVuR3llJZDPss9SDREsVcQrhzlp6Mpre1EfoUk0Lt9a3UCx
l9cx0J2SYiVyWHlppN9N6bQAbhCVPiH0uhSqHIV0k2MGdaUrnir2Oi5GAvDB
px72gRtfyeiK8VlqUAgRIZh7eA2wx9atj7r/Fr7W/tpjsBPO/Px/+l9XiQ8t
JC/ECYyMVBICb4m/yos5j7G3iOANPy5mpTtPQAfoyRZ3x/hYdYj8YlaDZmoz
6uAvq8Ca1oLTWXUl9cnVuQrIFI1oEK05TXO9r5INbV3VDOWsljpl/0zOKeSF
EYBp6FIx/Wd+TYqbFes2eYc7bXT8KT7lRXxmDsEHO4RNhQUfrzhJ0xd4+dyf
wOgqpCSwa3gO4AcUpiCLIMXoDeHFuq9+hAsKOnptqltzUA4Zt/3YSIEPpN7S
kLSUnDsE16SKK+M7E9P13/OXJsEFoWox62Zy33/Z56lNRRpX0brNxkG9CXTy
prxn85eTlFuIlwIGU1kxHHas1V+gf8gG7NvVnHjhWkN85X6DpRZCk0VRgJks
1qh3VdxOBBYLjsP9Zq36gan1ntdZ6OqfoSQmDa7fqBqlFno3nxsKvA+9EOrr
fttr6COaunZrx7I41mTHQQYB4fJ+bhuiO9gjwhIJyO4N+n0on5OosY3Jvb67
xAXm1TjMuZQ0xk4kebTurFp71cbBuQtW/a0oMCT11LAi5Ak9elasOd/XW6aP
acEVKJZ59CzBJzOtOGYFxjdKzVBhp+gfaPLXgMr9zqGpWAukMI5d4IfWyXS3
SwE+jpaQjWwcQDLdlL9oSaJKMtl+siUyaxz1gpplvT1Kre92mAHYd1Kq6jca
RT8KGx3WwXKgTyrQq4hOFoUebRTeNLL5KH40kS7WbV2XoO6PAcydQ9x4NaFq
/PxW49YrP2bR6cbAxloLiHf6pCcc/1xWyVxXRdbMvdzt2+LTkGB5UT+rQz7d
xwMKeSkTcDG10UTKXBvDlevhRgu80daAKkq39mVImRJ0J1wtXGxriB2AbMBD
HccAT7LkaYZnYuef8r+67koCdmmdhDyNkTipiwllhLm6kEA6HnpmnLkzh/1G
iKXV8xuI0zuTZMqzAxrzBI+8LoiEd8804AvWOmUa0zQoLKgHg/XO0oh/dvER
3K/FfG1ds3WaqjFQ9HfjpQxPY0NX5vVT/oEjK3wkp8csHu8SKDr5blVD7m7i
Zu7N3eLPMTUPPgXjH7TN0gT+bMawEiry+9d7wMRvtJhdZulMtYCjjcYIAu6t
vda4SxHSO/QFX+lQeAnagTBli6Lfkxpk6cCnMCe9QvW/wzXS9lJjCXlUN+8d
6571T1ZGMj6qlsrppNZX3CK74Uot0ZDntcV9Gu6j7RaQCIhECEqCi8q8On5r
r1O0W+DG0XBrliKTsExcaH4BT4rhbK+g24OKWDETgWmVJGmASde/CMfag+pR
tUjRAEB4f2OBonChmBJ0EmrkDnJDLgOkqBh3yc5ZD2R4KPaw2BoVMMeZFcnL
qDWgQGHmQ4n+iEzQF/X0hkUtLLw8sc0XLII0h39tnMN0uUqr6ZKLCtM47rSb
eRPQDT9WApaTzGnb6CIWGDj6WTDD1OyDuN4zjx7nWaccGqbMZs5HXMOmDe2A
7pVBcXpYvInrWtXuLqmoQrqKQlTs+4tg6pedmmS55qlD6gCl+ZDxQEeS17Q0
XDqy/alnHMakgecsN4S4mMIdqfrgUvkRYUOGGs2Rz8KyG/bYPBU1j7TTbgNU
DKmARg37IjQDKU13LjJLEWS/6+L4XHpbuoArudUvYEZ6wZPIyKxszgLVMN3k
yFQbjnjLE/wPrEvEH0XI9pwHQQvpyaYOjYXzbOnwlDvnUVg8/kDEvHuPlZcc
zeoQGm7QU4dK+/r7PgmomymhFfjqb6S8OJOVB6rXzZqOcKxLUkcniQHt6bgO
krl7s8YxeeLLJzwVf25Xi8Xn4FQaB+OkGSHDMENQvlzFP+ntciCY/AV5Iir/
uVy2M5RMuCyGIU08QNg6Vamep3WWALR7LVhy3yiXWsfEB5lnqLUqpENuUtIQ
r9bcGSgxgIoCX9us0kh93er3KqEDLdHBSqJzU601omXf2fQ6sjdwi0XHJ8yb
mTcRDn8IlAEXQGAanqjoUfozj5gF7M4BXVXFZYqysEfCrY6APqCMTGyWYCHE
2mqjeIw4hD+D2tzB/0Hml60FQzC5hdxQL3b3OImA9HfKDXzK+cULGrB8Oq+w
EK3gBxSup3MGGRqaZXGhbP79RRDEq8YYE2Kp3EVQjZ+2zTumbVPVxdY4eUQz
RINBbNF/kVJwCe2G/c3EPTqA8LylPW4e5YZUK67jhLQcpinHmq1YriGmhqRr
Ed3r/b4H7qdNpC01ZhyJcnu6Xw0zjnJcgRHECzXVN4D+E9N96uY52S2sFFrn
bIVzFkgDdayA7ChHiK3ReEvq+x7NPWtG4rTVZdvBuPVmh59ZPxQnxIIWKcHH
3z5gjGvUqn8AOeI4IbmX51vV29YJbDNY2vJLB3ObAFZH0ToJ5I9Z5MUY6fpZ
oyCsqJG2/15nT/1FPPrcPaX3q2IpCxaOfNsV9TWpEIfw5kLLvTYE5UuIduEn
TiiBOGpNrBQS0tZKke9e2DMDVKbA/Z6Jk8BcGElb2io22RzBLp+qFCUsh1dU
73u05gC0NnCx2fRcPYOX2hapBOMCRoHDGvlmaWz/jdRJaekUKu0gD2USqGtI
PpYUQj0W65hmqeXZv9/sIcE8qkcGFJ7CdECR5WH4VpGAEHy3wnZTQoA6TZME
6EfHGY30BcecKkHUeMILEY0YJZGbCAA1Ycal/SCNH7hW9GTiqSVvo1//O7FK
6UHxQANmX30a+vqUWEVrPXdsXVB7J2eYCswuz0ydPTC9QHLZEfSElHh1/TEI
jXq3k2odZbmOOrtBmAPqTOh2dVQqIU6+wAy19AvD8h2cN6nadFE/UhmuQ+D0
7ZOtwJMdsay/+z4FNt42lCPBK49b0Eh+DLR/3pv8+hR9UxEMccQ6ICXd2G31
xuHqHgJWyk31gumz8sAR4rd8ZIvWED/MMcLaU3SxB8SSo21ytFfkVPg+SKhW
T46e0JZB3bgoRFYfeYk+lvTGT63VXqAjH/VvUuS9merktoxzkDO3ErVIH7sZ
I9VB5q+NWMzBwfGD8kNjmVdJZMpyfn/cDRp1FbBK0Sn1oe7yVcB2xiruviLp
THYxzZ82V0U/vsW+tdygYeiXNtxjmL9UVj4ONvd+y9phyALRRL5wesP3qKtx
hVDPCo/3hIaVWD0dH5XUPBLb6uPcB5dvWd+kuaCQKVDxdEIyqC8Gq9/HjnVB
W8bP47y5OwyQOIBqiInUjo26k8pUZXWEFdcBH8Jchu/LYLM/4V/I+go3DIj1
xSOg0tZsiYNqKFO8K0bv7P8ZStm6ZAL27OYqXchQ4yjQzjSb5sAVx/+OE6vk
B71gOe8pSw0ipWhDPIqo0RRlWNS12vvNLvDJJ3pgec98ex5yt6rTjcR0C9qX
4S3oXdqbaUwL6CbRquzd7149Z2i0YxaWNesdrzq1FdDTEwF+RyxUys9XwTrA
rgpNkYyNivC5FzLWVTyZysdu8kXZmiTQMQhCy/8awXUQ3zBk4xh4coZCQhNx
5JWIxusVcBijJNsCOAyPpAM7C2vhqgpB7+aASyFGOFfNISSQZgJbSk/g2TdO
7RBuLLqyhprJk0WCIao1VJugjJl7t48WAwRvGuhGd7CDwvrKrqVX6+a1vl6t
iK+HST+v/6Gi8iAWZ6gJG9dfGC6SbZFBnvSAS47K/2zXCaVxBN/Ex/hIrrzm
dTPCEezNYfCUSOI41HTRzaeqv2Ts/SIMuT9CGebXjsY4yaor3ZkT+pky7jGG
ZokTlwNnqnE22RCufPeypq757mLhmjzkMmmZmBoXBlLfC/+QEuchnAr5GWAX
FgugogN/VOFpMFf9wxmSHypXFsfBFyHb2No1GnX9QQClmiWq8gbddDKrri8j
RPO82yTfNFbggcMscDLqU4pt9NyiCbh7BnFGrhYD4DtkQ6qWcC47SEoy2lQW
XuEicUC+TkK0DvzH84hV4Fm1UnR6/85TgJQoZgRR9aond8LZBQfu/FC0Vvhm
F4Pq0iEAiPhwTE4u+zq2KabqP5EguwrHnFzi9V0/OUnSokBBVW5oaWR10HBS
loWs4dgh3A3txtEpmdR/gt85FW9hwzaIDMpipmsYPPCg+dscVp8Wp/7OCKPM
oJH3wHFrj7OFRIAP185EhNo2YmXamT8pBNYe8Vr9r3qV7o9HHBXxO5nS6pC2
NzrGAl0YEk56uWEhBGYmm25e+L7HJFrwBzkNYmwS1tN1pBKelEoIdEbmpfPF
DSIcv9WrdArE++PvdoU7Aw0bGZJ2XCCCpsTGjYmshBgfKyBODxXgfafYec3F
KT4oD1qFP1uZldviiHY1wwYWSRU/U7cwxxgTfHpzTbw0++/rNoEtfIuU3CUI
40eGJCBSTvlBS3WtaZk2ECB2YVLihQMx8p3SUb9kQBtRZIkND64J9J4Cm18w
c8gvs2saUY8JL2AV0RuCAQXB/gGMh0d7uJdILT6g7QGEtIPL/vt962crR+S5
SoAGeLWEaCCjvyIhcfUfUddyGPdpuhVQp1xwWtpiLiTxxjR3OnZrQqv5e5st
V6BVgctEolFh8s/iVG497bQiEZeLoXyY32N5294xflr+QwaDRsjrWxO7xnIM
zqBM/KPhmiORC5UZC191O7Noy5GfKzrxfA/UTZu0JihukTacFWBdgjEijMx4
f2goVJd11/N5D37hhMbd8fx5Wd0Ikglntvl9tT+SxZzF4+knxS4zUjYjWBWG
LwmJMIzZNQlmtSWjQ6KVVQEPXCYhqGSEpkeEHtzRiAURlwhCwnquJLhIN4FV
ReC6dGH6aKWTbH7mdITkV9xhKvaxYw0j5QQFhjqc85xtq50Glqqj79diD8Du
c352syLFFL95gjQFDwtfViUHHWvQwUwhpRWBCdhKS7ODGpYTg42N/w7nS9x0
8bxhoTwiC5zvOMD00WhQSkDYoe/aayJMdvBIGhMYBUPWPEe9D/ZmBRPtaXWB
r4Ta8Y6NnPsFB/docuf9Lb4oAaZqWrQJEWQzLj2muitmtZRh9fjlmcTOnk0s
nmexzepohbx1Qx0Z/2sq3seHcJ/h1xNuWBl/M7BbGFpwOKjCQWiJ81rLCnqi
iveMWwgrzBG9t9nG/SBsV9mhB0zEtgi6ODHiklUqtToZ6hv1k9DKrjzhsx94
/x0FNcr1AdSV81f1K/u+J6ercIF0TEwloqirzN22Ry+H69fvMFnPKx46gdFC
YSZWw2VltvaNs7DhOgUQSapZxk8K4WO/1wuYxivF2E5HAlhMNciYmUqK+42A
+xXhqIpEKJTSguf21uj6HFjl2CksdEExOVVmtisp8eEpHIahO9v5f51T84N8
Hle3ZkaWzFdqRhU5NiKvzlnzQ07Hs5wo6vArf/X6Yzga8U4+EslsrHmP232v
UPm6k/v84/FqrceiYQ47gbcRRvPIQaCcBSb+j/PwVI+ceuH4x88cmNTA+70I
Mg1vhdXeJLPeqp/C2LdBxrgShfRNEtKT2kQuGZhJQeMM5wgpAEQgCPFpvtya
sOwYmAnR9rKrPOwOcKsRZzztuLIaF8jm/AOsVYe3CFRCtUczpWuVX+CnvV7A
fH0AjFMGQI6Xo9sZbq+IK6mRvylqYN7rPypP3mefrLJwAFHKgMMH+jjC0fxi
LElFaZUCglrEfRxZbkYvBN4Z8jY0nTAiPb8FW+Ut4dfGZb/zEjINruqIcNw/
Sf+iNHZQRFcg3oICizpnE3InYIkmr2sjvoXcHbFohdUJpEJ73BcNLw/BiE1v
WJdgg9GFu02lLNstkAuykVSjP0iizL1QsXLxLOBGQH8XW0II6S6qM0fvBUu8
zfxxPCwWj+G0PrCav5avZhVLHAEmlEZvAmy7eigiE54msJEDd3Fn8K0F4xsX
duGZhyvI8xKcTcP34wsSooP9eQ/H/44grMUerPraWm/ohIk3hpQWUx1jLVuM
4w5XBt51gtteJINjO71jEIwI5+WI+om8Viz8ABAlb0dt2Xi7/RSBxvwWzzod
pzRHOm1pvHXBdC72MRDMzTlN3wbO6TTe9FE4lAxUlM07xrGIt/fjXdsCYzlx
0t+dcnQ3CpD5kYXqV2lAkVsJuelQA7r/HG/EEOZtBzXGMF7r4O+Iooq1eXMB
hcqJF/nzElLUHFOs/sMVLvkWYoP6+HkO8CYwbSSrIsLh0XOeNc39VHxS8KiY
bOLtGN7A7v8qPJEJ/vqy4s8kgQgrIRyJUEZA8wq2WIsF02QzKTVxQVFG4p6Q
ncO4RcXPzIEUPzGXQJS5R3Eqs/69h2ePajHfN5Nekg3pa1hpLUjSw6jui7Hy
fKt7NErnWQ66BFgSbeUXdnRGN7ISffGeaPo6B6/lf0T49mUxDRR36fJvf7H0
YZSSJPFET5Sf3IDHRCvqki7W1dbYhioAC42+sEuDB7XpgZBy4JH3qoy8FyuY
+vZyWiSvUrQi43SKqMKuZxZZmXUxUJxGyHZcwzJ6Pixa4bl931Mw0uPnyPxy
NC0idtu35FG473Yy+twS64bbcFJqfWCbDTMK9tASQQEtyXK3iF/kJpR5O8ik
vJuavKxVXzTVOq9clK8adsk6fV5A69FX+ZbdLT5E1kxwivZAYxWueo6z4gJA
v0D8cJ63oJu8pu9a5cYZFgMxWPKgk4TNkFhy5kdfMdQIvdZJ8Wd45Q9QJEMd
3cCDp1HePGfco3pZXjQgW0GQEQW8adV8zIKTcT+9zWf3CTjOOfmEvRSHXBJY
tjLh5lJPlynzy1C5Iy6JwmlJtMvconXJLQ/IY611jfgdx88bMWFMXW/S5ekU
ZWhgvyrvg1l9qoG7dl2KM2wKw3HsBOv0KkKyB2aidTPV2ItiqL/0ZRuq0Wx2
sHk78zWuDx1yLjLvq5f9eEVhh6LIjBHCiLT7wlxK2GCPGHXzrqcBDmQiJmy7
2thn7JRmkR17kp/5zAWXEOPrGNtfOnzveYimmaN2XofKcWUqzjAXIT5A+rTl
3lUplxtRa7dg5OSAnXHJij6baHDswq0ArR5+L32v5dLWdrObgwHpUjwj7UV3
qXupNkTBF4pe+C9K/C7v8cOy84L5S6zC/bK+YKOwucoS1R85QaZHLsju2t1Q
vFG73g41CKkqea65Yk7QCwQ/6QCOANM914Thr+5AT2j1xHyJ2hk0lUYefKkL
os/qmwWbBhBbJ40srKcfWq+9kTliE3U60EIC6EZ0f4S+K7upC8W0TiT04GkX
LLQzJr+zRwDzh9uI8MOSQwf2Itxh1/90a8h9BtafUXNDJfjr+KMFwG0Lwnme
o15FhcA3BWtt+/Qge/7aLHByS+uUGduh2R1UUsoQRKDsVcUHjKRgI6Oi2+UF
oUrXTuv4SUgYslJRMbxB5rJvcvlCNtvS7E1A87G+GXy5o1eDd80FmQt840T7
G9S4AD0VJkq0CHMPUFB77InGWe1zG/k7M1XCUpwsEOA6FhDSxgEGbQ6U0LZT
CotzVCicKe+A+sSuEN0MlSUejn1EfCIwwAEsSDWeRnT3vs5mKZnHlgJvsKe7
d5tzmkK/A367Q0sBNEbcCYypostkOp77vLlE5tVe0mrEtf4Ba8LMiXYcjXQJ
nhYNx5DU997plt97qBdeCQM98lfRfrnq862WKr/QGvQfCo/f2Q1SaBU9TB0g
VEcZOfJ1KTpY3Z+buMNW6pjlXsaEgR9T6hH3ko2gUnfAsjZW8vnSUyhPx+6y
3pk0NpY3Js6f/BLTfs8a/xFuoF9Ku3XWWYmdaGgAB/cZgkON7QN7XJa0JAfB
mPFncPgGDBdUmYY3DXDuePcdHSLWnY9PU0PY/5kDpxvSwdPcP9Av8D3YwlcN
Nn/YQhkwUj2oP7LX2bg9wpI4wjgy1Doq8/0CBMmTe2XYN9vQpZ5qJlrVS2BI
hkI5pIqGy3cLS/mkVmEKQy5Xs2fylMqrw9GGrZxeVNlvoryqVC3kZ03Jmd4Y
mjbH1RhcnXsbnMHsikPSkbAsKSWjNfFoiz5PjilqKrVALGMdyib4xA1XgwKw
xINj8FPqQyTvTpFgTxbeKa+ru1LO9dW1BspXTmMdBTTWHpyO7GHwgkFy/jI/
FTTzyPyU0PK8mSx1Dwr6mdqb46Xfm5d4cmL8IYJQzQc+afXAcrS3QMZQt7Og
IWW1TBlPjUuDIcaKNAXOUmyyVjEpc4jodvJgzXWbyCfNKnH8ADWq/YWtHXcG
rZg7QrGxbgtuMNiLNjEhmHS3j1Ki+t2EyB4FgFUBpK3SYiNxDMowGkCyTkqn
sSbXfKa54KjGzKmJ2srZOX7YDHzsXmVQCyoEWeOjSz/2fww1ABH0k5D0Agq1
Y+3K248JWqf+ZBz3Z0IMqaWGgXVmT5JJw+LNQv/EXFkj/AHtcseDBydRBLQw
08VM+nMev5Hrsun4fyrHFRBpETARxGLsiACPQlJY/SqLpU9R1g/J7j2SVaYi
FN7Y1EuQyKNWQmzbnCz1ZOXfK26+giO3vXe3iRo+PGWrUyFnldtbh3l4kXEq
YqLB0oT/XmMvToOughxQYM36Ne7V2ilLzyWFxL1WE10w689nmYCU3LJj6/8L
n+ufGLQ7TjbwiT9BSFPBfXMopZu45kDAeVbFi5WIZAjQy9o+Kq0FW3ztBPgJ
tt0kf0jSnG+otKN1g4j0UpN6RoM/Nc762wbqYGKmEMrJMjRKX7RBXYYpMMdL
69+wVChBTXI1Gy7QqMNN1ak1xNezdqb02E4i/edW87h0cxekkblskG6bZeo9
5TjxvI/bATsxEacGakfctYDWHgS1eT7vKMAkaDfRivPqz68AFYqfRpftTElg
P0jN7gsjLzjpkiS6RURItPO5EEGsWO8x8hzCDql8AqZIv8ZfNHZEML2OjEvw
CeWhEAsNj+3BmeCwVuwlsjk6OkG4oQuicw3/SPujLYYAFnT1bsPzfZTuxep8
PwgBIrwyN81gXu3ZWaI2GAtLAe7ONR1jN3i0XwLx+vLNbVfibFxGV35sjl52
WjIpLgTgvQmveEp6flX5CtnPcnAEk6wUG05oUn4drvs0mvRNQJbJo9LfovN9
gr54gZP49MoSPSj9Wp879TM+VnpQLQE6yYPy0DVeEDqw1lJDLAES4gozFNAo
wQgwlvbznYnA5QdDEIPPHe83/jqNL9InxWGU+l5Rpujd08WdK2LHK2LQxIhq
jsiL9m4OHNEKZ2F1/SuF99k1X6pGzWgkJFWB0Seas3yiOV+D5AWNn2zs45Yn
ZbqOOxqMF3+pM1lNBnYuOPCMFkAAtHIjjRwH2z34mRWHLCG0u4Ye+TLmvfLR
sJ3yDqAgMmW5ZZ30EgL7iC+ULUPb4Zj/H1M0SM6YVLpiT9wv6lNbFd51yqbY
BC9zxUb5BmroH1z8AGFshXbMlEhnvy1JpTwMOa2qNTv5bPH36vMtsRAuuTsz
Ea0B7bWjDyl7uutMb0x1bLrugatKMEcYEyu3OeiXIlsSaOfpDwhyHWQZycXM
XL6wcu7l0lKiKOElS3WHQoVmgIBXGWfhMd6iWF1W9fKIz0dm0otPQkVsofKa
CCGprGAjiB5sEvWIxs3+DvShn/PP1QHZmRQWddx9QRqNNFfai+JaftPThVzs
3o5FVvo04bkguJfwPshmKUfUzq16eRopQMi4p9yp79DqQdyi8nTWFKpMruVd
S/XgVAdFKSNPp5xeVun2XsnHl/RKbKOtEZZg9XW7bj6nVau3hmevtfFz4YRi
fcisTAM76NsCvTN2+rJVHKksuAL2lLehv3tlW0iLUb4m2b7K/JA5DokGFmhE
g/mxSOFv8lpPuNYimWmSPYmTk3vsyv6M9LHJqA1E53rm9l0bqepAOvqoYoNq
5OK6iluOEEsuZxknoAXrQG445XbbFus/CMFyHO+pX0ZPWGK9LtIDI5VoYqh4
7pRl1Gl5kzktN6ttDOcM9ae/ojMbEoX+wn1Pe0YbOOO03tRxH5z2CWJudvhT
s27R0LUPsmZagys0c1DyI5Jr9yPjcs0UIQp0w+qd59vjC5h0aQR4BXkL0nSn
OYMbMr4xyfUDoPfpOM99eTFEcp3pTvKWwK2xzCx87oFeWL8gLKPYQBg4L2M5
7bXGe7LKZiHyq275TDmnoY9Wb9zdG8lfm5NduTNXm/LEbdjF+pcjqfIh9/h0
oeKsA8IgANTYdR5zEzXdqDb4/MwrvwMaQZB68xDVIdfkz4xwxvueBvGueT01
yknoD6VrjRoTGisHbsnuw2zHXjjCONICQH3FJ967YhEvcovtTND9HFWFFFpO
o53/nLrrAGMbMAlmXELOX9XHdIJMo3ZNnpCYen+dbyS8Rcqs7gc80yPV02ct
1MVPtjp8J9U5FDgiPU3IdSCcNJ1uie32Ev4rKANqccwqMA6RnozTqqfQSEmc
i8BV1uEuF1g6xKLGx8S6I9p/HK5NtY8+uQo0zINi0vxwBCjcxXC4W78V1EQC
T7J4Nc6D8a08U9AuYFSQdMKExE/trSELPZ4/eU8B8NLMB+QAutajAS+YsN5e
iYaYt44J9EFixj0RaxI3LDtw/S5d1Zr1+DeRRsDT5xbEC8JoBSPSxK4KFwR7
ovTX+HSft+WcgH8Zy1KkUYTCT7Nmj6ocfleKm1qMS61XlB9cfm9Gbi/dZC0T
d0zhPvqPIm1WYZLICNC4gu+YcxrH15ymwSHVoOFggRdR0AMVMiC+1+MRPgyt
fQ2JZ1mg2/un/2GFgkwhwWyLpgt1mVcCgbVd1gb9wjlJ+Wexw7X2YTmkWUy6
94wyxb1e2IQhXC2XU+7qwLP+amJA71pcaYXQtYqPno/HfwjkCIbT8g5t+dcK
BibO9WVz3qIYdJA2vDEqk1u7ulRzdObRUR+j7PGuLr4s/BPdhhb/Oft4ryhB
0n+oht0MoUZZ3EWhuyazgKiynZm9ZfrwMP8sxmTGOCZFQVzJ65Gqtw3XsJ5w
U7OngfC53aKDDhD92Zl1bkEQjzPXa0SFDnaK+OfqMivborLWnSP/ccq41wcR
TW1P/vR+/Ab+XX7nzFo2Th6reiLbrwrZUEHKUz7MTi992UJshTc2Gxxcvkum
oKKw57acTXIAxk/DTt/2rf6+MkBZg0FEO9bnDBPxPWenxfkIY2CKO9GfkpnE
Nd6paS+t2UAkuUvNdTLsTvYv9uYpWFv0xj4K9WJptoECM3pKdcJ/mmhFMPon
uAr5vmxYyJnge45jDIErPpTcbnby2C7Tu8O7L9KJsoSFw25zpxVN9LTOjDp8
rpGYrfAwUm1glI5XnwKXGa4QSLKrxzqIowbaiWeb6zzAFB4RStyNmlMnsffm
d3ScLvJZ8cWq79X0Ei40MJX+Hh9lP7Ky0QChmSX/yhBG3pLlD/w86lI4el3Y
PvGLQA0688xUG/eGTTGkG4GSFD8StMXsdjjZCgaIGrASQiG+Mf7C216IriNH
cRUbYbRjNQvOdN9TuBK0/0zf/5vtQDIDmf157Fp7pKhK77LIFTbFRxpCVcbQ
1A8S1s2Z5OJaxiEhhzgdb5KC7fdofLuPS+8wSG7aAls23eaP6pMRJc/+hmBr
mMASv15lI57e7cUu/h6p6c3rqviQfbKjZMldSPxZJ6WGHcd/F5RUDSK3jfnM
/nwraLWykbgXZj/TtDI60wmr8Iz02eyD6cvwLVcGWp77Kw7D9fg/RdBkypeH
k8Aaj2phY2imdB7ELwGSoW1fHz+cG5fTTSc7tIAtkeKa7F87YsvMYJtcICgR
UskLHTgglO1e8ax/WSyFs+x/6i9OydInuOaP4Xhi4Gqn6fB+wqI602NPKikZ
UQ5RIRq4uaVKR80MmKdivdz+vwn/2kZ69RydeHcE+NkRiqr96uKWSskyPdeD
4+8cDhH92ilv3Hu263yE2lzNaSdyu218okz3H83O/SMaw3lVUhf5xJXkp5mt
pFAKt/+Gcpg/jhxf4bH2hPXFJKzlwUawsvIjjuJldyeCLcQ6WCYf035cq2qy
3IEd7OC/AMU+tWOQYBJqWdjfpEzxC0myhRu9CpHJ8oNTvNLhgy9rGwExCAey
6CD8R8joR5KJq6YWbE3E9raHgX7niN2mw6MoCeRulRXv/F9YM/hsRH1HLYd5
EYnmvi0a3YYtKmpJSB7cYsmehDxmyjM4kvYvHf8ec6Tm4Yk19iTYN0vYFTDY
tWxkp8z+vVtxqfB8pKW88oSLGHj7jQe7mP8BNHs9sl19KY/fO6I3ge02yMqb
K/Cni+bFkUcrDAuULZ7eWBcOdImvP6lsHzidlnpy7ESyVvzG0bdwBfyOC1oi
/HC4bXMva5QzCvr5bG5sTGtCNl+EKUQZB0ZRE451b8ijLcQV+g9JBQZ0OQ4a
afk3bivAvkeoiLm81LrgWpofsMrQNGEwxfrvd2PkKAcTB1l0Fz5p11hkJrDL
HM5ZzkMpKQuVOWEAfi2IJU4AjTP0c7ukC6Avp/Uoqb6sXGbbaE/APjABS6dX
oGcFLFhqdbGKFdg0mPBo5z9hLGeXKW4j5vGhTlY/2isB6CBMg7Dp7hQ7X/7F
azwoyTgPb6c7Q05/2gsU6VPQmOB7zVhfEUhnFqzDNXXz8j395BJVzBJFauIF
dkSzFyconBb5s0si/kk+g90eby2H5e6fCJMLJXmLEuQ9Tn808VVMq0SqYUYL
lfnu2/b4oXhF1uH/glc3pjPgtN65wZt45qOwlA2fz//FJ3wF0aYI2as1ZMKl
Ef1Y68Sja+6LByTSv8TsX7Cg8BNFULBlzzxMBRMnC3hfgKwvjuxf69vCFPLy
+cRCwiOa2J5drMxvYIJTBqquzH5nUpfy9gv1NBnhBB3JPWsplvz/nUvpse5G
s2RWR7ddZBGT7afRcHmfdIAHaZHlIhlU+utY+H/hPKZe4HDZf2jBFe/H2Qir
BiyRmJBendVksmPPJoGcQDuIRcRCIKZA5VG7J3DivVFx3H6StEFnnLtHJnNi
LxKlP7Od1UFhyt3THoDC1+jSVCHkR2tBVLILZbpXKsvcQArqRZPvWu5uoGL4
U2na6qfeNZf/0bsz1q0IG6owbP2kOSq2eFFh267GcyaMrb2dfMFWgBJ51LjR
ngjiB1YHsPlVruI6SmxqS5pCRKM7P5pltRtdiSaJrYZsvRbR2OGN3AK5G3Om
MkAtGxyA63adHTBhteeb3nkr73qe+Awnmz0QYnHnplf6QYZH7JwALwvT1wTQ
cqU8oZ9bULXHe8Y6rThjDs3QQUPgsCks6UIAc4fNBRDsud7duokDlYt9Alcs
iB9TvxOyhGNipO91tkYsNPjfSMhO3XP4wI1KaEWK7WyPiXSte3grbCEIQ/K8
yqpMddad147BYK3MtUJ+Pij/ET4nsNhRFeca114QbmkiRKm13JDc0l9uXEnl
yciQlabPxqnnJYxPsFfYxyAkm4liOfO+b4lQ7M/2ptLgxvUGprSv+GsYXW8K
Qj7wjzj2iCZXU6n42doooriqpRCqjY5u4zi6mvVcTT6wPMxn03+4QPMX3ZY/
AhOLo+J4PcTekKYmtREIxQDKeEyFHhNJTBe4vkB13dlzRK1gX0R7n7cChb9k
JUcj/4wT/k5rFysfbbuD87/k+7WM/uIZbQkLX/qUu/YjbcrfUKwuo8AmpIzX
9UifSc6jzRTaefN+BfoOLEfPPmrua9OwCOQUqFKOzinLwQBnhH1S0YWRCc+w
+65HrRFLe9bfARVgRKgoxrm+0CksG9Vs/Sooj9c2MuKCTrfVYV2/9+IDvtMI
FXkHfCRwQn2P7UE0RzmQurPsSkQ8TVJg+7KOPT06/3Mt1xFwehemJjH248sX
wcAiX9qYM/Fch7qxUcwh40X3jGv043vHyx1VAKwBFgcsoGOzf2olly/OGRUa
l349VARgL6Sjvi2ti9FohUkr70VK9ifwKzYkmwehRb5CCtcu9IaWTWl+FCAu
IRZiTLn2O5JxSWPiptq7/gHW9crKscRSbKkYdfDw4Jz2ixArDIGvNr6+0ObK
5N13GkQPhoDQxXaZwtTVgoRAuMCWoWgAqTf1ef8pC0/OHCod6ndmoufg/tMU
e041LTc17g9Pfdq2N0J2jE8A5gze7VixUUzJFKYk03Xsmr/gCtgNtRmiIF8+
j8YT3HotHsrqC0PfGM3YnYdjHSIbDu5/QY9ha7Fn3PxV0Uo89p303LXlBKLL
knktMJNzFo21ClzY6io36CpjmGBFsVPan9iCO2c8kF7oG+mJKmVcpgEe5x7r
YrhcbZWgr2hlsTrnypC1LPLo8oOBDlSHpzo37fup7p+p1I2qLsVKxVNArHYr
T1WJn9uVQCOiBvAmMFqvPqi03oBImoxuyP+AN+Kvs60wpiXAVKT5/CZ13MN8
u2xzIY3VQBcbyVzUfaQja8BBsvMMG06e836JD8XVuftBmWNfb+MwfOzl8+i0
2x/4jfzKAn9MQRkGz28Pekmk3SA8x+eST21Gx4hgDAGT+yvp22YUKCP0GQ8b
92kP5mvAbbk9DzoSrja0xbDu/XtLabMTe7/A6vlxc0+ZkzAF33bdeuhR3GoV
mgjlEXD7ohbQAvdBuB6r2RikUnmttXBGq2AMbqWttbO+O35YiiM8UTi6yV1r
sw/sfZ76UDZRoWTVaSkyUOABIGF+ECLFhV3yUTLeAX3YCOGdAQ4JdVbqWStL
huE43v8lCA11PyeqkAZFfWo8vWBiZZH6yx1kGlLUfvXLQoF3dSCVglIWMNV1
CkrZyLC2vtw6sZUqjYgH/v3RpHvFDghr6pXrN0ARWlptuJMK8LTREHi93KDC
ntIIaWiG+i7DjcsvYY8OEHNPuv8yfPp8CIdykd8DNwOQd8lD/Gt225rWxlJz
NjMzJjyiYQwhGUBT9CIxTz3KT+sDraIIlvxHifYEqH9/DUQNzK2sHnSm9YX2
dFZRScx0IVXQ/8D2Cs+A1HsqA5u8J5twHPdegLNzkNvVZ1YqRv2/OKDUYgSF
W3eS0WtfHcxtuw56I+lHhgiSP74O2xu0j5dbn9xDzbSuCwfjZkAOMqyUwsru
STml/UVfjRRh/C96i9enSA4qxeq7VpML116q2GUEKizwmAW1ijQh5uVtDsSy
yriEsumwYjDObh5Lg2oVzA8t/R2GXDo/F/CZLaK3Jk6xRHQuJb1YM/16075Z
faA6gbuIvDZXZ+g7FOe2NT8JMzyKFSz/klxbkegjbwgD3DobKpM9QRHlbbwJ
vaAASL+RnfgWvP4su7cxU7kWz9WspNTZGKzGiizSemtRbhFhGmHktqbRPXXU
A04/zdEDlD7pNqDwg859vhtYLxf/shCtKewgeA1qioq7E7SpVq3qmS44EoFB
NtiPkbfJavN9uegIxosGUaAkFzZeP1dvAAheceOxTE1uB0P+UU0Q9R/3K6bq
DZSm6/dlDcFVkLq71NAgPJxwyOKZB9cy35vmmDOCjmcfMhTJ+WaLtScYSniT
3ofsorz0xsXY5MkkbgjOVcoAgZXbvCmqsEjQvkVt/6MH4MumzOAVVn7iyv7T
HewLAdsesGvlEm+eoZNKyWyMouBhDxwQJzu8V22UaFhT1EKFtx7vPhSzX0NZ
c26Q4V+qxm2dHRfkq4E9GiEoEahNdewYENuG2B5e8PUD91jOd3xhqGBDX+BZ
zl0TS4AOvai+FqJJpbVeePuyiJCcEb0I3ipWGqEA1eNqxlFEb91KJI4e9COp
Cyq1Zq6Zyi+fOSV53SIH/quGUj1936ipNj1RighFwF4/d5NPNcGhsBbColbf
z6bWoajFmF3cMl1PwzcEWwKp4lQR4AmStaZ+3nXRCiGUJTlXYtkFh/euwbCw
tJBHaWbsWkCgjR0MugVzs3zhTVKyC35bVCPcHkdYdZJXLG1rUndxGYvdbKPO
9TMAEbsPyW4ZwjapELun0Y5EB3Zd9GN4sFDBkaS9rpdzxqcEiqF1f0pM38SV
OXkIDf0WRgCsPv0Ar7n3niTgZVekEabzE+CeYqH+FdTS7+6vAMVzgYzlmjEV
9k6v6QBnAj5ev6t51e2IfI2CTswhWr6HDsYjyMGrkJUhIatGlyZysTLA+pc+
LacMlyVAb3URLlqWj7TmHJ4ZaNA8Sx2b6puo2HB2t0Z99eNEFl+bXLvtZWx4
0/rla8lS4vKH2BzHKklXHQIkdWut/sAggQELQgZHZZ2JnkBvE9FeUNU3vju+
BVEjF5pu1Aj4ZnendVVP4nBDUZvIoFZqT2VsOwSxKlD/77O52cYq91zno2bo
o5fEqlwUykTBCSHagQw1x0n2BNirzJIZ/VgTIZRSol4AhVIDYvadhPx0f58w
uhJ6puuaMPvjjWT3XuG7wEbU6Bz0hoPFfRZ0paVZLUSDIgocrlAVfPRiFZxo
J82+0lI4LnyRTmly9x7ktigA94Fu6l87H5XFhL0m+0iRc8cPzSFt9TsIl+dI
+1mv4THNgE7EwNfDahhmyDGna20wKhF9IO2ST0KnUYF9wRx2KTBO46+9t77k
PeJzSvsqndnSwM6gLtVYBfU83+aXHTZJjwqy3mm5TNqpHQsVveLhoksa9ZF7
6SptnxpqLzAB6tvXkzlWcyqrvi6pA49OaJtSdEZ5TzMaVj59QSJfpJz76GmZ
hPqv7BuaNR7hIRRorPb62sckMP5EifTal8hquObTMdZJaeCOd0xw3oTJ4ELd
lHgIIudD/8uPiN2r9U4X4SrLWkjVGUFVBzyDCt8n6TEZwucYgT2kulDfLaoS
9sVArYEm+3WGhpnKTN62I7fqhXYCLkOldNVoHquBz2iJfpPFySu2OzoLt+fr
eBkyP07M9YQ5G8sclpsjZe6Vx41Akow0Zoc9E2DrbRrrC4B80AKFdcF6slNF
xeD+CUvUsbW/rY4wFkDazJ6qaBXvnk7VOtwCJnp+is8Q0D/kEO5pL6Ureudf
WN004rPk6r4eXH1NfWNytroxiE6Xb5Lmpw3xxBJWZIKuyEWowM6uZVTcFMYq
xHp1h2fkQClLiqqajwK/5Bp4uyHmaENv7thgS/LuQQBOKBLcLt8yk1SjzkV1
F6gEk9jCZpdR3l+QrzNsowbml0FCm6U1ZuSjeQb6zU4fc0ELInFnkbMSn40U
CjpFcJydMxBRoxrOx1VNlZ9djRHrF09t/z6Qw/j4TspSgMLR6znUkrGxlbbA
09rbed8aLAbR5tuZdE1xUhB7t64tLJIavZHokCSZi13OhC7Rl+jyPpDoPaxh
3MZ4C3NOqDAU3ertGVSAgI9Yxp3eU0XiotNQs/LvxjA7DYXYxa72oOv1q0OT
r/ZsVuJJ8TyP7jHeG2s+OjJSYdmNhPtp6uo+QBZsYtwYG4Ev9J+529OXLinO
DdnqvWj54ST0kLEYpLFTdx65XyZJjIUKTcbDKhdbcFyFkQSByFx+0o/8yfi4
clEKPOWyRY/iNNARzG0VDG4EZzZXdM0RFgE2/ypp6JdeeV7EsF2iLA6Mn7SD
dzxUymcZc1g41+3PqBOCY9f/cjN5EPxQN1WPJj8CmlXnADfaXm+WyKCNMwls
tRuaE2oSdIEvyP8DjbIfqdyQD4URHknJasgFRMyFjJLv272jHsK3KEyS/DlV
hkfy12UNpMLwTs22Os+9sirPEQTrTISR23BSt6u3Sr3d1YExixMn0bYdGGbE
PyfBuu/zoCEXpWXcqqFhE0AHB98Rgd1Tb5Lon1wsIKNpMmmDML03QiLFBtPl
Od8rMoQ7kSMmw04yQhuPX/P+BPpCkgrV6HW6INEVFTK5XkGM/dJnI6bHl4EJ
LssA9L8uZmntaBWakMlg8YU+LfsDBhkyRB4BVr1uuU3KE7H863OnZS63R3f+
g6xi3bfoMFpasDAR9MU/7wl5VI78JNulkm1FAWORDXCCOwIkZZbv4M/BFFT9
CAsiHml2rsiLXdT8SBWPM5UnxDcZd8XbEFFvi42OXXJ2PzWDGHMeNae1F8ZV
0H1KuaymvAjZ+GyJrzCUZfseQwobyBuwRi4JjnaFLFN5zWZ1KraOPKoXyNl4
r3g629tFCHuD11XLkkYLU2q1CiLEgCECtRuEJ19vY4zWOvx2wE2bvIGpYPez
EjeIETR/AAgsun98jTPkKxKnsk53ZvYXsOySqmdW34Zg/Pi/Mdy6jiD6GhQw
VLiGRalvwXrR6HDAsHPkaxJtF/Uovtg9bJu+8gi3Wv6aMnehDjVGLK/FZj1N
kHUUWt9o+oibzIKjq5/tgwolc+az/+PI2VuRvZi9VW4vaRVbqaVm1e1P9qI0
Bk51pfjKShJGtj7L5qKTaAD8kQKgV0OKlghEz+NhLd/zYScx38a3bTDkxcTj
AQA83Su7gRlFf/JeiF5rreRucpJSHTMCyZ9Yy67phj6DekoEHFKtMe0wAqR5
AxwgNz9nmIkf3eIUFcGdWTR9RtBIzJeZ3qWxtpG3Ad2xiMbCO2hrtkCJvKH+
1aBwNX7Ap70My09l32bBiWTbbC9oZGZCWc2srJ5NOSOe8Wabv2455kyBvNzh
pGjwE3jCMx+mlW6HcwJeGF3u4pj8DT8QxAdUfQjG+p/tUblIdBVv6tgbfaMp
77oPCv/vQFNnsE6PlR1spcWX1B7b+OaJKFzS+iAPYFtJtLWjqZBy69LgdrN7
3EHhQRaNhdCXAVcgOCE+KsuCK1tj+FPkH9Whk/sQO5O/cV/MDLEK7tNsRUHv
gfiqvTNavsb7rs6He4jssNtMFStIpkYXD/spBQgKVTXCSRwK8plD4Al8wJix
BbYYvr93E7K98opybjuvUkAMvYuKvSfJ+5OvwY2/Y3nI3ynsO4zK8PoLYFSa
5EHbOGA3W70P0oq0Mddbe6pHg1sxN9S+WoPRiAiXqhPTUDPyp20pJxrN3Eww
ilx/5T4QovSitVNR/NWokt91cmSd0r2ubydLVjJd7823dU1gOgbQW8IxdBeR
Kmla7HezfvMppUQ7slWsSLwSj6GHCZpaRVb/Zg3st0rB7lyu2KBEZ02oO4zk
6Yf9eEaUPI6HgwhZzLFJTZXHZhrom2ezhZoUDqkGwujTrMmkWbr5hEUxBbOO
s0CilbdrkRTuYy69b5Mmp4yczS5geJoEsPliKAwLuim0sUac02YJcl+AkWDF
67RUs8P16bLK1WJ164dM0GctrCAyUop2kPsq2iiZaLmUygLVO2mavDxT5XOP
pfxzUwqtuTBxToHeJnig8sqjRmI+GSNSpymaHjmCpdN39ygZNinX7B3SIth7
8UlgYBjQMprS5Un+mfol37xs1WldLluE6T0SWfY2AlGuHpiTyKy0WUm+84Co
FZsnffl2H2ZNsl+kjpuYrbBwdGUy3RIdiViJItT8OzvhfIV/CHC+vn2CuwNN
aWANJmfzCzsyu5tGhlWCd66oWDpMpWscM8GHEBVBSaOFrspohBy1w3Iu4TSR
u9mIlx89CU9E6a5K0nbkvH5hbNwp1qEDqcoJnIggCZqBBkzCh16Zth7IhTlP
KnSP8194MeT+hOCNJ98oCJLPX8rmA1OUgaCUdNA5IUUbTDYHr4rQWbbh8m40
tfNjzir+Uqqchk/Z/+dwvU73OWW/u1NIPlwLBkO+bVYbHOpgDVFxrsi5//ZM
Aqeocuacu/tM3Oa/9ro5UGoccIjoFI7Xr/qIpaCowEOqP0NdfAAQTI6H0aHK
/0HZcJ123BHxbDm89LuX4Q6j8opfJAy3ndAx9eqLd16XnhQCg3lwfZYPrkKU
imKiCiF+yXRB3KHzcK4cmIsDoAvANlalno0JnzgvzNI6wiecnMR0O3T9Amr6
2dTyBP1vFA5EON6rwSnj1sTPi9ZJxkAI3nKZ78AcR9c3XeoZcxuG9cdSKyr7
8do8XuW+7GqxnZdYMjICjPAQmXjYjGm/Z7xDQQ2BdZYigX6AmWF9Cd8QyVo0
5so2bSXoJjtPyOa9dVAF3Q0encrj4epY+FfLO0GnKs6mgBZLrEtHHrzhbUl3
Q0ecYQZWkEjCIin0qGo2BsdawAZTisMcKBtmnn4wUSogV8VYzfPq2A4baj/9
tYeF48IHb0lAwlryQ0FgoWNnDWvO2C0nEl7xRiTm+uTbfDhoExJRc3JsDzMa
IxuiUJva5kfg43OJ2AmtKZzxaFKrxH3UyUHkDr2O71xJuY/Ypg3mlHXNCdfs
iJxTc3O6tgXYbcFaHBFZDOc2A2fCCSsmC9BWtDV1FoLBUu8JNFIUDSeFgvz2
PJ8x9GryQw5X2UzOIiiBiNMYn40y6pdfqdGSU5gagKQ6Jrzd+rsKjG6DqfqL
bSI8+jH3iAZ/03HVa9Mi9AvF176JQKDd2MV+jZJQKKvxlUuyiI9SE1CYqqfX
uoNbgydztAxLLMNMpi02Ee0MRkz0luwAwFjU12iqKweUcUxqhESjEapuYWVu
59xVl3C4etYtJzfaQlUYQQCZ3e+O+RC0+xKhgxc3/k/cUsXUVNv5ing5oxhi
cQPb8Vw/eL5FeJhazzPIr97WYJ1S3VQhxpvvCpRg0shXxk/zTE/YvnIm5n6A
Xj/3kH9MBgo/a3OL63glLs/zg5AEJg38TC8vhe8AKavBa2jPLj0yVvhBOcc9
xh4SVGgO019aLB4rM0MlmmoDY3erz4WOk9+tgCZr32gjc4ocmfWrGkrI+fkj
awHFNQz7OubQEFjeXvx485GEqrgspEgrA9nhVmEEu+DtGulb6Q4uYUTYIHc0
RQjYkqVwm8TgzjiHFzm0TOFFH7e4lsDltJAsYrl+/TDyHcNgMV1KeF+/2Xas
wq8rdqOfo/yhDmG1CbDFFb0Qz5dvZM17Tb+0aiYqAB8h0wIA+vpM5JqnD0Xg
TuO8b0EP1peVYQ8J/Qvn6EWeJqB1JkK2PF6rAbNrNaPsJxjJp1ZWDJp0mKDi
iDSW/3Z+V385uBMjm9paN9PzkgC+rY/qXTbNLI1gE68/KYU/qfjr8uHL0cYc
oAuxusyoTorAEcQoezBJcaakK+4/hS0r3QvSNBPyRB1R+5hPjKWtvxGr7Qgo
KAQIzUeo7pRXp4uIc6xSLmj0FSDxqvi7bJVI36XqhZJSyUD9xoxQzzrw0ubk
1XnI0BrdiqidGt52R32rbZ80eNF5hN4Ut0D2+xRzsa8yLW61PauMfO4X2oGG
Sm3xTKR+6ByqbrDYA9pDAcatg0BkJWIxgASMJAk8ekPQGyNKNmbmXsufD7x6
JEeLXDmAcTZ8YPi3cCMwURLwZU0j1XH/k8tfOMYP/5IJvKAniSlgpihwf84E
crE7iptge8KeDHCL8hsOsaiYCDLit9rwIhZDT9BdQpxnh/KAGkyIqC37PGff
ZkYBG/mMD/w7F8UPXTNc92qmjut5mC6Cca7m5oT5NDiKhuTkeERiIO3RfInW
vJUHT6G6Gh8IdVrHdUrlfknCpwTgXxvNieaDW9l3qOTxCgCSEjpqQa7Sdjed
umjJiq2vLo1Y47yPB/ttfo0Osl/nIx7Z327/4Kg1So1UnjmA6yyjaJz1IT/r
0kafT9hQoorLHx7OAvzIbJygN9nSkWYQ+B5uiEYiBVzCAzLYSLpMBQEqJHu6
FJoLZzUm4IS7iTORbIFj63IufeO8dhCyxInIpfNtI/62WG/bdde4VjLivbIo
SIa+IxLV0L3FFdEL80wvbr2aI8cuncFkvvZzVwhoswwG6Uo4lQEjQPi215Rw
CNyG5Slsv8iakRTZYpv03a3iNpPFAbRSQ1psfWi2neDvQyLs1wRcUxQM8GNF
2EmjTLgyQqWI7BeDrM3QvR4Sf2ikTTpOADpe2ZigVgdVYW9KpAHNpvxi1R2L
SnExoeSyYYWOFhQ8g8J0vNfMt0Yvd/3kyFn6G2ObUg6wYXwPqKobOUrvRDAo
UbBxeLCuQQANOKhY8PENs4aA7a1p+umdX5+Al4QIK4vkMfbE38mF5I3jeoHL
bctwB1qFkwc5Dm2yk1YvILzSSY3sQ7UkeOcQgf3/OjF1T9wIsqIS4jLoRaLA
Y7VosX+BfQM3YKgP5T48SQiQVfxZuFaAZeP+eOHwpd4tE0oxDoz7mzEi8GwU
6WAwvPyg/1xiw3+m5OgegagV1tjPrP5V2F/dvGPP/U7JBUkC52vccHuo0GEn
PLNjVwu8MBSMzHL6FL1dc2N0M2yMhGb7RdzO+S/7l/revABNnmT/c5BIDcO4
aesuj/6DcJmaBetwc+B8xKAH29E0eU+rplFGoV387E3QOC8J+WQdnzHFK9uu
eOBi3PFygz/qNwvCQ/wquYRDUV+VgQKPlUmoj48W72+ayVPS86LG+CwtQSrD
XD/z1fgVc1Jmc0eeOe33S0gy25NkUn/yd2d8Vk+jGrMiGDd4QrpOWcVEDzlu
REhr98+Xl3gME4Szoi6KpfU6wK+0NtyZrTP7zbzEM2ezEue6SCd7YQysFDll
pTRmKpkFmLTDSTs+aMv9KPlxzs9AamZknaeCIJHnkCRhF1kqNG5QyYMp2Xyf
PdE1VcvRQUUJungfwV8ksNiJ/UI35dXG6LMS+AxUalQJerO/fOCE2EYNcf/q
jYmxwdv5jdmBjQq4naVXQx1QTDCdqpwfJa7uv/j0hl/HhkDyyvV1USfk08U8
3Bh7C8DRUAYPtLLA4zVKv3DIj8mtfZacUpg9OU89lt3mUvavqU0SlnMvqDXl
7DzTjcmLeJDb332lNCIE+/nVHvGm22fv/i8IfHnTrm3/8SojCO51ejjpzI9Z
TKVWvqHiX2LNSLBsKTxOahNrTXZ4TFpMqYb0RwR9frWVNYX8VFz6EY+c+9C/
Zg+xZuqMA45pb7TRFQ1F5fCsyKWDcMkpX27epooZ/pGTOQr/ckJMgoP9dpdo
igmQZLEcjgCwC5xtHuBYk0Fjr71vS+9ZSU5kZ5z60uu4UahyWA/F9gfxiSIA
c5bLdcLZSMi8Aw9BlGeiEhceBeBSEEGvEAUs28Cn7iqmSq+/fJtDc1mPEl/s
JePcLWr5bvuOxdBIb5gxyMMwLdt60twtGxThStdVb5mpMsZKdJYw8B6VNaqf
iVTIefLfWhVJKwsKZJUroG1wxq3F5aHhrWFToQ5iMK3krT1MmYkPrxBOc8rs
MBlfG/wXd3jYgPTdxLenulq5np/zMuPCgjrvnBZ6fxIwHsBpVte4dWGJyJKE
CIYdW5as3vzdgDu6UYmvWr+zpiQ2YkPml//83bhAPG5IZv6WYc9vhl5zylQ9
zK+ytLh9/uuvGYdUTsKnOboguK7q6YsxfiVH8BknDBOPPN7NcvUkRc/3+fQh
apeJ7WOZK7KqGPUjMVt/OzP3RDsrB/FL4fR5Rwrqwq7YrIJoIa/B6282wlZB
bK6pY13K81QnQQdIh5KW9JPueAUvwAgIaNlm6d1/QkR8e15p1lxMnZhIEuZp
xFV1HTvdQOTzNs/bstAq1UEM8K4AfETIV60eI5s2GCiODrDo0k4fCuDNevTD
ttZBDLGZQl2uG1MYpfHe5yvEXYJcJigrSRNYkABs6ItWJXZn+NTpf4jkefMy
HWAXDK+Tu6TRXl/InUi94gfL00vpgT4vvX/6nt6XKa5joGOVxsnCP48dmID4
Zxt9SsNQdltEbSzTle5zPFnA9NkoxBtey3jqzkHJzIar4vV3yKxepGsWz3GK
QUbr9nFZja/ibLId6FdJx1n9zhnGXCSTxvU+k/j5QX6KYWWoyxj9PBKCc4Nh
yNDHfQOWHHp2SxI7XeFVk/bwhMyt26Yoztd0sUXbzz6JTjrt2d+yEAaeOTZv
YUUmNs+RAzdxEDqYP3F7kIcfTul1oZmaIyDGPYSregRUJYt7XnMZOcZb6PpQ
m80OQ/urX0Xwm8pUQnvm65XuCCiuMdv2vD6rJlRGDyEa78mM2IB3bpr4rjEM
l6WiMkPT29YAO7e+J5VoHD8hRt+PRckoWEpcZohQ/4RNQdNZiTrb1yPe++ki
Cdy38p/lH98VszuQfgr2SvdoySHUMhNX+90No8JIyPFyxGzbYT/JvuNPVaOi
k+5P/qmyGMAvSbSJWWrjiiUGAJ9h2tUdBoHqrqDaJMOiwZ2tJzyMHhRR0AAr
lJXJT8cxO8UMkPvIYLrW990WFUzLB2PLdxAifavY7/5N0OGjmvLf9nhzKN7l
ZOYbWX1yS0Vj1xgxY9S7kx7hZ0q6YvWScBXVSin4MiB1h8BiFxZvxPfoTQDH
pOq4f09btO1I2MRq+/x/WTpMXtNgRRXRhaoo1QFL8eCpbvw5e81rwG+XC0nz
uq5s4Ea39xx5RtTqtnpFbbU9vfSxfOj93I/Nq+fRll3gNwK9aKjjDsk+FONr
wJXdbDFcB6JcPe27F3NOq+uKDvC08IVRDly6IsqtdEvrP0q41MYKEleHCOR9
W8s0GGX+RYU08Oj/SNOi/WtS+DEZ2jsJZK12DM9SVLLA5QCfc4XNpAGbWN2o
N3wAk5jxHuo/kWbFDlI3lmkmJyri5N4QpAx0UijA9WGtwU1B6E40kEXUZySJ
sft38l0JlNtcQ2Sqcdp15xXMwDW7fgjGM880rlor0MiGf6a9d2Gj3256hcXn
ZCOH84TYUIFzKP1O69aF6rIfQLhVS6i0/rDQSpk55RJTWw3AtmG6S76kp4OA
TA+tQZNu1cil1YwK+vKwOmM1IbCGYCCWiFDI9FZTNTgy7z5P3bdC4VvmE78b
g55k7jaEaytNc0dan/mdTd7vtnxRcp58lWIHV/ycSsgIpYCQX66rJ/UBQQ1A
GdXf5KoYCnP63ogBOAo/IABWTu14WxrPWObaG8zPof7xfgyLQRmNpL84XUrX
h71tb1Y79U4Z1ik6Tn0OY7XNtm2JFqqSCbYBGItW3+TNrHBBXZZ2+XiKs9sy
nhwX3UmrEny2cJowgRHYXSPksRgALi5Hqwb8eZEDa6jHbYK4irGFrb9MrqhA
CGUfT83hjYye24wAfPJHTg/0wubYINXD8YK3RmxjwMQTGESYdvoFdGFZuEmo
PIPaouDFAOerDkDSrO6He3rheca49qz/GGH4kHvOl+3nZRjvNcpHMBLQg6S4
ShY4n4k+xN4ale8XuYk+0I2qn9fKT8DEmGh2lQW15FVy2MXjU3w+OeAaZrAZ
Gej9WkdcrJJFrU4VrFV4/Pmff51JRX4/AVawEI/vSKlkK/VwhITqqpuLpqDZ
M5enTvwsYE2OryTgxHCsfBU1VtEIFt+s7PVcuWnaL49qYnrvMqQjNJKal/OH
pTXWr4QaC3GsLpOVqwYFv6IFPBxSK2L0K+Y1Vr+m7S3wDiGilyzjukxt9Jrc
soiPcFkIe8bNSoew58Q7qfhtcYAxornaNilTEGqloIsRF8Brn0TgvG96yITU
myGTER3OQU1fpi3S/NlOtleQs1tTiVlxDYp3TO0kW7CK8LaKOFMus4mYUwSJ
kBD8s6mnDao6E7MdrN2qw1iZeJ/CjzO7vUyiB26tKHppiQ0LCSuP4Opyn2Zm
l6WIIUeCkkvDwbBzbHVrkzXUXAd7fAdkK6aOEQeLhM8IkvONnm3KKHpwcAk5
p6s/wqW2OIvtXE3autvFmj4noxE8XUvPbr9BBU5xOlWuOCt5l9HMFgL7lW6p
s6pDb8vyXs6ZBou8bZcWvzo5E7bVDtDf3k0z0QWPy+0mRmh/qZPcUcqt+vxf
QV+tMywjALSWuOrTiPhtqXJju6ULIAaQMscBpbaEBQDeVQI0PRlwwqpbjMPe
o3E9T1QpN32iYmO0/yglyRHqmUsd9RaQuyB1nn3fW0XPEmxvtdiom0Y1MM4f
u1AkYACi1Uhu2y+bQunBedNlyww+Ir5VA+uwsJHbSATRbnNnzFkueaa49g1Z
B9eX7b0W6/CCxCquTXyxwdcOplXqvdf3w9oOu3yqJ4U8Sb3z0CV15c0YFcDO
OSREcE1ebBSE2lkqucemRwc9uKMKwtsiZch+guNXJ+MBLzHsAU3p14JEyQi5
veL1G80xnui4TdHx0cnc0QQC22l9ohViTvNm5LfydkEVGmy4CrrrxOWkD0FO
eQqMGkZjNBXTGxsFTPQu/pk0wvOULahj9JgVIFPu0pLkUEZtzCwqf3eH/Y+K
1zpwUV7yGSI6Wl3Huv49lBYRkLkEssGNehbGJll1yp9pCJ9/sMUT0QEfftkA
ypN1BDc99J8i9K/qv+IFaiV8EMWzokbmmSBw57WU7RDyKf0rkttpLemy0stc
dGWnzxwhGjvvjOQ+RtmKlESQK7Nryl41oDuxg0E3XFc+v+W/rEpvlAR2acIE
LGo3nVxmoEaYAGfHyoyxdfBod/MRoti4oWO8irP1bkzBzufvoUVZE9aXWqhD
N71ezqa6joxtWItCy/Q/eIax49L0x8fzUbwPUaKDqgnjd4/m+/9KlNqBN/TW
7bmthBKEWBiLFv4njU53c8J7VXUF6bc8xrdkvmh2AnKwxWXhFvX3U29IwmYm
vr64ASx5JWPXCbONQJjSMT3Yf49dpVW1EvXlsv65NcEtjThvDffFRxapHlhc
htJdssgxjazKJIGRq8POiTN4t9lG69PNmQK37Cho4gRQiaSG8vHqF8F7iUnC
g3kLqiNeo4SpYespQ4Fe0J+67Yu/bCfXJBX2qhOSac7G32hbjUA4Ah79qVdM
171X2f27fg587YT0Otelk7aQmEymh9BFeBId9kZtcRuc0o2uE2B8pevWeetZ
/FMKstd3zH6SFtYie31adSbxm7uIo8/wyqAX7EOBmV4HCFQAU/ptKvYp0dDY
Wgbg5Fh1gfReMATmbfNVy3ELUyaUPpYVi+bFIoBTPyt6nStcwn/UMEZZLzLC
TQ1jTY7KyXV6Brtp5OgQWEsoJgyrNWQRpKGyCyh/b0S+OqhgDqdeofKuhaLV
LKGdd1/gRwJ91nBdth4q9DnxaYyamSPc3rGcdL1h/b/U1Rsnh9N1ZG213XBU
wd+/3gP4yZnLpKiEHOCXJBXswXOOQA00U6NJWPuvGTTPs+Wch6ThdevU8Kzu
DzGiXjNJ9Ptv1KR4zRpkgWFBfQ9WlD527zmysNax98IBYr4UD94DGos8DJTe
VGJat3yO6qkZfzwf331o+vnLfsI0a086aW4PrM6x6ZQVPs2jTKV13kuuefub
RTOvYK+4RbQeOJ6gg1um7UZesoNpddPDOfEMWz3XWY5iocqlmGksdzwjqWIO
JoMyoNP6Oj6+0n1uS3VbnA6DENaB+YIS8kAMwaGypOaQ9PCuP0VyGsPFDOLo
hLgWOVjzBH6CY6NlLiq6zbgndZwn7iYu5WwpkkBv1n3f5KvVg7pXU+AFfCJR
JdHf3xcx73o0+MXQ8Vororv7fOdfXBip3lmEaHzQC7sYYGjxndJn2kpl2F80
KglvAbYVcQF3Wtdw/zymkV8Da2mWMxtBepFSfwe8mStPhOQCaPDuc/+N/SPh
j5TOiRDdoyBmAGKDury1JuzkqFHztxG6u7SC3GnDSfDT0fuHyLepDVLlAWDH
KfBGYd3kfbHg4IPvOgKk3OZ4MJb2+5WZ0aeILeEmnUqQgsrJntXP7RxnnsUk
vj+CGDLEzou5tsmsb0zc5OvDj/KYGLDYYZrKDZgO/H7NX/1CeMRhRYjpHzg/
sIpRta50GPUmlGxEfxreO+Kc25H+wh65F20Ph8AywjcWKg7Hky/1NZmrGkqG
YVkNCY0fdChKP0fzgFt/AOfDcQkvIYapquL5jUihPg3Q+rNjRCwbxCNYXzk2
9fDGMzowdZVIYXiPx7GeD8Vp7hZOg40iUmlViyIYEJy2oSco5jsbEM8yBb+U
PrkMBbBuUHSidsQB8FTfwzi+CwSLVqPMHlAQ71tFe5rOew9Fev0EIgglzOiX
kbW6LSg7vydeH1yc3EZyCRxRDF1c+lfR+ID7Vapf0WErXIytsU8Se1at0k6R
PGPlekCeziziF4oEn4t83ue/zl4XfcCE3VKU3lEVMO/uC5Z6UOszMXFLV5AA
9O8CjpBsmgu3PwV8tnGm74pl1f5eA2RUOymDp0gPbxyPPX2LqODXco25Tvoq
aUm9N4iKzxK4k4luUJp9Aa/k0gXCo+UOCOQU0Fp4oKHahi+k2D6bsBmkxEnE
jJv4/Ff7/gyXGjwKu9FAu9btOSicoccUZLEph9YHZ5ZBrYHTozGTc11XlxIS
KE0pN7vyCOz0cxnK3tT/5/3+6fifT/rF5pGn1kfXAL13XMZ6tcucD+HYsAhn
mkndHWDNILoT0or5sbve3rCYJ37sAlQ3dr6XY1YyZz9NdbK8CfGU5Z/eMofC
2UBo2IGK3ScmAnzGsey3gViYoei6Y0t0FgXlZI6xTMwO026rrXyDBKxGJaHr
W3NpjyTZQVlmI8QkfjcZp3peuK4T4to1dj5T6TZIJSU4kuHGD9E0uINPl7Jl
UBTQC+TyFXRXxRDO7otRBURvwnMiHbsj1aQhMU9qGQ7vFd6C7Digufe5X3R5
FV5j3BabcS9vDw1WOT0rhzhapEsNarVsdEcFGMl4eL8qB1xSlG+y9gB1eRGg
Jsht5mF5sC4yLY2qe/gOJBL2RBwGMXZNBxVaf9lBSXpzkFAhHF2yHjbMjMwf
RvGWit4mV+XIa0pcWlJeQ9b+o6xb36TIrkyciLwzsnFAsIn1fkCxYdDmMzEM
0M3GUWJAYO6kDP1ChAx6wfTll5S9Zp77Sj9iGHqseS4WyosS8uFd0of7gjg3
esphVr5mZ4fpa9CyaOqeVYxwaYBnAK/PcjS2RMc7hYhEx1MJl35WYQCwYf79
ELomAuub2wJlInFYUejX7mxVnViPjyTiqEpv+jQVtiYBscYqNOC9RuxWm8qH
iPeAN8rpSNF0klALhnPvFMz5tJR5Sw5ptBD68p5ITVMxJAXD0Yv9U4a4tk+2
qNBvG+eLvobzs8gj8eB5kVC+ayaqXynCgBpkn05aUye//PM2BqKGMp9Mtfow
Oup4nh+iRCYXsh0nP2RZ1HpwY8rfoM5r4tVBAuMOXJkCfsuL5BaJ9vqciLu5
S6wfJEyALKWMfUjyVHjn9No7tc4Cd8diQodlodLUppEG8s1OfwV8KV37mkgs
Q9YgdI9sx2bnVuLxAqMEHe/ygIKckpIx5HxneHM94RrnHIwvj1kY4rIjua2m
wsMgi2KJlOMS7ZdGM0YEXo5mNaI91ex1D6Xh/S+GozrBqxdtuHjElwC3KRxP
NMqSzQpCIqojcky9g40ut0ghaThRCH+hHnU7Uv59ahBQWdmJEhbsHVUnJtLb
7YdXiYtOXwBXZZ+D7KsNVieJFB6/vEyhldOA6ap6w/TNF0IHjTsJMaJx86V0
LuOF/2ot1n4PIyHxIBDL5psSSFbJsv5BKICWlQDokrhvQlr0ZKuGOS9VWs7x
u8bGvR4LxO2qIHvJl3+dhMZegHQhGaDDAlIosp33vI46O3oJMAwjEJod25EY
nSIrRSkL/1BCZRcdaChDKX/NA/dc86fjbNs/GlBAWRlowbsXgatDbhTcUwDU
A5/B5ioDPj8LoNQoekAkuU4mhHH2JCgb/If6EdZc9LtCWxkhp60MzAH2vw47
H8YVC/B9IhP7PGju2t/33xA+F3+/yleECQSlqEhjMnKkgkX40sabm3dp3Rhn
bjBxRbBMd5AhBBNvVywHqj6nxL9UWK6j7vWmbNAWCJuu9gquaRZN++AKPXMp
Z/8AP/Y4/gClwkmuu0LwrGuZXtPxLLlQXB9Yb7doAEkhIaah2e33tbmDT8aJ
5HXyi1gmSfQ0lb+G502BUCkUG9OMO/7I/8OFUZoJrMlAioodxhQdbnaBzj1A
IjR9A3TNRvRhKNHVhcpVZO1RzlWQ46LAfLYvOCl6M9gO+7lp3/Q2bZftptS5
DBzZLXn14DLTJmBzZhby745533xscv36H9PqUjC0SfNlgUeWQIl/oOvYwHqy
9zHPVbiZ2qaWf8ZxSCaVn5To5+AV0+ktUbzGUpYv54IufsQmGNfnbOW+QJVH
6YIbyfMYxjhjHNc5IYU21yR/kpJ8Tcf/if2o8lkdr5cN/+UQAqancFV7Tksp
bODye0oiQgZl1F4jFUgGNwE2r2z+gqO6E5fwBsCsGEknjgnb2HaAsznmMRyg
6g9EKYM3vQ4eVrg2+V3+fahH8Vtj6a7kyt3du8UFd/p0Y8UJlJ3Mj9dGgnxR
L5rVbgY/OIwyp0cf8bNExIsDw/AOK6lICxUsEiur5HZ5Y6o7ua/YB7ugQhZp
iiWUCtduBEHnMYTyW0kd1Ei2nSCGuuZGYI2+1A95CBNxpeqQ30VB16uwsc25
VNPhPlRXFdDHKYU6pc9C8N52KZTrkVSp0KL3FOf9F1bmVth23BMXfWN2B+M9
U3a2K1zSNQy0ZH1XQnh7/Pl2y9hs7EIs9e8maB8VH1fO0mSlKeaoQvrZchBZ
Fx17pZj48/z/VMt2Uz4TjGMCODmK6vLqjCMLS3PhWziM0Cg/IqyohJwl6wPA
Be4cW5kGOQH1QJX6CaOgyKq6VFXv5x33I/hAIsYY9bih4RJJKDHhSeYsnoH7
xIX7mb5xw5jvrpuZX8Oe6OcI3Kp1m7uqTUVag4eh3m6FU0Ue1+w763lW5MC3
ddPMhmXVc6W1AXacdt3e/ptR9nkNXBQ47CvFCZD8GAQlk+HvJvUEo03Da/Ic
odF9pqQXKVw4cR2gTUl3I26u3YesIidzIz57/el9+pMFizVoHSsO9SYZ3kd0
uSjIjNMyONaWCDeHtt89PaI4jhdK6hWQHtyfCFl3+8TYx6Y0iMu0Xk4eKK3/
P7VyJa6e31Pqv2okMImYozC4ltRhWGTLsMi1scBrKGZtuA297b+gGzDYNAhJ
ggwfWcZ720t/emYr2iyUhm648oiSOfXeW1/4y2x4mxzZLct09yRQDzXO9Uu2
QssrT8jgA3XamNdJfExzHgpU1jBtQE/duqUv7yNXDDDWJLyswkTacWFzXWcq
inPylA9Cqixg1OO/q1sed6RUXwmrzxBh5fDunzjc+OiejEPTwC4mlRI5dUMs
MWWA0hAQXpD6/sTIgpO8IcvRTUsiW3b69+3mk1XNlFtlR8V+UUxjZsG5w+Nx
UyDDrMZIShhcO0ZAHJA3vXUr281arfars59/T4zsuY1c897RHNIo32M4llKu
cjHntKtnwCwS4qkvXEXBgJbcSy2HJVSHd3DaEkG887bjbyJAh/VoB0Bz3YJV
KCsHCRv/WrB0N3sDwh64Yx+QktvgKk4YfyZaU9cPwRO1nxzpPlLUaPWWK0v+
jVg3PANPj+SoX6IgBPTsxhEIDzOYoiE5/W6yoX9xZcsY1l1ZCZ+NZFHMdoje
0pyK0gzt8COFJ2lWCdtpg7/WG6B3KU8ZgnsPV/xn04h3taxMX5XeGrHQw06f
1pWWUoWy33fJHSnKvJt47v/KLt1nRMENrQwZ/c3rqUKv0cKFwj53ii2AApjl
zAnX6ELVikWLskxuYdvKC2VdbkCHledzSThaxf/pG8yFdUaao8Uap1nX0JD+
bNE+Tm6Oui7XzFP8K7AxZQd/KjrOEbTd0NvvZT0Avml6Xe+m1UzJ4HCU+IX7
2O7dI8Wxns+znYsY83kYFkLd9nLkHEkzT7ULF3iMnrLj6lSlmtGIXkz3CB2Q
DwPHW9kaKofG0s276m6aalEQnUHbzpyHW0pFK00/Bb1teM23KNZoStPEKFK7
qzDRW/mXHYE2fxa3P1ls2JwwGeIgDQAeA7Mc47yYQYXu/yssDaX9zLSLznE1
3eqpQL6pmnGhv8vqVPJmhvmI267LIagab2QPSd/frIwKKV+Jn6uM2uiZJwXy
/PW6hsh48mNqgs6agtglDLDIntjKRPOG8l0M7FU6FkxgzI3Bd7B1Nob43qwE
K5+V9z7Sn2dcp2afqeDLKO4Vvo4Ic6Nz9Fg1+pQcx4ueW92U8J/169ojt+6P
Zt4b8iN/aXWrPsETw+Jj6ofOSovwX5DkuymWHKRta6NfQ1ZuxlHS44IlRm+b
3Frp+cqv4S7x/pCyIcZLhdc71SMqVSrwpKpuSgLqJjZU205UzzyGygByYLP+
4xf2d2A6lefAQ18q1Oaxea55LN5XbN39cWRye9N/flLf4cnNapPMywGEak1A
5B+qGWHru83RhOQPwXynOATbAnXzWq6UolYMg1GauYFvlOV7342QZWX/AWTy
gHBOND5zvK3MWq32g/sHfXfj2scPNnddlBCOBEjSN2fbymxETpPQYZPM2GAj
RbwCglTi8TAok1GBbd2yeCCuVhnD/f8vr9q0radQHDE0b8EJI2yNhEolqzbR
4Zg6q4PdH9vdBIUAvxeQk9essVeQFz8xKndrpAYzP4TvyRZHOkk0Y+pwawui
hMu5BV01DZCvIMv9qbIc/BEAWW+wMFjAc4svpp0jc722bNyoLNbBb8opJMS0
1E6fDkGx9/DiXRN/KWNPHKHFL2YKSeb03oCadgOpwEfUgF3W/hCnugyzBb0t
xdS4uq+zOS0LEo4wW5a5kSeWYzMnL1wTjzXYxK/2+XsrJSeIADBSpYebUBrk
qwedcEeA3YYUSrTcVttKl5vC2I6rnnCkOG7+Gryq119mif1NGzIvBZgneUjN
DDrH50VmX5w0fuxVJ+h3KyWrLfs21U1ycBHoB7ukNKZvn2RW0NIKHsieAOFZ
lS64O/CwjH+cNo1tPEMazqxP/7F9yEZN0VPDhApaJIHhApHBVxpJNc/1disJ
mNJTNazrbXr7WThXj2xhUR6y6sDhoO+nc5ZDevQAve1CB0YE1cVFIP7W7qf8
yZ+S2BYQtxO3XmaAa9Az+K3BZZmXtwERW891OD6m1hHLuRXf45F11J21rkpA
I+l0XGaNya+V65mqAU94ZPqzteid12QIpicdCS75szUrqFhRZ+JZ0jirqYyF
2NynzfHKpm2ZjVPGNZYCV9+miQRTS2BvJ/WaUap2rP2R06OyYmO2ZUUOJ1iI
hkGlMNo8QNNUZVqbjgjw7xZKPrMxq91WOm5O2ZKLIht29HEXwNEewTY5h1DV
2HF28mUPT8JnylkYRYAJ1oRbjZRX4qa3t8wAmwnO4wvM5b3U1SyMxJG4dovP
J4oiXDAHiTSEBtMwrmv32RPyKR5EN1DtDQA4hZF5jioph9rj3ZdDnMrFBPSW
mKZnDuQaGejC/EH/QmSWiYvoMcO6YYNH5o/BF/kIcBclzdNiAg1i9p7W+Gvy
gP3Z+qTO7AgonKpGc/TMkW4cTfMZFCp/bGF8+DyJlwUSj4K6+s82IiIfCAzr
mVtm1cHktHsGgPEahBX26FB/4p7WoOqSOlXNx5RDK5Jmehr9mdKWRU7GJ/YL
tg1uEQFea25vG7p9qx9HWbm2Qx6KOR6rpFwHT89rr9I7aeJ876S+MKYy7bA3
1xjeE/PcEAUPvUzICYk6Y3oC3jL1qLZhxQDFssklU+Dj9kdFI7c2t7LCNfZw
c5BogVVnW4s4tmLQiJtRfjVe68w/KhLWENtx+/W5OPB5Zqxr10euHnSzqJan
9KnQr1QmcKIFuhYVJ/Alp2z+tsRHec6B+ytwDAi8hKvb98R12v1yaN7DU136
Nf269XIB+TnbQRp5Fuj5lPrNY0hTSeroO+KCcqSLJhXuZafecPfe1aWbaEjS
fb0RIkcihf3TJZcJKTmbmkukgwUxrValZLZUVEJLByrc1SaHZfsk51Qp3RzE
PnUJtXh5GKyTI6lfuo9gCtnlCvd23fW8CufuupktM1PfXbUNIRIvB1YrVtT6
lgOLIJUQeIJcba8lTP66KiJNYyPWeiieziuSr/bp6WW3ysmguYsKSf1kaTTO
0foFnKhQdn01sqpED0VTZH27/qU8T60xVoGNNbeqwAkj85RVxdmwVLahni8C
8ryKS/Nt0PhzFPGA0s5heFfm51YSl4sgk2Qw5rWmBT3BjwCvwd7H/kg9qril
1OeRNHLd82bIR5K4rnX6xEcVqHtDn472/F5q56rReqHXtm0PuYUDnuHrSOUN
zoc2NzjhI7bX5G2oGv/rKkm0uN9YmbMZE8bvyuTobA5hYpck/Mzm7zLkms0T
kAJRgtQr1Bx/D2iBs8ZodQR5NM573yXdFG94EmEgryMEG7+KkZqGSMe9h4vP
XVt8hiMMoeNVwGn3e3l1QpMa/GSgAdLskMW0jKu365gUrLSYZTT6vAJlfD2d
DIXaumPUSEEZEZQe94yinXyej/EG2Plz18Y6vBT0aPz0XN6tEUHBbSn574bh
ThpEI77jaR8toKZWRJ7IdDr4ZxAMmQcKEw4CZv9kvaY5BtzK+rE0YWtZ4s+p
cPWRkqA1FjQYb4SDy1cqNtYPRORZlbZtq8qX5mXl0gF0y5cxNLi55VETbl7S
Cp7K14gZ7jGpbMUkDZxdKU1nPi0ZFn7dcc8Pk5x9Axta/afeAocvCJOpSnxp
kp14yk4tZGUOCPbnPT3jEL2xKQBS/ejM6zfY1vuldlzzjQNyRGeQj0oLtlzL
ew2L28l0t2BMWncelcNeSo9IuaW+Q2L9eulB6mT/vLyb7k4MMerfdaD2VvUb
9T9oCKre629Zeq8OKUY3xv84tKIpBKndNVgjGju/DauTBHjjk6d2YxbfmuGz
bTEmiwscPBP1oQ1iKNwy7Kbh4UbiQ9pBEJMvJC/tPpM4XuRz7SecK8hHo3Wn
Y/TTbPHIki5u/VCSV8EGf2jxbIlvqKZ2FQoqoJcUPne6n8ICBbWRlK9DNrP8
z+thTBxvP2HQ+TQdMbCwXVs562D58I+fNgXbGgixjXj/xr08e9ortp6noqc4
KLEY+qJ0t7VM0cl+G54oyIA5wh5uAJRdOzcbW/SuFM/wTnuhIyYWqmdP6Xgi
trHYOv4yj5VQZd/uqq8zyngYMfIfX40jjivbglZKu5VSszT0QdPqdXe6Szfb
5MEsuGORpxHEvVuVRvatEgePWAyafBEADKfqMsQLpVOBtmKIJbgj1x0xnZST
UhGnTwW4jFVVuULHA+ecVS8lzHOTkBkoG+dzyhkI1O68C5XrgSYFMq/dNWkI
hewGmjUs/0BPQ4fjXOS85Addx/twx0IjfxwW0FymSfvjORzwBL3s07rHyT37
rBSWRk3ttw+zV6kGXkkh5Ka0ZySuzx3ZtYcnLzKeRutcwov3gMbva7Pqn2Zz
oKETN1sm7WzZ7UI7KH8+JdX+aOZYBokPE1+I0HLvOA2bX/D/kJJa1wDY7wBD
izoAhx6mCNEQGojgkRB1IdcrfrHsnfi1aK5TynfE17+Wq8hcPm8GlvdkPZta
YcvK1xhe/TnU9RrP1ZBvnKlF/RQQ9zDe7SR0FIq7va1lsaRg0pYWgxJzELRx
ezcoBT62DiHEx8lztC7rG3vwXseJpHZzDm0EjZR3mhaYg4V3hUc02G6NajfT
g1xyL6KO4h6axFYNM82/G8Uq30gO5QJhF7E8B2LVXgwB79IM4UA5gU5GdREG
lc2BgYPR8ZLkgjDoVMAUfn9KDvwnOLK+y8AVNatVFc0msbHQt7svAJFMMCTR
aeVfx/INzcFBxvpUg2rCM6WIzqXdebqG+MCUKyMpwowyZbjswTJDfzbnW9fQ
T54q3FazbVvIhm0RlBZ37nTLfBRjrO+Bc8Jswst+B2v54HRFHw690UA1bbdu
G0jRmj5Dp5GyrPG0m813K9U0eODGV5GffKjNbOPtOpcJCtmlHSPTNL2iA4Tx
Ocur8kI9EDRJdTihA5fqnbX6TGG5itr3a7m9NQ78Fn1uDirTg+nokTiMtXhm
aPKI+DpJjai8d+qKt+WfxHnrwmHkyAJjT9mgbR7Q3cXximlHCqnorD06BZuC
/lAF83vwU+4F4qpiBUA04Oqdj1K1qRR8l/xqm3GDw+oS2jTGY4cWXQB+nu3d
9gt3cOfReZrRVDUhz7zOhUrRiA9t4l8ofMANWTQfbHX7y5wG+k6s+0VsMfD4
iZ5A6+SuzPAHhTUpN8U4RqSnPNyCfQETVCOoDGSFZCDe0i1adWQsxhMmdrmb
yBSWxf94Br605eh9LHikkeVvT+3DQFeov2mlJXf5qjkbE4W24M0ba5ckAHzm
H0Gv0AQl9ryW+FKX6VA4Xv8OeX064uLRnfyjhUCZQoKo1bZVbzvGb6KEjtpI
KhmfXIsi5XoSDV+f1TnUw3pT8cWjovoCoHYlpJlIgRQsz0wCtC3k661gphHu
N1SNKPa1LMS49xLT17BplYBzwrFuvZxKA9EujjzzDu49iHy53NYgBHHAWJJP
6HjK2fTJCJiQkxZdnnQ6LeJfGurMTvuq1U+COCr9rGnJhMvkKp8qqdnK/SOe
w+iitO1/MKu5Rb3Z6F4oBVO3vMxZyaqPUxJsO4tvzqhrA6GdWwsOXIRNt1kc
ICHKR8YA/o++Kw6AnjGDu2ZseyQKYeQs45zqPwOXIhX6JTWJ6NIvhmSbkLS3
xre78PmHqolra3dHiFAH8oSeklYgxXJW7fvpbPgN4cI0ibqbQlyJmFmqz7qX
UMSKVIQfAacjJ6qzzSfJSgJ/gHuZRJAo4OkKXkC3WGCOj1D/JzoE55twttLD
FgyPkcBasU3mNt51Kamp9tDcldeSVWgUsecky/PW4BqtslaSOzM9YD5+WU1Y
HtES9/nRjdKswYTLqMgfkabiBpbrjEAGaAY3DNjPsqFsVh+i47pRV3vYeYpx
hiH1/NpwWa+nS/Y71PGFS240I8OjbTtlI5j6NMnJz8stCfv1MJGAGIbHD5Lv
qlGNBfjV0gnDYNjcXXNchlGEB7L656F2p41dLCbmRJqjLKx3oj/KrLqSeYBl
AuUChlmQ9EogYVmFo+s9ABaOu0JxAndHwLGiQ5f99V2YwtvRZULKDGE9/BHB
6LhPfwMRR8a3SuDpYCRLHMFG1h+5LkwiJVN4H3Ldl2OtAaH57RYvlppludUB
si+jd/FKsUQgpo5eHm8BihXX1xLTmIFBJEw3K50pmGkQcynnaZu4GktmTT/y
0RwutoMeftlXkbS01fd1j+T+Nbpd6ovgratlIlN/OY+Oxk8LSYorFxY7e8zk
OHEV1Q8xPDpGbyfTzmtaCqfCqzwvSQYwLP4R83i5ew0TdocAVoWpdk38U+Y7
252pDybKPRrLw7QLMkvSOqg11UvRH2kY/q6wdumHsaHhMyyz7o1csShGAry7
FXXQbQKwEDRpjz816Io7stTqlRFhrCtV/NpStRmNkom0yGwoTHaYnHMqHX3+
iIvCeSc21tlGyhwaGog2UrAuBDLPWe+dnhg+kGXuw+Y/3pc2iVfT1LAQPvM7
z/Z/dc+aKGAHAlwe28qmbtkW+/WvxPXEiMVAVtG501wtH0N26xUfm5jQ8fCG
bRuZXEj+TdmwpAALZCNzodAZzNNYnGLLJWzzdvD73T4U5wHyKFifgUH++Bpl
lLJxypomoMuV5DsW0sbMprQPhsUXlrpRbmOyaaAFcq55+UKW6nbY+zOOlQCZ
SDpk4GyGqym14+FeZOcm6p5GZN5cZ8gV0TDtxrCcb8jvqbhhT3CYBhdHoVZN
EAFmCL8l1ryKrhret5NyQm18fA7UjRWGBhcamNbBunKodo6af0jT4VhBIatx
Rzgh60av20k8r53a+onin05yVc2Qx+CQevd5Gzyxg+NFbWqfoNKj5jcr7tiE
VAmXi8yhVkfCo6tLRR8obPoAK2tPoTapUvIMmZhxAzgnHZ386yDdWbmePEeZ
ssb2tB1WuMzrZV8N7DdaN5oiS30682rmtpDRPgLJ9E7vlJ0HQH33cbSoVWXZ
pMBCu1yWe5WdgUGUHzTEISDmfhUc2JQrEOIOMQ0w02kZgmSw+1NBV18w0Axb
dgKqfPHb9a6yXk5ZxXmAOsXDf97FWFQFfl3hdMUyii48cgQhWc9r3s7oihjE
LX5WAYTsQHKs1MWvMvhdpfvdmTp0fsmG6/Kuu0pzAy7jKJbLBS3//5cUByRD
y7VgBDSHMNdPuPAQ6QPpQKlgf8Whe/D9OFVAYFTBZ/fUpGTwDsDlE+HvIEpo
v8mS9/aLwdq8+BqCdktJXbj86///tzSCLZtVuTyn7DbhF/MxQyXIld4aHDps
td/66PjL8AMtXLewIbYttgVqljqlrwrp5lTD3TYMVz7j9Ez4Ci1KW9v3LYlN
8wsf+cPJJNSnhRC1JiNDAM2d0CJ0qmomukSFZR5SVf3rpaxSRWRir7kF8kDl
iE66Ts9kVZeCt3njWAHsFzJHqklaspQ6RTtvCswsBIfvu2posohF5EdQ3v37
Wq8+N0jykbCHgz6AZuYqrM2dBts0dWX6XjweBGliTB3PrNs7RZBv+ILHp4BG
NfBXCvY6JsbWuLjDFWHjjiy4pUTUXlgk1dTN2wK8ChXy5yODMXienx7W1Ik6
RQHOz40C0sLW5vx3S32TJuyBcu2ZhcYXUBm9h7PghVnckNNH5shTVt/vmdAG
cslFdK3tkFdtg4M+EXEz0e8Pw2UgSAEw8JAVrJkECWQNxfIy50I6C/u88T3z
+xSSSX3M9fW7L8R+vfxi71U710twO2O7NnaHg0k1/83Az3+dkTO5YAfRIcNM
1bUEUoetYSSunZkn6HimpBV1b010cgK09+8ElJgmzYIWePf/Tt/3EepnrCrO
roNUjKgtTHqh4OT9xhIiaQVTBwvP0kwxNNDxsQv90fTGzx62V/uUaJCZTLC+
gLaYJxSX4mrbejSNwEK0FVJgbluNE/oDrRUqC6szqu2TCwVALq64d9lHv6OZ
fcEu+haeaK1tYDw4QF6hRpUDZf7FTAP4N8d/QxKW160JRezA8iZj10YBrYuQ
Q4D635K+VSu80B4/3dw8sz9fOOl1EdQfCNVn/rPUWzqDBa2t4EN/TQ0ONqxp
F74/azcSwBKRzHj62g4HKM+DxGSPR0RlxBsLE0+UQcK0lC7BZ/xLxPnXs4nZ
X7BYOAKIRyKGoDldKbEZ/2tfuIwUZJlWRY0eC3G7SIJMo1MORYhMbbXNOwIA
JhBlH7lWHwrNRfSLZ5lBP9NbPQBKkB4AbsGv6vrke8FSkXsJqOHcf/OhG4tO
2ex64TORmuImcO2XYDq7LeR8ijoyqAUo05+/E5cmgdUdEFevszFAGVrODFPB
QAtPF1MBk4/SPWK9orchlDV0gLUGwSogLQ1jgngYb0udy9oIdoGFOZHUqPKF
r2+C6Azk+FMB83gWPkyaKbJSJLYr7Yl9Z4tETkyKYQXkR4vqsI06BBu05pXV
Y2xjIEe/v6OIwQy+5eVeVrCpcqYvEj9wboH4/lMtSWFXFh8X3AbBKfnBaJlE
sUNP1KpTnaaRdt06ScY4/3CuFIbDwK+yHQdAzsJ197fkm+8Ly3C/v/G/h/ag
Tnia6ERlnF0LcVaehEx2+RqUqXD2nxIE1t7t+Zl5pwWb69EI5gH9wvwBhQJg
CxWMIcr68+xjMGEzu11KuwQtaU3xJy5dVUTf1YaFLt0XSR7UjhGT5fun/2jW
9d+WtcNv5c7SeMR4Me74+RrOha1oG1Lt5qU2U3+KTQF4YepLMFbnKHk5yM79
ibGByS5d7HGo/jM7XUFeAgjR4bEpDnKbxztsjTuA9xRYwsZgaktbTkq7Dzkx
WEhJ6fGFisK8wcfpuUuhI+tejCQ3hk4/XQ0tosRGMd5VVdITPRZKhTzCxjIl
sbzMBVn9xHawKqRmnKKnFX79b3bNQCYhfbuXmhdWA7V6bO+5JoSUI5yeJpg1
v3CqtHJykT9JpCUXY/K3P2EbjYVcE4lPirK0KMcuwqEkzvMOx/3MdZxwr6FZ
1mDXiTEQaDiW2wiT/UHxXViooZDKPqDLkTqUFRSiI9fyGqChEvLcWmIOLOfI
HKxYyXJfKa5Pye2N8K+N0J7bka0RnUZ0OpGs+GtIscRU0HnN9sbTmbEs0Ghd
uF8QjyrjuhGT5GAao2Fvpo7BrnQR7EuIzHPWAeL/jY7uHbppFSSHLqnVuauz
bOdbxnwkan9eoumazXqsoWLXrdvVIahZ81CrVAj0elYiVgb+iPjrmYUtVHMZ
XLB4Hpn0HyRsBw6Qzhy0pon1LpOZrJbJS1C76VoSUsPFnH4LxeuNZls0y9Ox
f2DLhtCsxttTFgYmRYIufFt8f1qmsu2azUsUttcx2Vp3GKpbPWN02Xl7nblA
jMVYnR53ehiGpu/eUZxsLvbeJZJdV0KRiu4SOmneJtdIs+thHDXx+s+kQa5A
nJPMJrCv6mn/jHJ4gDemRu8MLvR71HYw9ZApmVKGYsX/BECJFU/cEKAjfwwr
Yy4xjg5rsdG9UQPsFMfYV60IVNiI9ug8pJssufuB1IaVYziE0Bbu4HR4ZCEm
11t+iBfqg/t//CucMg3F0E2nC8V10LtWVeKYdm35VgGR5J/tAXlIaxDCJEEm
9QskgM2nEotlIX9r/TDEtHaPVbNk68OZd1mEOcn6kNbA6BxofdJFxuvpRdRs
93l5BjaFdHva6ZQqwbgD6MfIGeHPkL5KIKTuEt/j5L5aDzzL9ELX5Es+yzlh
bx9iv5ubmNwwdEAsruNydTaBruERBaJUgH9IMT74euVw5nkVPAUr1S3ifRIL
TDUHSMgVPuS0upMpKvc2T8rLbf+YtLqcGwusaprq2uTG7Cvc7vLz04cBkXAj
+ybYbqnkwv4MMFd4iOnflNnFqpTuEM42Ay2+2LFZBZ1tE/MpWrsR4NIJKJAa
KBwqPfheWdDLRqatekiJiP7Hfn+OauH/nZ58ujMzcYaLlEiEfz1m6mIzBGK1
rUO8JvrTyFSn0WcSGeP9Nfxa4zaBsvwBoMLTHUf+22FL5FWu0q/VCA07NIiL
Kijv/Nmt8aicOHIINB8D7At5ZGuJa3P6lkxUcyf4Bpu0Dn2TVQXimZqdwRUY
NWnUtBsf6mCgDw7uW96SUuqdlgiiMFzt5KDRAgaSOSG0pOCgUrRwxGgcTA4G
YOChym1NgTc3qMu/2/Vi7MBlks7ihCXzuMh55fHF9Bj7eTGzZu7604+gleSD
RZoidctzNbsf3q6NbkgBoP8aMsCNQygkVidmXIrUetxNarKE9y1NSX1akqRJ
IsfQyXRUwSfATdYpyb84izQTwg7CHnsefOzIgUNkTIfmrymX4C2Is0JmdGcV
sHZQJbr7V8P0+k6K54bjhcbXxAyoKHszBHaGcchUlqZL1nMowkE/1jacsQhd
+IcVfyr2yXTKgnUGXkBD7/zV+DRr8XfKE38zIb4dJgU8IV9Bt6YAW7u+Kv7Q
WvAISQ0itkdxJgffHR91m5M8bFuO9+8TWe4g7E9wczrVoP3RA1LboTl+PaHN
77oZq/iPmTtSOcdDutETmeif1dEDyRLa40HXaq98q11+KyXX1RDpnqvYzy1e
MJcOd435fu4K4Fs2asGsYX9BEkK3Pgc/x0pASrP222FuxKBMzqifwUuERoGd
N3Rz47JMwORUPLJILS96A67EbJtvEpXTy6ywnmExZk+7Q4V5pZBfmSa+r3nY
zBnjAg+z614ewxB5Z6yL1eQgs2B6U8udwuSwTPUStrL4Q0medRBOe/CEWzRy
cdOyRkxp/PIoZnwLvxam2sToe24IrwXK63NrHWy8/t8lirLmAbeGAGr4Apzg
zI5I7ShbxlQJEo+zUaFAuFgufIg1XOqJ0gTjrwk6cHx/HUKuhwe2+s0XUCYG
OZ3ewAlA149rJThPxR8sa0FpaeyElf0Lh5t7mGQ8vJNOaXMu9FJQ0s/n76W8
iJpMrcv09wy7lTnqy8uGLbfBoKPdx360gz5QC7mUpqM2afKqAbWFsU/0hXaV
N3BuWabyZQyEbl2QXeTuRyNalDgalwuVq+2Qt507eWXWMaN+A3/cpIeKGXNs
G17stR1gaMmrAqxYN7ECSaxKjFFNQ7xcx4ptpBl9U1mNqd2gtPfTikcGsZmk
ypk/hx8ViImP16PU9zPfdh7bz79xPUjHUs6RkEvQyeDXmAzz+sAnJ8nF9YER
t9Vu9wiCJZbVnuAtPTnmDK96ABE58nmfGZSZtwtSk27+mBV3ZaOubxmCsQRv
GTqOIjkMwWw1b6fkK4aN8qNAX4aeWOFZV+XMxgpDIJtDtMKxXRJirA5fWyo1
hIwOVPdsUUJ9ivccstnWe4ZHYmkeyYRDo4oFTdxy3wyUu/h6qmW/UqBhRjxa
SJzMl9fBxhf7UKjkgSCCaSe/ff31+NrNvdp7hm+AhUcSx8mfrfN08m221Ktl
lGuVMaLaZm+/DMKxrG/qFIBDz9HGV2GH/OmKx7KmaTaS0rj5HUacGxiDi6H3
9mvL/UdCZogWlRvX3HB9vb0X47WL2Qu2jC4mJAvsB8li4ql3pM5Lw6qXhwFg
yESBdGcE95t9d8AJTHmoEQvuHMe1GonUcbEvJ4n+SB3uSqHX505QwppupePA
jAxYMwS7slRepXgsFkN8ha4yxHStgpn+Hm5OSb4udyO3nt7BJrBJukV3Y5mk
SEVG1aejSKlcsxXdE6QQP62IdYFmWWEm1c0gS8kjMp5fUHjg3yyCk+Ikab8G
/L/AJMiENvqnfAdi3AYhELu02X+Wmir4hD4y/NAS22lZNjNDC3QKABHbS5q+
281/I2m/ss24uJVWS43fU+04sw+8jTQfN1J4HpQpPFXNpFRoIVWPIv/H3vHT
20kAdfkDGmNSEKSSXiz3H7dhxHjnDbtMovtHLn3X1sIeSHu4KSkuwA8ny4q/
LiB/mqI01qk5ciZUIsfAzVUhffceg8uHOQxgsR2rkloxDgLFJGBMmdAtMyci
n7WlKWPRItHFAxg72iYVg1DfRXT2U+wwFnx4Ux2DS40ySg7VYdmyGWbD3A+H
Njz4VxcxlSgMs2LkuVGMqFaB5IRXSclsDSnVfpvz/OqD4nXOtly4rlZR1Zo7
+pd00GZJluYnXdKc7We0J/otdz/2vSxy7Xn8vDD/LxFQlmhxtVDxvkj/w/vZ
CHQzLx8Ou3XZ64QeaChcdWv8gD8PO76J5psB9uf/+ub+pcvMt0H/Utm01baS
Xv6TxFkitTIcrOnbtSuqTOwfFljs4TN8qgI1iXspyDxJdQ3L5iWZAahKiqCC
PMARYqKzf8BeF54zOjDKCQT2cyVnJSdMAbjuzmtiIoJzD69mt3nCZ2ihA1L5
dTBDhDrDxxlpRWt0l846aCYZFxjcTf7oeHNza+mKIYBQibv3m2sSF89eDLDp
LpqbtjVPmy3YJ2WFpHEFASK6scKzGQiIuLbyqdVO2RYCOxb/RdSe9gGONdPD
xGqrGiLe1u+QqA/U9rfo9e4uluEdLWXv+uvs3ZsbNC2GuV7cMSaLIgxXh+n+
out9Ze/jH+x1qFcc+ggselmPD/1/RLhYTUwf/FDWsqo7V4IK0dQ/MWe17aIJ
3X5AhiVhOaiNzba8ijH9pjXxi1jq/SJ3dD/FTdrJtgbOHdiYk35VV2pVf3vM
yFxSUr8ICklgwtnbbjip5ZdHOFibvmrEsvmFQB2SISqhOlhf2sCUaeD0Kkni
qe84im90Q9aFMp75ySFY4KT6pvxbB906/n4amdqTBRwJo5p7zJAqCj8l4Hu2
eMAVloSoePK2md0iBfLNljgrWOFXlJYCKtFRANJYucmG8GkMGdIx78D67Zep
2LJl+wJkRI5ui1OGJkTCqnHOUC5qLGyTwoltsAIQ0uOgqQW8qUk9Gsi9YNO6
1yq0IkMuPJzHLnbt02Ej8ITnyyBnZkSF14WUIAzA1iIZC91SpdZFK2Hpmuu8
YggpnSQlCgmz9PVl0zS+bfVlPzjPnhoKmHmqYaQLUQjG+MwHcJ9e8q4ZD370
F6+RmIQjlSftKEeO6yRW0AIcDNkwbzCE5O+ghN6Z+Z38zs7nlajHxqxlcobb
7d+RoWJ5d0bJJppBqXIXEszLXJot1IpE4eq0ojTlc6l1NdWZPRf5DZZhR/jf
KIIaVGkuKrK3ybXGjvM7xdaIvk3SlVAYpIvC/heJrYZnKSBwXbzpw8PfG6BN
/3lfCdEc+Qw/jJg2jLPnT7Fj9jcyFP6ory/exZer0aj5iRhujVLBglqiYVbl
MsHV/12NU8T1LS2unURybODFtvlLmjVl/NKwR1yqckG8+rxDzj64ynlxDXkf
SwoCMuK0IrOVvdG/LasTNAzXA/bOkONEhJcbsxOamXb6JibD+ZDCw95JCAyn
r5S5pQTmE2mo7772RjfND3DHCzEchrnao4gfsfdvdP19IGweXYhaRVck0NFB
9axwk2bno6p2IUg04QQhxeP36pVHCkqgsNOH/8nhBRGLzcbafX44C3mz5K5f
1aqicIN3xniC0oCJ7+P/1t2tUEnZdwgFnAgtROlLwfKKEg7sBQHuExlp/lfL
Ea4GSqPSUSqNEh2gZSkDJ+c6qZVM/CkzhRJhDLEkM/kVQ1JIc/cosoHKf8ky
sEdDGprH+SWSLLkGpd0Tw/2MP1Vk0k+NyYH9lYtQNZfnhDLDNNT4VW2SLaNj
swBRChN9oUWyAp53TGogG4zw3p1BHqecjdB17DjFN7JcnJx/rqK06umUa06B
riUC4oriRR7BY8fTbeBsg7tLmA9OII9UVMKyn0CNIiYUcoDqv91SiK7gS3tw
URaNk4dzvDWqh/46eoE/YY+R+zpvgsUejd+4vnuGr8dfCEmJagU9ZbdtqxtY
v5pBMf0o+hAYsSAl0L97jr1kfIu/yJE+/Jjc98D2QM6qbVqr0LC3NVGHb6OQ
f/MR+F6FwMvi2rfXkLcmNg1GUVhi3OhVsXO3KGnTxybmpiEI2BK0DH/R+LnI
QbMFGBJLBR2OheWDos744WEDTrrnTS1zdVYQWBltvc2469lEsvHFkqqfgQ5z
ysOr60X+ZhEJagp0wI9E3JRBMGYn+AEGUH7oKWlxF/Ufc+dhfaJDMi11Ifrg
Imu2yjb6Nv73VnB4s95cTNxyDuPQO8meZf2Mbm7SbPxUd31zmFBwxcdkm4RW
tcWHQNlEppnpa1iWjgx8pjN/ctKqUN7Ap/PWoBrjvI2hl2i0FIkRDIYgpGPp
EEUXUSzJHJtm8nQ0q8efZ4pOS1PWDvCPu8O629SFPD/Ov/oPxjL6ObYKKIUD
2/wrgIhvoLZnmUyjR3Bw/Ywk/4ENEeySshcbx7HbRyYsLweUVdKOrdji8flp
Vt/n7vb5I2u9xEUIdTKdWwzdqTZ4qs31A17dKKUA5Xaf2QBNU+riYfpdiHOW
zJQfz6+mhViDeN8R72LRL/02lBzssFYA39h81WcejFLMGnxOnu00qTyMNGHz
w+Mfn2zFrYVjsOiogc2d4XAYM+GP6HREn0Ea4EkpgA9lE/9ntCQazgwu2huw
jtTePZSxS7JyzbwqZg1CcGaH1nDzP/0Ciq/SzNci5ieVPF9bNYI/Rm24wVAA
cTgC9H/CyzcJ3TTuNNs3eC6ltLyD9GKYqnjU9OjqCs9OGVJgGGWThBSm2qJD
hZmFkPSBK+xObsgJT0kjYbfdkaKQ0Y0Tg7FhyekGgUkkMp54/mfd6ZEeTsdw
zttmpPiTikxkkkUHmlKiuz+L6Cv+PF0f/6V4suuOs2+sMu+00lwhzU1vfCJl
CKakrOrI3S1U0wAY0QXEscwOG9tZerX7LODA4DbG1M/a81IIBngOyPsYbMcB
xhAiLE2HA4c9o8tGINfKldeMplNjGUU+HBiGgmOeVLfZD+6PJcfNrM95uh8w
2TfHz4w0ZqUVkwW1V6fdStzv/i0rOYbAFOL5lMhPd+imKBnphHN8xz2sssK/
KAq1nfubT1TZfcj2p2J/2ZFaed2HBf1194k+b1rdMR6v4Q2iOb+yM1rlAmEf
nsMSi5NzgASf+BL/tQJSDVJ1qghf6i84NLMutRKhfYWY+j64nRYyJC+aqtwx
8oe+Aimom41+dEwvnFhUVKqF6tOY4zf6n4Gyo8pijI5XCtNfDoB0zKouxA+h
+tzTuPRfYJxPLXpeHdbDwXiR29KhiH6FDpPEfpBAlIK43ri/V4G31r2rK1uh
X6mIYLXUmTH1QlCUcBqdWKOZ+npoalzK+9bKV7zRPpz/jBvbLhZ+fbxhgyDB
ZhlFR2DqPGgGoz4lfKl4r/KGI19hVSHE68dd9xdgpl3Koqijq68wwlTMtp9M
Xsu8Mka7WL+5NCxNmBp1zjufGaGAtfEx9KoYd3nU7OxWlT6pBz0pQDaGYcMy
ckT1IHyUsLByNSMiCTjkbcZRp/bBAHIatq/AsOJ0RlZ8v6kVTYHiIV0zoyRX
JQf3Mxho0UgrCSU9jN3pr+UCTHkGBuyc4l5XPU5RVqO3KLH7doJ/S7yS0yBA
F530Dt7eh7KBp3jNQ+kh9eHXuvus1LrMdJJMjPozHN0w6jBvxThbZEuhinHF
ViGLYw+BqbBwaZXZjtFnfZcR1oFE9K9oxJZ0gIIkDzg23gsf54J0q5fG+N4i
HSzLZQ5/C8OAZOVmuG1W+3mhcblmWACwSMjsXibJI30kQreJqNKUYc7DAR2N
a/g/40OrvDckkMktOsqStyPFNJObwoudHP4drOo3gTsBIpEPZWweeZ+y3ryW
/08dNUX1Oh7GYR0HLSzQKlPNHDKoYj2FtlleEZUZMrRTaM8zDYlZDF9nIslt
J9ix9l1drkO8p20dmEQBGmHaMTbGNUbgKEGaPQuRH2NoWMUAgngg0eWrgoPe
qFyf20io4kUGXgJ6ZnwmSrndTbOCIZ0LcDR+mBXrsYcWl3N/wz/XCOnanen3
JgPuMmQ8PfGpqXQUMrC/suiPt9wdX1Z6dahHk1wu00ts6wuNRr2xzvfbzkmj
At0PeGGIgbsUQqTvTL0OSktJi8iMW7SIzfOWTPthUaj2G13oCUT0RjojLyJO
WDAQqvtzb7QoQjrssVvRS/ejwiAdrsz8Sdl8MIQN8q4S9Z9+3YdSGH8+/it/
9z0fWSV2c65aWzU5GDki9rHGNUOZ2aORn85cLC2W8IINMtGUwvlPoD5B9GsA
ylx2I2Ov7Q1aSRkbY+KtF3cfyNlUvszOsPajQqmtUOppTX0woZICMTJKBkyR
yncCnSUCCPMRUo5Dp5oVbzyocUsm5wqej+BZHiz5AssQScOpX9MG3JHHh6x+
rGbAIHTImrvN7C6Kv43OjYI5WDFxA2Wip07vCKgG9B8RAmEO0QMoWd7OMcHR
cG6ybbA4QTwHj15B0Wrpr8FhqtbpiSLhKFkF8ll6V5FgsRBawrRw7HPIijFE
1i5fRCuBc4iI4s6RcJaazwBdZyuwOPbOjlUHKz/wd+eruQTNoV7sXJ5RtodW
P/oi1xuWu53V3DUD0CcABG2uSXSS36YtzmSlSHe0/Kx91QyX2gIlhsZbrR8z
Yi4eLawKKe+ciSG1xEJ14deuBsDYZGPaJ+K4TJ367LZt/XAp7c7nO6YBP+CU
ohtkTicmFxfWETVUBWtZ0CPUEJHFP36y0XzpTEal1rdo2Tllk53uRFNZikdy
1oulMhcBndLkO6yNw7+NGRoB1Jtq1AFWdNdsXPnph7FobgrpstFfPyw6SoSC
Qj1KDQh/inTDWe7S0XTTJU+DQighNPTDQLm12kchweqRhyGhz9/6NkTEod+J
DgTO6R7hEBtD/1NoeOta1+PslwN8pEJybEi5RoJC2gtYKQUXgnJL+BWEmF+D
fNHcVStUlDfVcBupCj5z9sLEwKVjBWNPn8TWbyHXytfs/+GrJPvDlsE7fl3e
MYZyD9iOIopB+fAwV1qzzpSrtGfRtenlAZBn90WsWy2ujkvxSOPy7lj2+hwb
OcZrCfeQO6Dj+7MttVGoz9e0UT141YkbwOUD7kbJHrFIaDsrbEXH3Xg2qa1/
BnEixHDxHmaL38YV9Vt9gE1dTpi9cbh3NuKCxNKBBpELPInlclkMX0VJ9U9i
+SiSwqa+yqbBQ6UbFf5ojWkmbQNUyOxZIwTt/vW1IA40yR5E/FOEzuBhXwx/
QZDYy4MXwr7HBVqEPsQokbwuWrGOlI5/f3DWHrOdkxOjhteXeK7a68PZrnlN
gf9+fJKvP///LUqCyLj7lxyGADcFp0ES5jpUUacWLdlF1TIwJI9D6RPyQEfS
lt+2iklSjKduKol3UsvnEk4BSaKOrdaHwhZelG8XsQ2jmPtvkp+Upby75nxJ
5Wo7h0ADtSD2fJuyU911vGih9eOwFaVA831fRlVB0iBk0SxiUPDLEkRYXL+c
Be9X2/UG//E3CDFoMbkBHeuIYim+7nz2OsAx9Fp6zRTUzPQu+LlnB2UcHLFK
POJ0ghgia7InpVBbnoCedXOFUFp+H75sSkyJ5eVMp7/ajecCcdCaYFC6wtYY
SHSHXFe/8SC708gyPpGEgEiznuYWhyEKqKu/VokMsCqYkDGqP5y0Uq62pHan
vu+DMRxGH2A0KmtZ7kswx5ucP2rVPHg8Nmv/4+ldJgJsX2O2GNJRvzQkoEzx
3Tc6Qiawpd/HCMlX7Re8EdanxXzSsIdsBUGrnJQvoMD4k+eJPDYEY7mtmOtu
Ld7eU9RMLA2oe2elo6q7OMvRY/Hr4V6dyvLxR/FOprzbuy7mrR2lziD1FR22
KbyVtsxPzFbBZndqX4C3u3qi2O9AlVPVH6deeLtRr0kwDvp7rhl8OT0Jl3qM
lGNl7PkooKk4IwSuHbor2RvULtpAdbPA7PRweN2i0uextIaPc8BwG7n1YXox
qjPkR9+AUBx6HKX8FYpPd/ieDgVDBjcPRHav1z1Hw1k4P5cm0HA3hIz9nzsV
evhkRKvkPHyvsttH248JC7w1Q5EHfCUeR8NubBoz5DE5dHKFSgqCrO4Ixyse
dwzYXan18TI2LSvsHeLqK5JX2Ges3LG8a953MjCp7Tcl2XzutuMjiLjVBYiQ
Q0cIjN8QEUs8YR+3wYAW3/aI1pfXuSw60YEuwMNBJVKUig3eRTcpHcPPQIMz
52oMfmvaUmnX72cjPYsTcOKLE8sRSoGfMzGNZ1/lSY9qPq1xH6ceTgXgxfrb
a+2oe1tGR/PCWwek4aqZmnTE/unqAhWZZLgfDly3irhIVfywptcJ/UHZWB8g
E+LZ8WJZlPdPyagdx0qOM/NYQ2aLm9WpR84lvnXkf8p2fPIu4lriSvIqdAGB
abMqLhgy1rnoq+CMcn7NFWoiehg9ZgItxg6z1yw2skwRPfqYEz+2632kTWVu
bSBUBAA9N8o4EEFSwqkdva2M6Pf19n+ZR33BauA35DYxWpZ0E0xGK+4IAvZC
OHM6ap5gfDDCwSz9CidoT6aU1ayw+Ktwdy/L9+LYowjZZBtsiMJ6cEa9sCHE
47D1HJVulz4K0WQbkI5dL3i53pUqvdkx/8ENqeTvi8X4cSsDP6J65p1iSmbG
iLADKw4v/4O2o7ZZy1tK8M4VuJNjFRaIYa0OhAbU8yz9GupnI4essT+rI95H
ko+obzNtvymhSinD8XwoJzgoyrIVlmaCJ7/DTHtlZhBLlteBC1b5N/Nmtn60
meyks/bDF8h07yQ3G/a2U/6U3vfzmhJpoIcXNVTKUuJwK7f1vgUYekAmB9Ui
XExRaIPUuRy+2kl46DjDQ3FfYsRTOstvZJenux/qtckU5YuXLGhUuXZ/O1ht
Hh3MF6XyAWS9IbvKVs2NrkInQbPuIKNO51Q5/rgcBR8aU+iZacrHJt+dTuKz
P4sp79rv7NlMr88uPy00dkGsqS7tEnzUrbKNBJgF24nTkbPztHdxOSwXjsNc
FFxPPBtSMZXkzCG0m9vG6vH39QV+LWieQH4tISoTC30+kE92lblHSho+MEzR
1ZSn0A0mitMd2qS4G9TuMY0LZBVeZF9yEqrKrJtRLJEW2BKcpGA3ohRz3JrL
JbNOIz+lZG2MWY9XKaTpV55YTKRViflQvE1BoFCp7AaADb8/HgpvT/McS5QS
4j9MA5N1FC9hteAYUhI5Tdm5rmrNs5xyu0Od6yAADfRUpfuHrc5gJO56dlSJ
RxGJGv4JoljnZH3Norjo13ZiyoA8+z+NWg/lRDJ0zzkDG6PuvEzeC6+iKrxX
hjBRpLMxzPytF24QbsS1qfvJ836NV2jIr8zPljHT8KnI+L8gdPmJ8dQQG0J9
4ASyJPAZik319xj7JThWRAPznD24V5KgUhaAgu5WUH5owwm94y33fEKaPWTA
Q2bEfjuEv8Qix4YxECmcOm+Zi2DIAYWF3hhTzKqYdeH4xz2V7pAVlzh7FhIR
ustYWFL8GyhFAZy3o3OzlMugn6YhznTo7Tx0S/ht2Vb5xOqRMyf5NILodZrp
p8WsMPbAH4zot1O8rnskuaTqH+Uvks8mdHvkFzEtJKGC3hgRwoXJIpH6Uh4o
S4YypMzKy7eazfFySkASjE0J0VFzk7+9uQsyisMhI9t2LCATkTaW0Xdla2j5
Mf9lYn1XWIT9HPJ8HuuKc5J7fy1frqM5gthcFGUDp2gnP8hUFIJ4ZUr9sQAL
ZAzs2ZKAdrG2NhQUUVFS/RHc38n6v7z3M5RYj2fZm6tft6R+i+t+XvVrKSD8
OZ/w19Axf7UiP9jnZPFS9mv3c0j9qVeF4156yXHINLJymMQ625QKElYUaf1K
kEyXe7vrDF6hKMsKT1rszvts1y4VZ5zB3noFSVY6weo83x60QDfObS6hIzpt
AbQp+tmqzgIBvze/0w7/90kBZGUWo3ycPXeZJhfF5fPz6UXMe1EtU0PPV009
V3Z2JsN0g8tgzSlhxet6BdYzqYhO1fScOoJOb2Us94CN1W1jXuVFOpDEHGwy
zuccQ3mCUMGLpc8vOnHqjv0ViCL4DVMuV2fB0Zwi3DD0Mdjfq6TCh/OV0/31
VqdzBd1JrJngF1d/sBY66AUQN/OvAkEB4fjo+21eCXq7pB4KU2bWabvWVkgd
M22qxTXoGaeqk0CKeveFPXhKhlPUOJ/qagjsflPjbQ39HkOhVPZaCsE6R+u9
VV6N9JIg8i/EsK6IwgnN/HUNs91I8ysUmhS73rxFPwpiDVhuAlOykyTFNxVO
nfktpyHkS1iTGYptmzpg5MS5t192Xv1OYXMsxMTMJKvLnfnrQ4h4queRIvYt
QG7Q5MPjsbaFnb+lkRRMqy0KvOLvoxARyCDk4ZfzzY2enBdg+pS5F9Gm0k1o
zEzssAVTKY0aNDyQMznQ68FGm3I6Ur9eEl/CqOel92rET7OaPx2pB9cssPBb
27pX5xtnZMY8QV96p9bZJuYZ+nAWTueCgeTNMA3kd1R53pKKNkSoVngZO7Gm
i3/PlDXWMXkvepgabOesbaKO5/nrUoxk4E0a0sqfnyL63Ehya4GkOJMtuJAa
0UPKn0oECIFrZq4zF8A/Rm/iThRCXERlQjUNG7i7C6DhOauJwg9MU7Hcj9Y9
ZFzSyTzHqmDVS1UrTAy7krFKt17TzTnHrQIrXYK9XXkAl+zuAaVGN5ywwxVk
MN0fErUUzpyPGmDnh5Sloy/hFgd+8SA7iUFZz7GbnJc3jddrqh5Dsyugo9+B
wuhAgGtrVx+K39+SIH2oKDhxchLYNCrQlElmvdXJQMwd/3uK4Y8H9gRnst2G
tvWby8Y468xlcFbuxqojw567AjL93UZ91+83mAr/lujg2VynRbV78xtA5tGF
YlXt8obtFhkTJJHncmdXwh0oowMZ+Dfsw7udqeF+pV7WcGFVYHFkz9iS93LE
uFa9BiJQ5SOTl1UNR61n7VeolmyFWIjqjGcIuaJEhdvYdGvZ5sBe0UpA2bus
H6Wm40hYxVuWi5LuRXceZPeDTSGZ3yXMib33X2+0A5mjBzNO0CnBHFWVugkW
Lfl1zdxvobCvcGg51zqRiC7j4ZbCbE318WUIgAtU1GI8VxkSlhVVtpIb0yiy
HuPiRbrI/taGe82QZ4UOJrZIG4Xh3nwBhV2UvhpgYuUDOeHEIj25J55GRHF+
K023FxMotpYP8ejl3Dm3jLp+KdHEkCXyLGVPuY8tmOXNDhJMFnqDaHROZCEt
jucNFOXyPFzFZ4o1Z2JfFdYKv3rgqtU7ACVwX7mZFtz5ExuQ1BJ9ZO8rQrar
hzl8t3JTJAOUyEo1OMAkowQSAZ2bsa5ME7Uc7pVPSs0gAEze+5itmuAD/fdU
vdeZ+R2g0WinHZgTPVJ8CaecXgzqe7yV9NqyriGJ6amujPF0T7W8+CE1qLup
oFeTiP8ufwlxGNAWgAtrE4q1I5x4cxEX8hn5CP6GX0oORbTG0O8qRGU+xf7W
jqCSXdKhonmwYUYP6auweJMYhKjPLz/pMOjqQBZkwS6pIrnnvfFhEjsVwMN4
cD07DrR/RVm3fnNDL0IQ0HfVTwz/D8JpLxTUpQaDY5FOhXvnuHsI0iZQFa9i
4HEqyR4O0ydUVZlOywsZxx6lwhOUXULlQf99Gk6zRzjzfZDfH/Ii50NJN2Pu
/28gKqS7dv733DbH/jgyEfquJtD0i+cFE41pqd2wFlkPRYxCpclgk9Q6x9ek
r3ivY40uwFZex6BT2cx/9Msja9j+LqZcYLUsE4Se9Bo7Jij2aMQhEjCnMVT3
anN14N8jgm3Ey52Fyum3wamfs7G1xlMPm1WJzO9Cuhsw/llxNFU3ZuO0GeFL
tz18xacrsRvjekthaSy20X/8RodGVwoeS5AOH9D2fzcfN3/uiPZsxM2rrXUb
eLo5eONEcNKGtkUKhJVkvZbVwEx7eNOsfVSou+a8dYh3AKa8az4yLg3OrIKn
ZSpvEZP7RtuwXAaRsRaFa1gneymttYzkMsEY+XFIZi3mqNs0m4tY57d05xBO
bgHQg3KnnWai9KeKSEpGO71749/u/x1/NxOp6paUttxggpy6puoEG1vSn5U1
kXtPFO2H84eRxzE4gwpNROhIbGhym7Jl5YgTbK3PYCM+y4c7jd58doQk3ur9
L+OzF9smMOG+02mN8VIW3qxhxe39yH6h806SPKFmlWDaxkeuoGyZ6n9hta4x
gedBNYoXaV0SiKsdfacN7N5bz8YIng91RC8pofg6iXva93JB+Z9KjijfHXE4
HJuivw0ysA464kgLjvW9ziG7Hi8s3vGbZpTaBk/28wG8tABdAjCHkx6DRX8j
iUYApMnpHgbA3rhI11TJHR8pSdcsXYGw20dSULOvgOmc7iGasJGpYEh1ryjp
J5PWg21Rrrmx7OTa4+t/1ZuyJV+10qXoO5wuWFGX9gUjSdmgkzSRwgHAHU5Z
q23wC8sfFK81rxUf/eiZHa4mwCwqjdQBTKCbQkOHbkOquOVckI+wMK8Wqw3W
PC6C1MBzAHzNxw3Gt1CS05tdiVPGjQQGTBx5TE1ZKTHE83puR33OC06S+MOy
aqT2m+D4tIHoGLsOXlqqadE5enghhdPPUyNRClcRnSVAGmnx7NIKlKjgnZkD
tJEi2PLXyDH4LxCI156FgOvu2KMkXviVW2gRk6yfO1sr0zFCG7WSNVsTqtl1
j/UOEb8MIGlo8162cPCg+ZGK00Xq3++w4ebOMDI7gyG6v+usvINO+8FoVRM3
7EShZrcpgvuMRfZ5T39QZgTswpFD4QdLf9sn7Fi5pFgcs5fOLOYBWXOPgg4d
ImyYbQ6Ib0OpA8q/zECzyyEO0XzHxS4bpiS7tgD9yWk/uvRB3JXJ7pyu19b+
xfBD4vzRZxfvrAhEa2fGhvJJ0cc2cwYlCUWH3CXIx3Oy4n5CmPoP6ndbPn8V
p2DBje4g9W2dYE/ED615GjuvXIcbjOjfhb9HYakdMiLEaPicsITY247Ngao4
1DfSnM/Np2zCY5luCTKgIThVNQAxg9hgkvSEQr2/a+xhOUYnyGZrMM9glk33
uvD40MaPNk0mEG0kIp32m7bsNw5KFoI5FEGpigotJKuYyiMXlCYilovmOr4/
CbAUQlrbi030M1PfFl252noT+VzgjlW3C540QG+MO1BliVAxm9CIWMZheXef
rV4YIAKM+nzSKnRXfQbKIxjI1Illafrk0tVLIdQfJoqytiFg7NtnLIIbsaYU
qUVsDWvpxA494KFmLTd4eHjAxt6uus/+NxhkA5RAqB38iG/MSrar0DMm8P3n
P1pvpZjFBcHDkiBcVqc3xhgvwQCTVgXYK47OEDCv8W0bpSnUPi82T2DjfI9U
s20fwoNu16kUg6eEZh1ZPPlmTWimhn97tGSEA0EjbAsavLtWEWH0XvOdT2fo
erofS8BBtjmp9riPtRm1GssWskD3ke8e5LYHlHvWzHy2SylHMno87JA0MB/Q
YTCgrN271LBMP67j8nW+eOJLC2h4uKMpfmn7K8lZspEGHf4ciibm7ozfieb/
pfZ3Hy//L9vnl9XXutrFyHa86dXO5McQdlqD16pBDKONjltc4/9PJ2qbcnTE
S3xVL/YzfvXzgCEvV1HauJ9KBO/SrfLmDqNOg1F9LAe82BcuFSf+YlWL3rbs
Snymp+HgzdrKnJoW+I3kjRF3nz+mfNjhJvv0vHuZXIuOUeQCcDSI9CYnLog3
7nOoKmwAYlJHP9pNAIoEQG3qzwWLpvqm3O7jdpiJtCJZ0+O2popinFj9qu/c
y5ZwGlxiW4llsc9PJg3MvwMAlNl8kL+yXD3mKdWCT2Ng98wGBshejAwUr0D7
VHQZGo777Q1TlJqHz5kvZcoQOL3w8PN7RbdnZcBaIqaZmlnlrhCaDyBJJHIG
DvKENPUgUk9YSMg6t1BFZ6qswSw/v7frzZNCv1z4nN3vbP5Cz0IeujN1+VoD
EbbDqo5iJBUkpaU0RaJPycoO6ZVA0BdxDI+2u4aRx8r06O4+BX9ia7ksv64W
t4W6ieyXKS2So8iJZBfKLNkFLh6Zvx11KnODyxg9ZbCJGqMSiga2yNShICuj
cMAnhlWrna4h+YxgVr7XwhUtn1VynhiT5J1GEPEALbpkEehsLGzBJuxR4Kuz
RmF2TaGEt5sbzbnavExUzgr6Gsu5EAg1ez8RBauJQYdKfRAHZWVxHsCTJttz
z4I0ht/pWEbUrVVIsjsy10HwfMjhOoB+6ZPl4LnVurcB/QjQgXC0eOpAvFXe
j2Z8Dmy8ybcR/t6PK/Pfv3U05nUqGztLs5/1h0lVoL3TtgM5N7LvyBxRjFpN
1m9q5DrEl2gg5zfALHUGgeesUF682v7RWvh56r8Al3+Sdpmaz247cyksdVnj
exP8RAJ0Lmk24hO6OmGgezrJbuMZdVZCY13aFrnJNBByp+z97DKfmUrKKAZE
dnpTmNYOiLkEhFcjvOgq3g5MjWLDGJtnNN7xXIDxnoJ3vw8J15rI6s70woDY
NRSe/KF++m9nEGnxK8JD7xY7RiwAJpoPHqJIh5R/AKlzYV3d62y6Jh8lpmSS
rMNCoVUHQrkq2RKLjgHxjVdP5lmWFeSlxqPNKo+IQYh2VXO66vbdfnoUWrxf
WmES8bEYeCXvVNbhKQfBYnvT08G1/FVJRegUNTasXOM8cQHyNvoyNM4LQMFT
bf/j6t1sNz2fX89NpaGqZ+y+M3JbkEjejeREC0HlO5hNwpW/yeX0ZfZA2O+t
tA5cj428o783dwJ6bVUsbPwXSv6SfiG3vRxssJcKPWeRyPMGIbggpFTPImjB
QbFktuSX9jdyh7hzxcHgTnS2TTfPMNrnoAo+omumNO30Gp8p3b3Xi8xhVeVn
FsWoZ6oTvIhHkKJCXuBOnse/ghrdMqrcEBJglSAWtlZdic4GfWZxS0iLlUHg
NfpCULkiJCk1VyBtcZRtX3E0kWbXehk21WoT+VjvVbDHR3DNCsV1MlCJeCYs
m6yAb7oHStMWZOebHlvVM6yM/Hl/EfrgKIeSzL/Wc54B7E3uH5Tk4Lx4Jvpj
j23lo2cA7agiSXm23K5xJRPyEaxJdCMAtuTFud9xcWspbc2jpg9UIvcjZYU/
uxJ7wsrowNkPKyJ5dRncuy7Aq90lbo+HFBeWDlO8/e5mNQlIng9uuZ5iJwLC
VO8BoCJr7FduhCJQvaA5YJxEm7ICqNdOQxfVmrxZcs4Q9NidR9eWk0QLo/mL
i1RW35EaNWp8TfAmFN1IArXfxKgBq+ImoEYNVKSCK582r2uQnlwxuY30rU3s
fvrgsFRiVVfoFoqfKQkRn2UwsvsrWk4i91whPQ++b2n1Eg2/3diIad+BazSH
YqEQVs+V4Ao2lU+yHd3fJfVNybCj4x8xmvunWFklwL9pveDNCGYUQR2FLwtY
fk9PsQ7qHnylaxnXp0f6rLm8UlubEB+6u3U3T3tCPQWcsnLICJ1wFbfznYJV
oSyx9eApDHQdUNrJyI4DVEfnzzYqqWFOE4vDEyliOXNeeEwOxBOjeARgIzOR
ueQWgGqVdhtUbq/mNvOc4v89YnjsqCiVWt9dpgCpcBVulH7BKwb9Xm+XIpp0
a/tMXLuWrQkhUrJAWWdF+QfC3a2PcuN2BO/qpIDYPhobNMOEVwiFMSeoZf5k
5rn3IsZ2kLTvfrkHw1vNTJhxDncEcsuJE3sJa2ewQfAd4Yw1eyJ/oIDV+Uu+
8Mn+cWrjAE/spMxf12+ZdFgLCCBzE/RAtQqi2RoIwNkme7TLntQXvM8d6okO
WV9HkkuHey/o6sXX7UKoh08YUxc5DXsgWtpnHf4+ChziUu7YYzcc/HbnzrTZ
Ph6ZcQIMRBVe/Z3zF72IN0jhl8/cLDZ8FKJ1bUumvoRlmEu57PDLfAilursl
+Er88Ws2/VPwp/8vrct4UM1EEPfAjU7vzqg2v0dJl8NBp8s1JOGHod5oR0WH
RAwbuvKazcx5dE47355G11tqqQjrYhqxTFUuYTLYg1YIQzt5RvnVtLSYU2yX
6BU1gZRZ4yqjpfJjg/t1KZv9frmR7aoWtWkx0jEBESmiFbq/sWd2v2WzGelK
Y+SkDHWR9A4wrUnmKh4qYTyyOUQQ34oPxxwi3n6uaId5cBKWOLcrUJrwmk6A
zXJ4GYF0Bgv5Lk3FS3COuyodTF+bdbNnuy01hNJTpseruF4pHyx+M2xTCXdu
MDNr7p8gU4Y3aBE/Y3KSXYUW08DTP86/heqQuG/j5lRDntmHUetSmzLA5qJA
aQjQZhjbGgtRc0JCsFsbt16LA4n52yrpMzmEy5dsHcvxo8xKG45nRqpy2ynW
YoQOvv0eWCk+Maq0k0+fkFClz0ouD4No6+5q2JrYOzXYrFIG8eC7fPak8ew0
0Ce1Boz0/KQAoY5QIx5twrMjMuvbynV6sAcsOTwbbB8UdWZh836NMWGbB35f
fjliNE1v4Rbn8Suobqjv4q3brNFjexYYMBAjKDCQQVsgxEPijp1kN7qowYWf
CDYes4BaWdA6PAPIq8kRZLrcEuiPVAPQJrtezttLiDdy+Sn4ZyUvuV+Fuyz9
jmtqbPwU4vinW9S3LJxZiA1zoO8Pqc9XOSWy2D26n1rcVRKbY61SuC5Faf5A
SeGChzopKznsXK0xvPNZBczWUiW00LjOKePMJwE9RfBArJOJ0QWflr0KZx+k
ViGninBseITfk1wcjyZlK7tURT2GjCQbnLOa6DLQX2tLzhN5J7MOQwPaQJzR
aVgGx3gpZAijNCyiQi7gc39DRp9c3HL3O8wEcCIyF//XfTC3W2cGxdI7rkGd
edBMxMPsL8ghX6ZTof1BTw/1PKZlryKJ0d0Yfl7+SUJrfk8+uPcQ3tA7a9KY
gS+fjK7fovzw4qn65xmCuCxXlAs9osq0zKhVdPmHHn6ikZkPKf7P7MruBcNd
oTgKqHl1JwceLHqm7Bra0E978g2o3BK8yidqg0luGHVaQi0diEVTUeYhTBUj
7xHGu+UylFjnWvwvR5OkzJ61A+ZYv6x7IR+y1deRpR9so/J75okmHf/lm4at
CCWzneoL9YOp7lF4rojZ37CwgNqCac0EcATNTPbX0Cq5yFlbEbUueAfS8oEl
MSZTibVcCfpSZu84biE37aAfgi2+th15m/Hs1FKFcSfTK4rE/kZoMEVHafBE
RXCmyxx+BRk2TrEqzh9Yng0WR6I/jvrhunmjLAJfpsDm8D9doXV9S/4tDP5f
GJA7PTBk0sdl1FOdnhNaAGX88vlddm++O7nTchvrcdcr/BhwwGrbmviXPnB0
Vyt9Tbh3sdczkrEaLETKOB8wfQ7HrzqjaXrecqzwxUuGjZcmq1tNCPsZnKzU
06JwURfIl890luHtkvkshHbkF+BznSNMjKADpSlj2TjwiQLHeWhglzwVMBPR
sjGdpQNot/qSw7/6/RZcpFvX+C4kodyj9A1tc6IREMzg1DCcRFMkPJtsc3DS
1ACZbHAKIQNJGb6eWGi10GxFafIA2jz/iKtwXJf5l3kds6bOtIhadTrP7+az
qkXwUtEasWnnEk3DZYqoFP+MfdGDc9sS7DlNbZcD7+GoTPQogPh4BsdL6wzh
fPyja+2f/aIXimDMXdd0iiq+QOjHZWUcj+MQ+hCaPuLcwNUC/axEUYFllayS
ZjRZR7UtzpMe9hXuFFiAoTfQ3cEfNaYLKFDmSjBMLR38bzLBuF4JvgNoLrcn
pMIqG/aNR5OLYsBi9R25AyYZBI5Yhi9L1WEKqW7wE8CE45tVUtHW1C7spOZQ
ujMO6qJ4KoQaU3nIPwzDc2N4XvTG8/xRtApcuk+C5OnbLAPECGsBdCsSjZ58
iBmhrMiQCNYXD6As7wPOqhIvfx76r2hvLaIDDghm0EZEapH/IeiPYTRw8Bm7
d5/NLuT39uCIE8mAkrMiqGpR+cHA1PznVrzHVvWPQi1+sS5/i36ahEe5CFox
1flf/5kozHwNL8Jw3J2Z1xBWv8Kxfy9sYgPRBWdyN+6LYCOU6lBBib/mZttt
ODFLn4ruEgfFTLzIEVfmqa9/1EONB6dBrOa5+2I6aRRVNIgF2TKQFceCr0qg
AkEYiI1UWdRJRbtsUTaLOfum/a9+RM/iylKAD0Yg18mAtAwbpFj1tZflXcyf
/meIrlhRR0QCowHAbAtj5Cbb5d6NfvuDz23CHztP8y9kilws+Vqr12j8cdyA
XxNmg4cYa5Y6xNwJmxga3mGMwus58/4U89wGk6oUv7cJPkV8hLdyImvloGuJ
fwv3M3hml2drnYhzmZk+wZxKlA/o2Yagkd5rPzcNJgQDBeDesDQbNc1zn8+A
4dLRhxNljajBbKnsvvdskTpJ0a5LsgGHYVQQd2Z6sLLCNqxlS76p8uzDTxbV
mZ6hrbsUmNftWhEaq9G3mmCYGmTzcHhijXv+9HixRLrsoMyxzgJ+I/kmfWe4
xTAesjK5m74fprmABzSUKXP8/2nbASNZiHGbR6vNNbUYvPBHFnWArQPQihEw
0CQSmtzlDGwwBUPWpEUtDJUsSwgH+KYfphw/haRPf1TDEtINlTQdvCZRNi2f
ygiTGMnDEBDWZbAF2RlpZ6miT6EAazwmn+L9g2AHfV7xljKhbqut5Xk4/kLo
tH79UQya+xzfgvA9lc/TfMGJ1j8e/LcUfgFH2Hu0o+DgMzPmWPy2f309IjX/
GvAfVnwNMPQqjOb9hJ1Fym6E3sL+PljePAvD/uRvmv8YmkaUr9Zf4L0QSatq
JDfV0Q0BBu1uSHciD9nYrAKwfmMdVYO0kIqXvXCgdnA+TbG1ImfGXN5HVdrw
H8Nn1T9jQgToME/nJoyoZAstpqPT4a6cCSo4lUpFF2mAGHDv3d/tr+yOEhFW
98+cipYp11LU9Gw0tABgzbeEm5EPc3RcqMqXAkv/VPZzA2vsP6fBpzfG0Kyh
FeaHdPRdA90ATtB4jGMMpq/QnVxcug9LLS+sklb2nzsBz6DWveRI1uvg1YUw
NoPyByfvnr001cFwYlad1WwcEY9+2Tc0WCMRBMIx97/m4kRLe5Wmirt7PzxJ
PBDuC68wDdwVwD7opev06fFA2qhEYYc0KgbFk9OwoRxj/mbqO5F1ERViD3Xg
UIo8CXGign0yAcVMVqkL/9SlfIBT3nz6d3LBiPl7N8wQ7hfGqeFBqrA1ohEO
pln1kjQM/y8vgUtIzXt+jeuvKO2sCTHoxhSagGoKAc754duhq5f1jsU1YeNs
BhPY8cZ5/oZuXT6iWYOUTcdwF1sOLLlJuqOTSy+oaiXMHtJYR4Ofa+JgsrNi
GIH7NNAG2nmJfhbuRA6bPNKB8Ii11Qrihp2QB9BWSPATH9dh7Sof1pmFy9Wa
STTOSIIEMgbs5W2iNfG186xPHHPFSmySWcgVirC1ZlYyQm6p/hvzzMccmqDD
WvkJNyBRtsgBOiHX0zID1u2vNHpNebehudo9NE99Xttprt0qg9t6/kKaq2ly
3S1IbPHOAHnSRNZVd9mG78y0yhWJFtGR74DA3Z5L46HSbgnQkhLYAfoIGYZL
LwJaq82FECgODEOEB9R6jlH5ixaCc0tL75CqjmXbtxmEolLBw5hA5RAf8ZEm
btbGL8tlqqa/Yvmcece+hMrR9/aP0e9iGl8RJv7Q+2fGulON7kFcvLWCiKPf
I4TF5RjdiRnD5Y+2nB1/1rF8oCTrHOv2Vut02lE1WuRQLKU/ilShLtB8XOf4
k2ctBZepViJhOU0T7HZpugcXEHKBkLTkeBwaKJPm+SS//JZ4FFFzQgrrirG4
weaA581AHALOaG/q5Co8juAJDnHeaTOXhel0t6m8Jt/f6sMRc8gricRXORMT
4U5ECrfdk5yQi12ihSHeCegw2ECCADFFScvNBsmmTfDw3bs5IgE5yQYWx0X3
4ppz2q9bWfAzLpmHuc4ik2eEe99Im6cAwoMa1IoK0Wc57/tfYeHjNZ+xRlvo
aqv3b1ym9KJZHLGfIX3M2BaHKhIQ+Q25I3Ek+3TsDBs9P3q5z3Xtv5L0uFxC
/HgaXLG3EGt12jYT5HQyh1TVoGK7igpmwsGtMW0Ek8GpoT/53oW2WXpUhd35
D3fQF4CtnSjnQ1RLfrBazWwfOs5L8Xh+Fz8pZKVvA/4qFQayDD4CwFumDari
ljLo0afTjxo2zUlnGQt5VF/vnB+yanNyRwFWQkqcUWyDPuHxe7docMcG/kEL
VpF7OJtqZJL9D4J4ZNb/8E6CX5Qq1TGPm9Utb3Rrv9YNUcv8k6yK4+NS0RJ8
nhRQCx6daUKvH95XY41lx8vRcFyVjV7MvDHPwpN9DAr9FyJ+YiHHOgIIHgIc
Ygpq2LMSnfFFkiUUAs27HUG/NYTDYsKSZjrgEUVv9UcNrFojO5BA2sLoGrBX
Zyq4w/wTFXCkMGV6YKRXtMlvgfosraVPDnrr1Xl0UY/iRL9yPgLDj+vs0Alv
4iGHC67kJZ4hvHHb8ym9T2uHekxz6VZLrZv4o7ELox5rdP7UWGuNTJdt9TMp
OsNfr8VBnl1jF4XiOkmUBqxSOIcKsA/Li1Ft8jf7oUZOTW3/O0LdCQHhehn/
WTFUbxFR3NCzBhfk1eoou7R2TPIE/2iIGhHCs64Bb6q98tkBz+xE7M4IUCy9
3UxVPWNqTVQPib1FrZcYno1MDB2nExoy91ipw4xxCmPp9TnuXVBptWvN+eMe
RHARElGw1vWCLxZZnaYaJRq1ZCjlvrmoiuiKhn84IM4O0rPDLi34VcaM/FK+
8bhWsTjkeMMBtDkEYQKhNB6M9MS9DA/jzYZ7p89DL6XfbsNZn4kvExI22EiA
qn0QHQditg6tcAdpYCyCNQaLabg=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "t4xPJbmEH6v4SVL0gN6FMeKrn4IhP8uxgDEXixmWFrfkRmUmHah0woCI0NWn4jNi29PHRr8qC3E+56ObAVSYSIpu2luY1Ux8HxJTmEZp8dfWiQKOAKoquE/rRpOs7kTiASgRERfy/4yFwiIwBiIeSiYycsrshs/YcSPLGlUvkeFONkowA1F3QkwXAeAdMdMqD0IZHCYUiyRDun/uIWwwqKpaY0MedDAF1dXVq3jdOlleT4+y/XZ3xBZeW1LelES8J5OwvQbkXPZiDaEzRhMSB9Knzt2+EmOLs7irnp2ZWk4wsZlBJ0vd9i7/IPf16dQXrUSqH78DHvSIQU3/FzQXL2ro0DSSTllNiq2PLAR1TmtYOTQMSwG0Dj+VWwRP5MmuhyfkzFov5sAAk/9Rn1IkgL3J3pTlvE2QMUIomSULi5bCX23K03Svd0ulOWF+DMmzTHMGnJuIU/2wHCPIL9INC2mRC96ddUOMk0VBqLz9zql1slPK5kiTXTwwAvQ3ZbM/KfQKxhnvZUfdBNHZ3WjK/S6K14bDUAbajKHILVcIeLAJUFWHQVY3UAc9XYYxwFbkvx9QMjZilnuOdLg59T/URwiDNh2uOAuGiE3h67/YpxWg5ao88wnQCbioznTpr7XUWcYfXXxsLeAB87+5lkwcth18FWWDoxfD+HMcZ2QhxFydpasiOpIsh6DTx4hieIgMWJUGhEAGAOibAkILTf/n7kO3BvbmOj6g+BSH7j5JkkBD4Wq8l/NLJ8zAH66Rj7Wek7WaHUaPmXnK5s4RESBZWgFJm0GkOfGfWDVs2koXAsTpph2ekh6lb/qpNd6yNw55p29+JeToryEZVIX6iTkuHddO+lZDDjMkrmu+hYJKS64tOMg0bi2FXvX8mI4/DWevbZbNKlwG4YWRA+uDBZWBPF5WcNUKm1lnE/q0PkNNjBVq3h4awVuc82cZfLO1aNB7YRT+EK/y6tCXJejmeQiVfBrEgZ9TrvdGbOZCOI1pVqT6R5CanUBOpUnzxPHT7ZL7"
`endif