//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jd28VKw/ax5Qb2JzBTOG3OFomqCR3s0DTykkhPIu6eWXsCiERZUylvTmy12r
TmrRd4oLKAyb216YdqqO5GO2H/gZ09tXFZ/i6Tm5MnfS3ATm5kBRPWhlC96/
zmkXwDZvuD8CNAdxe0trxUkCMQIoxg380NmfFs/GsvNR18ZN/Y+B/oan2UrP
lRcqbgXshdUezPcrHeH6M/+H4KKGt6Wq385Ofj3j40fZ1M79V5lTYt31yLKo
iqLeMw8pvcEGMI8iwf1MpVA9aX32A19UPxhLNg75OSTcaL18YvSS/xPDY5S3
8G+5Aqmm3ANGtn3zk5PVE4b89/NfxVSBHNAteiPCcQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oa5CFMyYq+mqfdAuy3N/QJ2QPssHqXpXQGzyLxQ6EmqRwX3Ct/eLmtaYe8Wi
6n4sTUfWWt4Z42AJPDKSe1Mdn0P1iPPyNFP3ppFe3Ph4QEYXqGv7l8L5HIgs
IFqc6ZtrVSaOGhT1UVRk1j9NMvXpisUPQs7bJLJ6AmT3GMDT7ZZBIjwYTJ2n
gaahqdsxABQM1OHVlBU2DXppliBr1V0J17MxJtik0TijEIYejU21uuFPZzdQ
jszDojdI6a6wwo78PQjmkjPNhv1qPEjpxo59g8abfwIb6kTX3dkNhZhBvkrm
QTqcFOmnJD0J4r1W+dctYFrMLGi1ogDngSOhLWlFrg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
HU4NS0BsDDZTmE6KjiXimTEVDV56CyrBarUolyK3HljcJutPipv4rTVV3Qln
XO5VtDqvX83JV3lqvMpVaHUtj3MkvY+6JqI5d5oijPc3pJb22hJ6SbE4pCAX
2iYBAQULLvzD7nJdG0nA/+SfLK/e1jyGT+I9TyqLc1pB+rhzQKcxE1AgetC9
Lrto/rnUGQ48KICJXf/8jcpdPOK1EVHzeMrmxgO1FU3hnQyxcxWjYPGRzvVD
+pLCkDQNI70r6sIO8jHCfQyXPwe/lCwXZbITBHB0GUx6pt7nHNjOcA91PJvr
6T3d8kU2NtGkNRi2jTpXqEuNS0RFjErusN8t+gl+Iw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nQmkFj5io+REBbIiBoFXJuOxDjokD3LOoL1aQ7mVlCBHw//swGUlpdex7zwD
BMpGq/kI3SywlVPRg3mc4lPksQXA3DGzItUeCs8Re2qXdaUkKMdKApaCLc8R
d2vsOIWg9+TmF6MF2qnRukIWMbTGB5Od5Q1GjXqzPmCz5uKYSmY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
UQ0AtuoeeRvvmjhvyTe4puo1wARMunkY2Gr8ZU44dyBl24ignglFipee6oIG
KeM/fWFhk60wfY8sIL6VVxFIOwXgVN+o1Tren1ALRUWtdKj7mcoGwIQF3Jlm
KRMgsPUuIcda/2lTY1ozvpzhdGJsbUKq36UyZdG38ShE0XhD8e5aWn1sAXAJ
6uonNawgTeQZ7Z4MYsC9Lewr7gvCpF38NsUXJNDOejwx1RRW/9SLYcisSmEF
AhbBeMXr2hQtdVuJZe8Qna1IIH++7qCQFsD/ksjzFQF+BT+i5lbUC36VAJIQ
eczhhn/z+ZX3bmUuYVNEHViiFF7o9Hpr8SfjuFauSyjq5C5iavCj+NNIXjG8
naVrQQfLve4Pe1p5uhpML23a/yY7CkejrGi/utqhDmincYG8zLUaaCuSALW6
kt4IHKxb7jRo8UqJaS8/QdnRBu8qygkF31x72CEQzrcoIKrm1zEDB3V9vlGc
Vb7XOC4vqgWat5mKssGEkcHBliYGikB6


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dv34hmUnNc6MNRfxm2BGOke2qB7NhAc6BS/iQl2E3omMHylfFmK2lOHhAkV2
VnW1ERoG1793GN4sBgYTMiFZvoc3x9io7bsbrpJfNPFrFiebeOW/zt1Wwp8E
e/HSUiTPE0a0UfJz0Drilu81SJMCGFygEZ94B59wRTS1SNtTFh8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YH0nbVMfMCpdqG3g/5UblzPj/hf8ZiklmxCjy1fE7Uu6EAo3T5p8drY3fg1J
+uPRIl0Pba9nWRm2vmAgW2iN0Vm1uiL99EYyKH+tcG1gWwmBa/f7NdqJD5qk
VIXLg/JTE3DkdNCrbW/Qkb79te8etsjJ0aDt82e3gTw29myJqaw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2672)
`pragma protect data_block
CI5C5SjKM6ntQE9ho3hGImh5Nt7Ys9EGKSVBeWL6kGEZH8AHJtHCXTMWOVPN
2kE1pcJuvxZc/WYKB38FYPpCEWDFJAKOvTDqWSIPjS6tqth06ud1TGpF0qqI
3c60l87HRfY38vylxeD7ZOPIf4KaoiHushIsEE3k4P4PUNr15rNMVIuDopjn
46uIS/X3hYNEIDyCNEqDDJMHXU6IAFjHXCtTFKcwWHbtM5lAKg0SCroiZkzJ
K26t+IJ7XSqoj4MFl3SZJqVrQv6JkQULaq/0UBllmEPM80rKbZqN4Uwj30Ha
Xzz0G14WKRnosgf215Qh4XHdObV4xy2j5Rx5N/7ghg8RjJgeZT1ckpEex+Fj
0tJjp4m06HQwm7fd6rlSvBD/83FUaIo+/YLi4rF2aPtqnmxJ6IC8gwnoPWwk
FRTA/h8EZwUNox+okQonyFeog0+Pcl3H1gVmmhm87lqo94P6ueTCba2NoJdw
m6ll1K2Zi2W6pzqS+DTlrZ1z7HefmfvzdWA3A6j/IFzwsGq/bAJW/6A45jSy
d90o9nY3dnVVZVNEpcQ5DjBanqM4YM9dRhAZSVvtHW4VuUWnZUtGamvQKxdZ
DtvI2rwLwXv2cUymm5R22/5nb0GoIaUSUIGGnE1ERXeOYjl8Gh6l4ftWa5u8
nWEhgy1UOVPfx9fRF8lFddYi3d9M0ZOUBq+CxfCRsl0vEwE/+bGphOY0U2pV
PTP1yv+7MxFPFvj8qcs8C7DeGUaYvnSoBUJYbWDa+9KevDqpzUR0p4z/59eX
YOd2vu4/m0xNxMWYi+hnzmeZkgqp5pXZEVSfQSDaC2MsBQ9hvb7gdhlg7k3a
8Twg+m+httrGEs+L69eR1CpTiYOntD5j8Oufw56hzPTWH4dZQ0JEyciM9U9P
AB+8hI8qNoaV2HQBXDhna0ZkIqJPh8Ph3B/mGrzNj8gMUzmajLqj+9Dz5aKR
6jM2fbuLOj7GkdHOQh1V0IQnnLC0gen+6yot1OWSa43zH5V7cgMaplgmVHFw
C3Yoy1r1CkWpUvLXC+78whK/8+1PSAzV6Hi7KrdmLZ77sx3DaQZPmyl7f41P
pH5ocFE8nuLnfp7MRnEatEPvNQFfnqc1PY9Az4KqlEBNv0VhW/mDspt8hie+
NhmR6Xg6sbLzksBZP7vacZuxVW2KpFb653zPiUZo/epTPNu/JRlGdDCGsIvb
x4H8Eet66t1bfBGMRCm+4ZRhS2OZuuTSYf9FRpa2KVbDqTGPWXHn4hFX1WCz
+EAwJiV7DpA71FDEws5oA7LLU/LErPcLPGbWzPGgmtcRx2zRJ6SWwcbuv+zA
o9ar4j6UWN5ADaxenVPNTyFmA4xs6nzV5eHe7ZTiFIWXZKpoyjjufggq998z
EyFvehNrGW83ncK7Pm5FMXoh2HCPHAavkieH6YqDlCymKtvNTTG9xy8hnRwy
CxH9SZgTKiM9D9zAqqxzacsf3lhJU42g18/kZHhJdVWgQBv1hy68GILverRD
dLSw3d2MuFMqGSwamlqFXfGrjIvYKmkXo5TCse8BgMynOtU6ejcbY6MMlP82
pNeWUyTgWumq04JKxWUZAisQ+2swsNfWZFK4mNpt8QD+PcIrjfkNl9kkURrh
QVaqDcXHTFtaxZPLQV7mrrFc05pSPREIWiJ5WWovWNf+d6BW1S+N1Z+0NFVi
jh5iDAYsf/1P5QgJr1LE29Z+cQ88/XV7ffrynwkSbetEQv59xofdOkL/tTMH
dM2chnxX3sKOu+YbOqSYpS2WdgLHDyt/5VLIeL2tvOpQMC9LqUjXwJeQoe2H
+FVVino3x7MMxdpgXsyspeY560eMZEhfAiVlmbpSI07uxCiLiEFy2lNr9OMY
ZBxD7rxR4ke9WTwaX9AARYu5H9lNCK6z/f4aZ1LhEtpJlClgYAoknxOJkYlo
v+2JaP4ASR38e3UWuda1/blZI35n10goFEQBm0jI5bPn0/nu7vvhsZ4W058r
rDK7sGAm6UuZPEVS5NhZy0Gy/9VHgSvb0xgiU2EdmUVsnzKL+kQEZNSAc1j7
dNZtyezAudiCPmf7BtC8pteCm/PPKkYOacMYMnFjqXZ6ikBFzP+9/49kc6v+
rsw9NLzDEmHv3jYEB7uwopqoU3ef8Y8Cqpn9ZqnYe/tN0Bn2a42WeI+xZ6Hv
mHRq5H/uDovCgfrxR+dVO2aygyFi+pI7D3HS6H4iDxblpo1YFJ8VECBoYZpU
ULDhTUZSXbBO7QIypITH/I29PwmJ6CdTQGUJTOXBNy3HLs0L/X9/j6i4sUfB
vM2bLmMvt46i/JM5xF4e7+rPRyiWXzCLm7f4ZNeQ7k3awe+BS31DdiyBw4pl
5mZsoy/7OOtW3gbi6wC6b/xyCoUNom11ofIjL7ORwpPWOPftSrytJXfSJAhG
+OYjLn5cKVveIEynsFLKGCkpWfqn7WTxv7vwHA7ke8ExF1AznWH9hp25m5GV
FES96VTbOMA27NCrnXCqZZo0kdnnqKogFz8jQrj4gopnFlvrjelu2HuzwRvf
CxNatvNqbfwjmxMdEMDpwPeMtXNwbL3ZJTc1A2FOhzQFxKYU24VsK5TMY8J7
XzmHdWz5iESyUUsUdL8BdKe2rtGbWFeEvNEBi4M2lYZnZhjFDLLrEZK7H6eg
3dD/7DAX2s6KmAX8hKDQOpL9ZFWZ5MKZJ1FhlkPV0UeB02ADFouF2yfDnry7
DqB3PnRO1CSOSNxXvtt8SUaRloKPLa1kl8XzBlbyRLE3b4F3qnlDeVUzcT3T
vKgEVkJfnt8yFnHcjIa8tojgXgj6qRW/b+puZ8roO/yXCOEEtfOnDYKnth/d
U0DGcXCN6lSPskILJD7W6cM1G/g9wB9T8iWEEAW83DZGUUcGN/XHjgk0roSt
j7xJQ8Jm9thG9FmdpMyrNJfap31U9u2loyrXghAcRer8KL2TUTyjPso8ec8f
RHvgieP+ubHp9XQezvuU1HVGS253ygjju2CDuzTi5GE+tP4djKsL0KA3WazF
o1RgwGneljQhqr6rMNiFia/WRru7qdaodM+9SgH/ZYQew+HQ+drv5CITyq9E
nq1rVPWDK/d7M62F5z4UbpR5zL/vE+ENGPTXG03K6uLnWOjr+DkuPgQg+wTi
vuu9TxGDVEMdVsO06VK1qjZIoPDyaK9rKFr2W2RMYmiz+YohX/Xp/2/XCJ6M
pn9q9Zml1KMNg4s3hJtarl7Uhzq/er790ZAw67nHW6thFmer0veU+oNEBYZX
A9I56y69BPE7W8sdZMQvjjMNBkN5eBA9pi+ZHCHVfjRoLZCGfBDaOrQv3xTl
eQQ1izc68zhxCFMFFRL7V+arH06n4wodYztS/vGVsiqK4qvi88lMLBn3I7HI
n6h5jc/yify9jErg9VXTen9DUPScZzAmffFbg+MyiMQLbtsAvdz7mBqLRrwB
FBkP2PNrULLbZNHMAoqU9yJe93ANBkt8u4ZWqtmMJDthTeUIhAyGr7BL2UDO
oEYuAKoB8G6T9KLNOHE99g00AteKgU6141BnW6MFBV7SFBqu2ONlO69GHclM
vQkU1rtPIoytI4+eZuGmKKY=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+kzOfSKOcJtOuUMJ3sA9pfvCiRV5Z7MkB9fUTNHvkuS76OQMsU4LfPUl0m8+Wij1YUcvbIpDNp2IOCtIDqCHc5ZFuThKQJMb5UKKn4IKnNiTjQi1ghNGiz18zyAcHM3ud4S7dnVRQZz4zBFSpk0BNsJI/UayAXEfFkynfqYEiysE3Ai0XrWs99mDWzmx2+X2FDoBRVJyLuTKZL9MolOfEKpPdg0oqqebI3vW5VS0I0ORbd3ehd9NOuhPADIVJPwci++5HMWkhezVlF7FmND1yyDRZyRYjsi7Q1YOe8+pGpt4OMUtC71kgZvzyzqai6YquK+2AA4BxF0qzMJbYtpbBWbma8dZNHWyhrgq8oZpYX9wAP+xnLYy62WmOxL+adx+G5VW08i+jI8DrFu8DS1dwIccRPAMvoDf5kQlrkMXdFNJWWvpmhWqdnZkjZ+4ni29Nxa2h6sGUBLjBR3RoE8b3ONGBvaeMc2qr/Wv/Q5/TPm47itrVvTM5eTnjdThN5ndTrhzN6aV9xsCed/tyZbFmo930so9FIStuT5UHjjcbQ8z4nng4WeUjZbOKiakxbDcovjX1zgaSsLv6vSSi2hKwCsFbAATJTg20pj8lt+Rksw0tHUcwll/V46YrVNdTU+oiq4vyl6/Sp3hzGEnJ06uWp3Q16CeBxh63dEuYFNFJEb5GaFa9Z+E3xrgz1K1aKpFGc5DNrnx6me9LXRGWMwmAjJAeAWxHOtF72f0s6DJturuFcbPQvNnC6xGj+u155adGK814r4UP4QrKObQBWCnyMk"
`endif