// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VwBB1TjVGTk4aI06LU4o5Ak1ByEZ9ObCrosQc1gu0DiNT611R2uRqcR7lDLT
VISqHn8gfRjoZz+aKl3rH2m5BJtQcsnx0Fpm6mQmUm8SR/traxhsIIsL1Wwr
zBIj7dK2/dTgdTrW7wBs6HZzP1w6qADO1d21Du8pfVlt0E0Vjqyf2kd5ocJt
CJx8Boy7BZe5orDfAxbkiAykbhJFONfGpu8HWNt+yPJdurEMj1EIhh9cDm+r
Xu1c3if0Ng6agp4fNBGBjYpFxMmYWbePDjuDtW7qs+s8ef4bSDWLFcYHo25O
npOBq3EsxvHfTIpxSpTzpm+wMP45fFhepsMgsGkp8w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TNuPQV1kr/z2XZxAOTadXGEMXrwd+FthxNAxl+n7/scD2Qq90VHTauni398L
yGv7GHOboVFoHsBB+V1UXtOxNNPucixu8g2xF/ceudf+xDJRA/CJuEulrvQo
k8z+JZr7IiPrCH6TA6wEvqkVbslnhMdC7tdYNsK08zzWGIs1csO+70xGoqRu
PmkPCYfbLzbJbYUUDU/lovi5xAUDw7psuMaulgLobvkIjeW/wIcHmfFzpqmP
1rLjJd7zmiAidUNnBmTmQ9T163YoeWFn57G0j3DRKHvmyJRcmlVz/p9RxJHx
SMtYU2YQOfjp5HhXP9LHsLNJeQgEFS0sw7Sf23fIeA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DDmi3lCWvAZkHQwcOCJrTKZPSjEk60lP1KvYiSecm6WK6Bf5OCKTxaec2puo
1DrAfvSttvuoo14BQL+SWZaaSXlPOvwDmUIZDOCs6aTvjOu6rAQ/8MeIZhCw
QZu3yGKgdROFlZoBUDUET2qnn42L+HMR1Cw/tEM1pd/jGLMG4lZWXmkkKb8i
EvPGvZlrdK+0uhwEKu7QkCaveH31XJ8fXjczaf3JBmPPs4uMYFmFmSfIFSxO
z0w/MZA7f2LuLn+zvyL0wBrgwrhE57SLErbUEUInxM75KiXRGHMMQDOBz2Qb
YzFsQANX5u/gaNHszM7rTZLkphjtJbGg239TNj7X+w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
EjcNtQ+x66i8RmA9VAeTHUc+ABQWc2WE4j/3oSM0+qX9UxK3ZobXyMSFEDuz
Uc7L6s1tX3IHMpM3bSiS32OnJY4J2YFLxoy3dffKM6JhPgW7pm3T/XI5cyf9
S5Lt9MtyaHZCb0bTKxhj0G5Jwg0KQzx796t+UiqqjhxBtNKMZhI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KlU/NQMLw1IOVTgUVYuH2j3B1iRVfQW7gDVeopjc+9N9+/JuHxZW3EIV5/+d
/yDnsYeHDhotv703PAFOAoDwDhQmc/xcOhDjPvG8bnQ4cuXDnGvIiYHjmH7w
92So83BBhm9MpPqsQ6S9Ejq1BetyJ0cqbjRj9c0kvelEBpT9SoSRUPW4SQMo
Bz/XrSQAV8MjyZ2/XD3uXzqAHJW1fHqjPVK75ZhBgS+CSBW8ZpYPFTVyYlcs
vFi4xeX6aWgB+FbcT02AyloQAcpu/6GLD7Vukl7Vvw2VQuflvzBLM0NxmUer
SEWHmvHDwy2NIRRTiz37w/oFtQYUBbqNF5DSYisKNuGWWPNrPAECRTNaIWNq
u+PvK1IDWbtSV42hhPg1wQEuflM26OKPfKKvD0gFVlY4nblOkH4kQhQ+jbh5
EwfDNmv0uBJFldbC1XPEK+iezzYxtgHbfoFa1gUr4IRf34nrsoZhbqTI9ft7
yzEb4X1xklwMUtaKe43MCBwM5yMMxxaw


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
rTWnBQyb5yDxaQazhCCDamgPxB8X6++6ddMxB/5O0HLz9CadxNTwJNWbtYtI
Nm6Qzj4pi2cW4dvDmraxXfKni+nZgSTQAV556NtP3s+7qwUOMV/WugrSLvdi
i1wzEExyyBD/EhO8CH3CXIKIv/qlyIMxYRK5/BCyLSZwmiPQbCc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RYsAKTJ+78RES67vhUNLWowq5s+fynR3Lg3sXqNjCWip74WazOtDcMHi+YcP
y+x+Bq8w1DmNtk0nIqvtOkCZX3pEDnStcGGn6nWtGCRDAJOYVyREpA6C2Fmg
iokTC1Mlwmn0WiSiC+dhkrCROi9kmAxolit1zgoy8bXBjI8JaSw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 11104)
`pragma protect data_block
5+OQNmoanrlz9wxR3LhbBScrJhKy0VtoFFds2vKqSiJJvVbAqWFss5HIXotz
HH62fPzaildMHyHCeTnhiTXrC6rfZZsXiw6vWU0ZXKKajQCYqJlwa1YVPII8
v8skHjoFd1LU4jlOa1Iir1HrasCCD52kueNoK+clQdrC66qVBa7xCm4Ucr70
F9T6jNSJHT93ZZgdFZ4kuTrQsAkS2R+m7m5REeZ8w0ZCKuqgUQcHHeWTo4x2
wUWx0ewANGZGgFZhUG8byfFqcUo3yYUcVLYVa2cfdp1b/LiELUWmz7IGIWbR
WBFTmQ746Vfn1FcFlO4a8fuv2XnGlN8ci3YjJj3ulWdqIxxdTNHzDgGmcLMp
DrD26hRcpWyp4KQtmIfAMVpkGkSvSBgFp7vJxJ5USHK8WXDQDhj5EgmMSSvg
oxvn3EcoNeZWr3wzEd4Jasjx56HFXJePNTaTvgTCnwNiiWeO7QEcfFj+D3X1
6qTaYPN7ZM31kDnwCTySE3w91Q1UlSwlKGlP33XbxKch29u95V+/M9gsS46R
NyQL5j6X4Sa8GDFLSNjqtDCkl5Zp5DZ+X5RRvc7+4+LA1tHTjp0qwO4VgNkG
ciRNUC7GrerdaqAHnrljIbFiEmF6viZC3+fo+COD7G3MjrwK1CqXUDseODP8
U25famAMkE/Rwcfhbn7MkOiVj60pUf9MqVMGlgh4znZetAZjJHIAMI8vEY/t
zmInZRebG8DOcEZ5QNsnqo9doba4BTW4hHEY988Js3O/rM/0YaH5Aajz6XLt
Zs0L0gbkypktoRtlkLDyzh0BOV+LJws+D7exPATkR9ZENe1IXAzaFbgXqxZa
ARcXNn72z5EvQcnFem7Uag/KsRRQZ6ucVr19fdEApjvtx7fAgiZviIhXUOyi
Yw4ktISubB6acKgOSc4nodidEGK8yoMZgtsFU0o/nI52UUukhBAFzS4YZTD2
0Q7dCyqyNadjWQJ2lJfsexP+rTP4TvVohKaD1kBSVxBI5w2V9UR38jRGPj+E
RzfUKKioAUsb5ItWOOGsgzRvqCgknNwuDm5KmAqhxgDjpXg9aphh7PUIHtW2
dQ8Lh4/u83/cihrB/iG1L8qWvYTzM8hWm6+I9RBBLZYdzn8Y3L3u5X+FGQHG
/wUF0sCGCl7rKkCgktdWXGEcHliG3pT/d+Lnfr+rsby878rwfuDJHESD5lCk
QwaE3faW+F7zg0ZoXVXpYSHEQvl+OW3E+tUV6FwC2kDjW+FlOmaeb56t5v3m
nveiHeGrhqPhvUpj8Xpfmy9vU6W3Ld2WjHf4dCeJq0Rg757QLTN0Ev7eY2Va
8+8Lb3KzqaF42EswNUMluCJOgMn9sAukPX79rd4UNhmzY0m1YCbRekpTGdNb
jGHRB8h1iMb8PjqZ2TfTx34JYKSuOay2tLaEF6/Xs/NutgpqS0fue+kshxP4
LYpSyGByZDSsHrG/RoIV5ocP6iKx23KZPxJlMwqNC28E4Jr8ptKoOkmOx+Ug
ZdCjhHRCEPVaMou0Abvpn9AiALKR/+nr+KXg567QxedsaboEN2TM4LMycR4f
If6B1Odxo6zqBbtpmCkH0x26XDTEpmMhBlmyd7kbaCtn1Z9TQyUoigraa/GJ
QEUy3eS6U4QK/fregB5Qmf74iyC8fVTAFGZoaSPUbmjuf0R4Wo583YKAuuIr
PIYgmy5+Z4NkZMEXf7oh406AqorLiMCFJUvCAC04rs75mEIgbWI6Wy+jFyDQ
BcbHoeZzBV8H+uwjlRP7i9LNXseDqSA3TI7AlXz/PPK1YUBTY7TbPosM6z1W
4T7bOZEQMreRS5yE0nRnYK91sJybJiUYZH8lpzypg2dg9xAXq10ZFWhmV1ak
rPFw4o23mmOM5GKS6S/WocRb5iKnlk2rQvofC0YQ+1GM8e4nCvlmkBWzEcER
qDVDsjGkoFDXpq6m1xmTCI0lQUW3MVqElMjjD1YWzf/Brl8o5GRr2Cc9t3a9
AQJudCCDcTg6zOFV+HCLrcZ+9umdO9LqNVFqklbvHrapQxmoZEPNqt33Ayl3
hToTkpPwWfzdb9NlKU0ZFtciJBbVrmiiBA2Vcc8NzPmzYclrw5k0j2LZ8kqo
tfiw6wXI/j7epRR5cNRvMVWLD2b8vYyKJoAz5fHYtDMJVB/Zljmkqk3gw9Fl
8U8POMX8UIrGT6IzmUavrj0ecZ9JKnZfoFZQj2gGrplmKbuDlGMN/vQLlaIL
JlAQBTHSgdVe6J6MFcb1dlemy9hqVnKqIwu/33jFYyxUFF5+dMwHJBMeWV+8
r9/4o0lJKKj6Ir09ERAlirDxSIabPPabGMtgbBrcrpboGOiACWPEm9AxVQZa
YdMx6+nfDgtg7l5Li8uwCqNVd2q/ZEmrzC7rC+rNwyw8MpQtL2HjTn4b7TBk
/GNQj0QyiA+E7DRVVMQ7eQkaZEEG068qf9AhR8mTNNw5LDbnIsQl4HWthI2S
ASdQtm8LdW2YAga9oZe/zub9bjMA9U4wHyG0LrgH/ZOgdk8rm1JbG0rOeu6R
yKrqWd0vXKnM2QMFnu+MEljg362NtsHdrUrzyWdHQy2qOhWLc5zIwa41HEnP
4LiOW806jGRDc4NOF6XfR1iuqwO/gTXCcNyaUg/xXWcTMpNWHcUiEJS46z+b
fhvl8iQVuYT6ojDXttfXlP6IWAdmL3kTHdn/r95HedNhDC9D0g16+kZbdxUL
Of/ODa79NFUcyCdp83d7t538EuLcHldHjaqQgF+4/5JhdrNn9O7h2DSM0OuH
uHFIzS4JKzwSq9+VieLeiSWtywT8Y5uINzB1nBETnQ9ZAXF6V18rdkMsZbiw
Sjpb1cBdBoHIUcqQXvIWfNP7ohisKdWmxsAOi42uzjaChibEaBCfETnD7p4u
hRK81T7Ee/6JbRvYHUjcww7ofsCgLMDu/oyaZmYqKM6mloUjcAOoKUS8m+31
St4hwai0uJH/uVFsfaai14kOOiRHijCBjctB2o7BXjilLB0VamfWQB39DhSt
AD4sPYNV5YNVEdQbgM4/3BFD2z0TUMFpfL0m+hhzz/DeounC5+0jwP5xiT2U
91zbu+LNT/CQl1miXRUttaZnQ7YHKLe9N65O9ED+/Im67O5ogp9lTNssRk+c
V5hBxFUJIJIrxvL7P1OUNutnRX7M47/xH9sFVbZdw6f5uwRtnlfbNLt8yklR
AGRS/ewNPYhJjG2RGYjKOLMi0Bp1ZXnYGcyiA3OatUDrBE4ZvJLln48sF+PR
Zdy1FZ4KHwUyy8rsjMtI+gxuAT6hog8H7Cvy3RfOSSUgNTN3fZd7j9V424tC
6Wg8c2nuD3PtzJBwZrrOeCOR/nxfcXdrSP4bzvJr0rZS+77Sdpre/yQIiW33
MiJmQkbuiuiLDGQYoXTBf2a0xTs4gXSzd9EM7RbKFpprW3mTKyJT3xSczNEU
Is7mZl9EDq9gbpMM0clwsCPvMy66ZxUE4TNF6CGso+YgMMNskkK5sx872PUL
+EHptewyJ8eNjn0Dz2EICsp+KSNJp8Z+BSWLMwrYQnrh+9Pse5D34aZCCz37
PC/Sgfwbt8g1cISYt7ciaHpET06wxYFcV3luGYjeGgIDDyeGSzB2p5w3jPKp
haxtnE4v4HO1cMrznyIU8GoQM8TGuQW5b9+TFlhxfWAE7uEnLgqYA5Eg3hcG
3hAVXgBERGhctjjRukHk9tolR+WHSzHbqgTBd3CY6sXZeEzf6xfLhT65WQkj
8hfVedSQ2pErWqNbCrVnt9jESOT4zLNI141qkFRmG0RRZ6JcGxsjREGGPmqr
C+wuoBz7bs+Dxhp25b28KXaIF4RuV4AwGI4FnJBAGUzoew8OAq0cQ/1EjpHe
vMDDZXXBHI3Kt/gdaVfHeJr3Q/2HXdYE0KdbbWd2MFND2/ejRoGk2p2M2+YD
KBy8FXH+hZfL7zXi7qEpxHZAFVRV0BxL4wCv3ODVHGTZ1Vr/cSl+gV84w5n3
Bg0E3C1XofEoQuwbN+J7iYAsse0IBzP+io2Ua+w/80YEC1Oj3UUn6dH1NGHT
pbgoEf46WpLy1O+yw+GkYm3f120xZdFLBF8VJB5SBGd1GzJXAL+pQHpfXiyx
SAJnjYB003FNMS/aR2SXUquY6zNu8GvCQYYbDQ6uIIJpQOrlWQUgpL14jwRq
zFK1xGQRRd4X4Mm+jy9E75goVDnxYnK++nvWHgCNSG4hqTjBc8iWf9zK1VEO
KISPTl7aZQL+Nd9LHg9F08w5CcLJsspDdC0DCbYoGpYz1EPmZw5LxEC72+ft
+eihoDsZIeQWb7kkaYOsLCq5/BFRdLxRDgNwYR7uUmihpf8JVVPFdIeEAFBu
ur6e7LdZr0dK0BfmjQmS88npY357q5fAG4iyEqmSNY2n6LiID0pY1yVfZkie
cWlVvyyWUdUUU4cqioTRx1rv7PiWhw+RkwtCAfikIslG1N5d3/XwDHAoo0++
i06iYyc+1qtmfMYFwGYBS7mkWfvo8J9UBEtrLWLoesKdxHrpekXfmIDQV1nC
vBMgDVwm3Trxq4lgHSMzw2CeNM3V6Nh5o4xbhmQu3qIzeeAIxYuUoFIn1C9d
zRTvFWhrXV1dZ9TjbzANAZOL+5tBdjZjg4ES34PqTNM6VpanFoMu1JJRX9Ue
dN5K18+kEyCGKsUexb8rs02wEXQMEPVcVkZARRTQ0cwHkPiU/bqoxkpFo3Hu
Qtw308IN1nZ1mjwrXWvwSbIxy9+qSlybvx2Y0jnAU9onHAXOSPAccXN9zJHv
dEhb+YG2yJJg1MjNrqO/5vqWHj4WERJmNm1a+HxYclktUK83Nm7I4+mutKcC
OdQrN+4NReZNvcnlwn6TRXfJeD7MKj/3cdo0XYXKi3CbMe18QiTDMJkmCyB4
Udj5NKJfux0aDUzFsg1iJtGdP7psgGNxQpKZAz7Q7KL6hFOzTOxD4Rbt8lXM
WdYEQlTHL3wEffmVI/V+RbAVlM6K8LwSWW57Q1r6vBa5KLbAgw4xHMOSX0tK
+0tdCwSliBmCPmlLkQQoU9luqdEkvB/XHN8GUzGVUQlmMcmI+8A8ForhE67P
OMx7gT/CvBcB4+olku5mXtLyOpTnjKO4GDS9UQWgz1YcQso1SRI3sHnBPWDj
zJNaGlnjztekBc8qWYV22ceAMCAlJnU09wEZz5yN4XyfhzuQc/4FN67Reg4Z
99qT6oNl77hHvSjGNXvhjrNOs4bmjZ8Zs/6j9PWGcXqfDkb08JNEpF0wFRPT
9EJZi2X0idZo/l1VPhf2bRE4WKi4bwGPrYaesq9cMHxzXCNRzZgeULI2SsBV
zf2tQA4fhMDPdJZRm9xDsyHTysLaCsOlBWlIkhjAQRBeAZRHm2wJvSg0hVbi
g/e5/DmW3slCFuZ5Olw0oxHW6lGqcWAChvVs/UZ6n/Q/9sBu4OpDp5MC6meS
uo9GIu1P0oeO/2bBaHTVj0h0jm7dVXDL5omY7AlBLkfgoIt+mwtQMl52MWTS
X94N1nxsnoZieA+x+r1SOWOt00uYqKa/XmoO7k2bTdp/lPhoHX8W+mhYuOWl
yy3ydXkbBCFkOpHjMF4BAi1qeC4S4yOyo5/BlLCd+V6EA8mH+ZFUCGFOKFwG
uwdJD20dil9ywAftVlBPQk4xTXuTfae1d4zbIICnVz5M8C2lTX3rRvsmF4Pv
G3LfTYIpy7sz+7tvJ+OCmvar+9QN86cQ+FYAojAQXxOupf/WSUqTJP+P/GIl
sz8nhrDmNayYR89z37N9ai4U5rQu++G9RUKIEswXo8oOunilZV06HDygSrzq
N0Lwg1mblVplbOcQ91qjXqZprPxdjmxIJeP53GbaTaGGCMz2ZdqSJnE/fAnf
M9gRxrN4X4e77Qpy9TYJv+no2/sXiXPcOiL/t/3+DDU4t7S49p/Y7ckDG5a0
7/RPss6h0dqccy9HRAswVPBn8++Rtb9mDeV5Oia94ZM9Jv7H+Dts3FmM8pIr
D8Bzve0FVxrBCHSBFH4k+WOEY/u+Z8hDIMmmEPEBMjD6rzbQhs52R9SvC9Jp
wTUIJ3HYHVyGm8+KG23ZLdrffB/V5YRhJ/ara+Lr8Rug7fS/Jv4OXI9APH+R
a7Qa54+qFSPpqBkoXU2olGKNtLPzJkRFLNamo1yNjbnfODH+eDE2i3NIXnGd
9iZ+cW9YdviEHw4lTv/9xUFgZgWWI6hFPl2YxDOcVHh20oiFnmEBlxpnP6kN
2MIjBaYsyBsli0eczrPqCFnPDjeSBhRGXHU+sUn3t30E8cgCYk6kPFJ+C6EY
+Z/JKRXNGGcHnXYz/iMA8zYvIyqW0BdwvJjthMtS5a1RkOOKDv7giPI4SH5W
CR3X2JwECylkZrjvRmg9nt2pMU9+swybuxjFFhcNz0/pCM7in5L98yW50XuJ
Wcx2IgEjsv5ebyYeiieOMvRFqu2NbUlwwkHGmFpWLtCDNR3HlQOHyL2dkicG
VDCNTSttZTsK724EjosMimEPnFTDNou3aFAHBPvuNvz+HpvWU1ANTr9+M6tM
RUtu+cTc1oiDlmJ3F+WA4ELX9ZAq76Phxy8UAAn6jXbb6y5E0FIicZoQtrUe
cVu+4zSAjTtHDUDZs8IFbgGeLu6EnyOqg0mYe0eKctr/zmY0iCtiR1pDn2kj
b+JByn21V3bMG0wTly+D86XG1wKsOJJcu6wwrKnGCOEiTrR/w3oZuEhmjEdf
L2zgJNLV8ssTwGRD8K0SrGLVM8foG4DMCurm/Nxt/gy6f1MqcDXUR0MuM4sC
sUCbJn6GMkuAynC0BXnCGHWl9q8SV/mhK0EV+YmuTg7xpHZUQJRuj48H8rT4
BJIoB1eZEqMSrWF9DQkMTaVn8H9D8wyaO77NZnVC2R/0fbdBFLzydvvrbIlb
Ac+iP0yuRMXtgjNxOiGxK3BlsQk1JcbCv1lzTnZaHsrQ3nFDATZU2UhTzLxt
haqYTJW63FW+pGGJlObSI1I1ZWXCFwbP5+/tvQoENq8EM7pi4xa9oMhWp8LY
+jFWU41Dvu3CdwUFXwKnyycbEqMapPf22/bgTAfx44sLqrpOKOvZQl0OEen5
UprlwNwfbS24K/X0IUKT+VG9Ksue2HdbYO6qeiYNw8uU5cfMfRP5W+HFombC
dP4A4RJh3iNcIG9Amjo5wh75/6E1NgAAGpS1UJueMIWA9PBINS1sGyeKjF7F
SXkFsH06KFjZnDLC8JQIyrvBNx4n5iCZk/IMDAdQerduE+oAXysqBJqGZxt3
DFLZFQ+w/qJY++IWDkh+4H3V4J+EZuRIXGEKrrlttb+JZR5IIclPPrR8aau9
hBeeCRPrRWkEe0Iemo/VtexxFqfUvokJJWlc7tTIAMwjdvKQloS1Uf5vBiCX
c94oP+4b0eMp+0XQRMsZJQLOq4kEAl/mgOLURTa/R8RZAATnMMHeW9rTpyrg
I3kKFs86QjKhsmuvQhBSuzs66WUQsL4ak/Eymd6BB+r4iFE047PvOxfBsHVg
KWdqNuR8mZiUhHZGJa59o7Q27uztpGFQp/CygHRidWZW3oP866ZXliR/wtVM
tG3SEhUX9ZBdAEiYgEp4zVx3LVamPvGo7dpcdTqXd7h9Rx9NnMJSggiLBbuk
9ZFagqfmNAX5F//1bXTCJyC1lWV2EZAASgjJgXkuzTtkoEKdrSuXG/XT88lM
h6ese1u1bupT+MMPSfU9r1C99PCyWo85DfrPhSDAgZOR7EBv84rMwfy+mIg+
Av2v536oWoDyKu6bnapgZT92+k1I+XTDbR3xQGg0MeXBlfKsLyqErT2qBnAC
J4DV6TcHxeBo3rIWa0PhxUImuRsKaq16wx8QpanfKhJu2SmC1OoIwtRozjtY
zGv+jYg52pEChRsroshUWy1pNVdgFKmWy/JYOxDF2OLFSuHBhV7czjtkAZiM
WaYrPvJfxpjxwgMRRIc4urrdWgp9rFhXY/iwXdTNuYVwKzwR4uicPTecRfRX
xmJJLe0MdM3V82mzQZxgbR1wUuxZTehABl3G4F/DbP7dTY44QlfMFRRJsArD
qCw5J9XG8hJ8iKrt3Bb+hazISu5LNm4Irmjg9BclgEBwmaM/7WHL5NZ5DwKw
/gTXV3ZBLnxVyuDkOSQS2cjBeStalkMGI8vXKEwMOJFfe7gIEEnG7OPpsCAt
5W5son7IUkHk0j9xfwgTX88mEp03WWFg0utkxmRgDsJQpSb9QiTTVzkau0ys
V9/6g43Wekm1NNki+8+8fVH/48ONGT96wqM3O28V1hv5Mgbz5NeL0a51uOzg
bQ/vkO6TyT251IUK/P4bNgFTgeQpkrh+wTE8KrH5eLd0nZnfKqVAkyctyA8h
yvhZTmeL/tccLj0/nw9WnfMLJ9Ls/5ykUP+ZfOWPbngxxHDaLbQNyX67xDeh
Yw89pG4j7xIohTcyRvbsfIEDsE3ivckYWNhpgLKz8R0kqFSWg4u63Kz2587m
ZJrGrg9BIZu9GJpmliZjI5MWY5XjFHvo7FU1wL51fqw/DgTKtQN8lmUgcer+
+y6TOP3DU0krSXQylrs8CjNGB9CAOgeeWMPFKuMwaW2zqiFjHAvqEsXEu4Eo
ZFR0rN974tcW5lhiEHvAjOjOC0xzfxSYgMihU6vBlKLUU0Ac14InDjGO2t27
7PZPRZobtEhq4SJHoTqsEaPWy6IY/FQTBGoDB4u7IwHIarp6ltsoQ6Tuoa5V
xgXQM6Cr8qSbbfCRkJa9P7+z1b5JYR5KShnnVVHqggP+getUmd1E6StsrWRC
6F7juYqh6UYnTGG9J0/CdxbVqvQU8J0L2MgrPo0I9eV98ay5MwUsM+7ATzmL
7YIOMYOO6sO8qo/yOrj5diBP7OhhyZdyK4ndNU0x0vsJRmA24f4ZFYFenlJ3
yJeb3RytPEL82ovWoCNA3c0sfMnvmi8iYkW6Ve3aCfxSQ7UDzDaovMwp76WP
SIjh1uoh89M89PXs3XGhQ0PE9v0GLgqoKLmzuvxGOs71xWaCwNoEohcvOecd
EB4s1qApePtPm7XomMFNEz55OwGsjrjnxVXjj2IixkXby169twWx8rXXJGqv
uucmuORZw2z+hAeispaUtaoJd/o+e9RnJmGgMzUrEPgwy+Ad41yIykmKv7Uw
6fAP3JekJiEQLNHL1rAIsAz+V5JqyrBXhtNJzNtvks8QuY42kPSQREP26dcT
S8e7sOe9GA4SaY4sLnLYCU+Zks/UHI6cA8FCBFev1sTrGXs2RPnlSuWunHzU
0QRWrOP3Wkmx7hHAp8cg8O38cZ3vkF33HtoICMt1voCPYoL0Z1Wj71KPV2Q8
Z/0zBmJRXZT73hxitaXKrd33pMV2y1mwX2sya59DnoRjk+UaCkRZm7887ZSZ
jQOnDU05Z7bVDQld2Fzj8GYhSSraVwe9vyrGAW3+7NXVtmO9q1U2hw5Es0eU
kbfEnouaW/cXHmqN+bfYePG3wyKllVV2F5JBs/y7sadh6oxV9wKzQmp5MD1n
JyuJEjyotsrV93XUetcfZJJyLwPZmPz0hSXHiakbhq0sDsmVeVXITDDrwXJC
cyImvS5+buVYRxUNUMwXb7QKMuT8BDBb5NaL7SStMQmx4EP/p/JfQSezFXWi
DTg9nseKM9HKfCQql+Rc6a8GqcQaDDhXuw9T5U+6ygNmy/JRBbzW9v7KP/Nk
DpWRy19am9jxDnwiCywwjaL+cbMwRRDa01jp/vayZt/Si5mo+1vj7h5SUKvo
7fZKTn0RGEhUasFHomL6Js49qoSx7GZ6W4Pg56B6DjM6dgtNXUA5ON6hEwtJ
JGXn1yc2xN6B6zqRkLc3KH3sws+vp7jIrVyBRhIeRdwwOuzzfna1DPZ/gDGE
2Mxr892/A2MQybXtHkQCYxNz78I8ylZLTiGK9bMTdUUx/peCXEHX7nvXz2bT
+dtaXyJT8YrCki0njQq2+AB97WLTDJMj2zfnBZmJ7en+12F7nDn0ddJU3hcq
erIqzui8IXbrfyppzFtb+b23CSJvwygWOLK3FNcZsNzlG4v06dUqrD96xgxP
A1o7aNGeUlG37iZQ7AQgsTqXRrXroPhXB5JOLpichJroODOK5KlVUYUNNBpZ
g8U2/FBTQUg8Rg8KixgDcfJTF7XtoniScizKWkALnkeFc3MO8/2DR8tOz1FS
Drr6Uu2xyVa/hpZBxEu+d7eqR9nKXihsCDsAbNT/ItB9VnX1zQhEBRPC+ezS
3PfPLq29iKgDC7brxq3lLg7H7zuDPsN+tFZkhPeOvjLJLBWubccyPRnHdPRO
16hlWWaVVaAXL8YWICRGnGMpLjJC4iny8g+2y4+0oR8bA8AAlEll5kFiSep2
EmVoodkf2hFp67I24nhlzy3qz/hQAJ2utv6jugNmGhSu8E1LpEorBsuUODDp
dwKfWKnpjcHy5fhUXV8ks3oyQ/tZhLL77IhjMqMW+JdUEEEeheCWxVlf3Ljf
gGDu5dD1wZUcHR/EsUO5JH7aAOBO6nIKJOCpR7lfCC3iAmYRJ8CArKZIEGpK
mdbS31ZGs3zZtxCZoAS89bjZWGaaC5+vuh5b6ZQ46wsNkvYaSeK7HrpWe8/o
cq966zL5ELQWisPe/X5e6UAYlvTcg6DQcTYXuH+GiWvjbEuIzOEeR2wC7b8F
bADKqvFZBz5VHAqCsqzja/JpCVB6V0A2zFUWPyLyNeQJqoq8kUBUTLxJhpTs
Ges/MuwjIdaFcwGycz5vJ/90rm7h886jFsbUU3WTd44oxCQpm85tCullROY5
Rtdl/zy7SJBNqXKQW31XyiPWklBxtCIyR5vSsQ9m/DszMkpDmFa31aCJ6bbK
1cBHmcn6xNHuR6Q4JD8gyBdZCY3kKcxr+I1RgMLARupUexSW5vrPcLrw2Ngu
2wru/vmoXoBTyfuPKUAOiI9+TYau05JJcQwYgk1BwnqYn+jeDX7/Cez5h9Ac
k+tWXBu6LCyWDNfYWMuweZTYTTg6hwckgX9GgJuyn0nQHYXIbGNMsmPmGL0e
MSwlSeofot8ZAeScYwG5TZrJjPompE8uYM/eU3St/kEy6Jz5Q5Bap0mtH1yT
oVNerT//fiX6iOSfhOWcz2utkue5mDkbBGGdIAqnzuTDg+QtcKLc2Kkkw8l5
F+RuhoVZxOde1mykWSYaGWDuGy5DVBCEa7XXK6j1pDM0+OeXzBcpTUHs4qnL
BjRfReOAqQp0LG2JNJjQGZ0IW/33aoNT1Pv/CZzi2pnbuKfPRyeWfIj3UYym
sNKVKNLbPJppwwqaNgbirMcWuSsnucJiloLdef3lIcicX5+4w1lWE2G774C6
bs+P6NSK3ROIdhkpMy4ZCLDwXf9Qs+A5T9AlFcm4srwpnoPiMl0donar2iHg
yt7zZxEPxOyrXgQw6nBE7BRzNN2H4zaFvhZjc9Rxk5ipzR5lrIwstBYYGFYv
ETUVirc0l0ct2pKGfEDI7Jbo+xIxww5yLTAZC10HRDBxqNQpgJhIa5l8cC7L
aZ2BB+HIErdQDEWyyJz8ZHmSK9aNQIi0NJgrlXcfS7r59mjtp46osS8mU2wD
T4YPkSebz1yfxQPrbItGnzpvF2JHqU48PpRRgjOHQuvNt+eXAHVbSxQ5xMxl
R3ouQDFVvQ0p8y3RoSiTBUh23j84du830jnR/4sPmXEnzjQsdARTuHLYezAP
lVDzQl4Z4pH8Kn6jMf+AE/x70rBRn3lF/182d1tymu9W/zXT6KuA27jNmKzG
H+is3t/kJ8LG+gRFbPHzzKdKTKVN9zIln1n03cqNFbd6pBoKVrBqJjOFrKMw
+kpsSCKlifUYHRLBqUXMc4eYG8gGJq4uOHxLRFq6gd5K6nfoamPEH5adBpUb
z1BR7ZS2834vz2XoQuN8faSaB6RSBQJiyma9poX34ckPlRPNZhtq7KdSFYgk
jHFlYIN91bHtq2/mFppvm5FVfOGUEPixd/ntPGWKE6n5GqUAJACVVgAr5r5c
sbVFXU5hehGfKmBxmwq6L8FjFxXGmi5EvbW1wMqZXEdFM42Ojr9295KYuc7S
mTM84BgoQRO5IL8xvccdKMdTwt2m6J8YaNaJGyA9B7tSwvgfF8Z3kXG6DgGl
73xTlMjKZcM8RkKMJEkiGUpN+BibTmRVn1hvTYcz5uYwQzg2Imxge7AME6Lv
O4cRIP2Qnq0ANv6nnYkYiYCJHQf1OwM1T5Y6FOAZUo247LY2slYdH34souBr
wwXYCmDpP3k8+cWlUuTwrHVIw/rQ4qQebmJ1jYLCJipOhS76TJRCZXxqQhZq
erVUue6tlAMh4Bh30Lw2H4zIl4w6Z0TINSvVqL0P1XDRz9ms4H/nzuASBGKY
t3O2uWByT09M2ABkL9TQqufLfFqLAt8/+eL7m4EL3DZEPKYvOpzZ5kv8EVPF
yA9crkp4vcs/U95g7hczt+1a9TGyOdP7NLTcGxS6QqV93LTVqSxrkmvwzCSN
h2p2KXP/sL6MJSKtNwiEkVTyAYbXl2p/UUIUGg0v5HNU5RczJmnuZsJyI6Ol
at4aduYSBq1FBfqC9m9cynAQ4bnFsPKmr8mXpvxZxYE2nYX/pCwkL96WPvHp
6o/jiFfpwub1eq+H5MRqTSsEyy4S9g5jWuTBhymGX0oAse1tbwng30uJLqqC
5k4uFR5xCQfEGLESf/+uHCobUkKP93M3lLlxxnBYWo7ETPBrVdULH9aWZBs2
XKGVTPOcYYRWejngBRYz6Bgfr2ug6fVc3idHjCNkZzum8MKxbSvK556+Qp/V
f5kLrkTBofI47F3AEPlck3dpywXjUKtQ7TaT9W+InSIZCuOEoYHRRLtDUYvD
fev4sWNaMcoVaHhAQVJMLW7YP7NXWPqLtiBOYRVNbtdLBiI0RaNE1u4kFoRm
c6JICRpryTexXWHOxzC/8G6/rXDhZyFPKjMv4x0Rm13phzgeAuphSOLLGvZA
vMaYo1ooAS11d9Kvua7Fta0aaSAwTm8t5U1+AyIxdZ61ztmoBSD8yI6Umesx
BZBpWIs5sam/njWXzVuMLBEHmGdbKrC6TjJB4mbngCPMCsoIhezZW9fhOrNZ
WxIRlRwbFuw4Yx83wKZV9b/1GQvoN1QQqx7AtWDj9f03qD6gLu64Y0IVreOm
Dd1fjrXKrkzZnGATWjzlnY5Q4xx/s2/TF4xKlbcToPks5KHojYnwe5ZY3IQd
JFrctkQ3qh7KncZ/ugW6YOxePfnu4N7cMwi10IJwDkoowMScMQsLuKS2jHOz
1JKj41lnSIAlKtiMKgdJjbTOx7BdcaApDvX7tACjHR8qAHYRFCNsePy9jPDX
gwyrVeaa6jjE1KnlKjg+EssdOCqxw/aNZZJSqldTRSwJuq0y8Wmlui4r7t2y
slS3gWrRtUz/URR3pMorz7ougEFGFztS8WkLBxIV3vBR+Lxp3joKvgsKXaZR
uCwHug0pUqVgPFju5uGzWkPuRVNbYzGY0DX0lWGi1iRTt1foOr+GqbBSB4Ia
z67XGUXdSxu4i2U3D1yhb+k1lO3EopKZ9ok3VbCXOg6r0Y4KaWsFGi7gS4Eq
t0MyiGHqOXdpMTGx3zjjuRXxd0zpA2bx+RSg+Iu20LPSsJr8jPDkn3/hKFN0
SJwylGs3KETSwkYznRdiedNYajxq24zp5aBrL3cIt+J/Jw0omddJQTwkuAqp
I+s7SThxH21PpkK6aylaVKPdsws/N3kTPeN97XdwB+ozcX2yKYVXtzhQKU5v
4TJW7i0ZkBV9Odw6RYcXDjEfrdEdDW8+qY85EnTVO1zzVfsg2O0CngdMKCuz
LJJEEYt/9vqrSqVHGyEghqUuP7YccR+meTmkm6JsL8Kadv23U42iHUYjNtku
zuRiC1MAwwccdt/3EdrAqRSAMJB2vHRZNR8ppKel/Kdn36RYSHQBo3egaO5E
09lRI5T/Tp86EFR6xj0sxK5UaNQKFq5KIyXpF9x31o6Wc4/XfpZs0rsPTms3
qXmywvYf3pOiXiJ9UAusXTIYcO/aZzVGEB9MUjHZksvFJOyao8BpN7P4KZ2r
38+S9xxQX3haQ4bxFbVqJiPdVdx7q5lhJvn7DQLT/MslL5mBrb/6sbFqTkps
gDUykvVmx2mSgbw2IjT483Ne+e5bZyn815jpikLZi2lngmoAQmficpx6/7b8
9PVa3ENL6nOtRo/u5470vYqT0MnyOLygXjfa7lqNTaU4Xrdi2EGeWXRQtPaN
unrtZzULDUS5ZJ9WIsNRpWkns0uARFfXr9SBV0NzNn6NVa1IDxoiqQudH5hv
xsJHA8fmydZiB1zvMizrvLPZjfRnUxEqwlFkWcQoFemJ1HXUKF+yWKEsoHHz
/ZMu6ukop4j8jmiTwpKQfp5bZdg9MXX6Ylp/jiK0xfe0QqRBRnbGRVqUax8g
TBkmDw1ddcykbCc6o9Hz7quRpXTY/P3cOlLVVpXM2TZSnfpcKYCVk8D+E/OM
QlFDiD2KQGeIOKtCMe9pq3dSuJIPhHdv75qzc7I4PfjG98brkMJOnQog7jMQ
DL6NDfbWnpgp5UMoXF0GCMN1XQaY6WgENV+0m1BanYh3Zbl6HT52wvsNTLLv
rZYioHzjjb3/2GLYEr44McE3SBuvcCOEgY3obr0qkyfIny5RQefCzuX4cjvS
n5gSbcezGFXyJCf/+RVW27Cy6lyLmm73JwxXKPH2uwiGWaG8yrI9GO/YCiEj
lyHsOmbkGYlbOwPPQkrRnAQNzHnSfl6Gekbmp/xhVx0CWMwtJhOxmirzrNJ0
AElmpU0BPXegkogDSX2JcUowbAxlbHG3j745WwlFWfPVRlLzNp9CIFoB9ut1
b+TgZhSKpGuKVLrHRBom8+4gTxPnIDZaPY1RyBuWYAOTTHeqhUSrfZM2dMY7
ckuAmq3JrT7cyULLUmq/SHF+QGMgzB9BWHcJJ2JDf1vLIA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfQBBBEvxQ+KiBV84xpM7wlX0lKE1Yunx/iLDr6k2aPyF1b81+6PGNQf3pujIbxRcYox+HE5YqOOMxgZEC0NWzPhgPXOKqthilOf6eRFTSlDXCWpsZQPCZD91++bCXyZTcX2UsmSBFbiJuTXLI1FjUoy8xogh7rhjivlCpU3FeuHUDmXo5gg9JrvtzP+JU/uO4VxkCQ9Z+szEOtcqXCTnW1IOf0BM9rW09h65bMxd2tLMqIkK6P/p9IhNROWufQ9iW31VwqfoNt5pmGu/ogXBDmPwaPUM4vqvc0xBQTX86bbXu47tafZGHgovQKRbfXumWlX4Jhg6RCIqC7sHbCZtYYAX1utQ03s1qOxMADvHAhaT15cgUmWqeTenmy2cXy8Z/pg1NMOVHqZ8Ol41m2/tF1EC4MSN8tMn8etpDLuPAL2j34HaQKsKOkTuDYKzDdQjYQaLCnUBKENvGQ2RRmozOAcq/awdb28iya6cG+9Owuz3AX1Ql4p6VIiVV9pW5Qv9uNvSXPyq5GYyrhydHayECrhJuFt82ZcGDFPQ5GLeD4ck8da285W+Taq12WZe5yPty3nCXhH60pPGXriZU7HgPHLmq9zkjkmW9Ej/234ZAiypxuyZyx4P5Tc+1gothgi8HxXbp8I4tdtGsN4NotU3R26gDi3kNipPX5PUnONpdNl4Iwo6tx7fj6pUT2mIFT8DbHJDMA77v0TW6UwIQc+76Auoo2ht22rqaGwOTUqIJsIcQS1zm+gg3oylWGHLTWOEOZhRyZkCZsISQxic8rpeTr3"
`endif