// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
zemIglLocLIUAdOLXvGgHFMEW+1EykObrnGW1kU9sLuoJWYYOPXpFo7J95g9
bhKqdiU0DRCqVqZqahkMpCpo4PHEO+0jWfPMI6am84L4G+zHPOakg1J4Cy9r
/km3mxwiDNETjB1h5bdJSzn7pr21IssDUdGR82R5PPQyCrb6USmAiXu2zIcl
UVs+MxP7XX0ainxDBrpInsLP75O5yTRUGHY8d8Jy6lhskFTSHrB82F6c97tN
/EG3b9corc0/A0vgNcxA11t1NQzk7irO2ni6pou9ZeXmEqA6wimEyQQ0HQpX
aFwljqwyYMFBVjjfGUqPoJxrWZflYktI42sNEaspJA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
S6a4WDNePmFY+ujSfv3k5jvgLPTlsPN3TlUmvsD83i8EyOyZuCXsqsRrx+EK
ow8DqV+otW6KSBJPreCMs8Wf52m9569FRrx4FY2/ZgFpo5bxlzvC+O4wde3g
vUDaAUnolX+F4MuNYSgv+Qa2lrgGHBtWG5f524d1g2nk4zPnj+FWltlT2WnU
pg+kzAPtbmCOlViUwSZHb4KmBMZtn8eYiJtdL5qTXQ/HOELGfAh25gID6utr
AH7wHfiIFSB+cm5EnyDWNIjadCXT/kU/YC491mOAOj+rIhjNxQcLzYsbEp75
N9ZNOfdzVaKC0GcjFbEt6JJ7V5QjdoaZUEVOQzai8Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
H0Ruzn61pw7+PS+xib/BUKmyuhYXkdiMhYOOkEriJsbHDyhgFUZ7pgOvYFQ2
/AqTrML93i10d+2k6NsRfZzisTHDTxS6LLZqQbMxlD8TcQPKZoQouQQhDVQ+
QHOSTY0YmjHfb0PgKYViRd3VD8d+i2WJexWXnTRzJNqvpIqio8JdGsHidYvX
dUSMpb7Hsp+OxIdGeZPbQ4q9bX9qQzYDF6somm6JDeUgCMzSPI9Q9wuZKfQe
LJCq9M49bp72iqBTXklIVRoPVPsGCZzIr6yTeCKvWInsKBQKdQ/dwAWYaWZ3
nSGx4ZJ9JSWJGsz+feqDRcyE++XBhqqXbo3vWIlNvw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Fg9kskbGRorXQ+XOFDjWuulFNf8XgxRoRHXbLVdYy/YO6Zj7T9e3REzUlP5K
ECYLnl0FeOaVanxyyPeeTBDJeuo3cf5sQ5qBhJLPGNI4Ggxc82Tw5vffzWQA
atOxetm6szoUkY+U4qu7g5MZRLNNy/eDtChkQPayJKhiO+kkYNc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
krFDa7ng823cAIryoRIBCJZ6crfW0b0Mbv8z85j9w4WOpKMTh3rXitxcMUzv
7CHhjETUNoHBB24DrkJte1GvUbBZrbfW/qAR+a+7N3DI3EsrgUGDj38sJy8I
Wzy9nkoUImmL1Is92UepdomvqYtc8HZbRejVEQpMv87fffsZG7lJPSLhHg7U
n49gYHbMO00Bf6QG9xYwX0j9vc0Sh1MAZCWDY6e2FMCaV1bomXlSKvLN3GPI
LbESObU+7UKoTkxv0eX5+O3dyt9/fDuCzPzZ0M9zHr8T35SuLGfohLi+3omJ
6Fy5AIezbKenBZp/T8Lw93ZkSU/Ov4hVmR4ExFZoewnnKexkU5XoCLaqSdQO
uUHO5s+TGHF8LyKoOm7zPAcjEvDgajDEgkZbFUfo2GAjKXvMLi92g8pXrh2F
I6md4QW12hfw6Q8uBVCyUWKmss1gQjX1iq451yGYGHKAuZzgcVJG2qlznP5Z
1OU+1da4BEHBOqi3USS8Jz/xIKIOdagQ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dDdQAGwlqdaXYyIJMoHS3OcM/fGxRNM7apdGwi+tHB1sE2BOYpzb25kbLZvU
u0rIL6EpeDJm/7nGcekexXZAqjsy7bWH1BddE92mOKpBAbLzahvip8Chil0K
QOXmt5r6SF9iHnkV3uiLKeVMmmM2y7T7CNCHyxg5wRE7VgK/rDs=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
WYyO6UgQnf4cWz1q4tqglMw54Kd6938D/r5Q2cbAC2D1S4A38S5YM9JYL5T4
4rDE9py8Ptq7/rs3wz9qtUmrPmnMc+jVrOVIdpWUtDhdB7+gkUXZl5xS4nKj
BHTc2V6mVTCtYAKWbDHRTQD3pn9FhRe8Te/BcGwM75sQy3a28kw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26432)
`pragma protect data_block
/ezYh5Opwer9oDbuvenkroncekilgWMQ6nWQQtxNKYrRyhPReJV3JB4yIdbD
dUIMxJOm8ilVgNQnTDlzW9cuEXINJRuHQZ9+JcIKqr4RXPmrt+W5++kQRFUP
3GUqIaaBk5wzU33c78ukrNOqS2sb1EqCGXSKhmwqzn1ndd1THVZHI9alGTor
FRYCZib7yt1OcfiKX4k8+Aq20ZKbF/la2m1Q6CzSPRN3noasFZWxbgPbVL6V
GiMOGY1AQRIdMbZKizJyh/yhWYKgNctpHe+IfYqNCYQm4u5eaqyOVIev6ykw
IU9V/zfHUJWxmiFuPqOU41zJf3pO7ixmykiEX+U4+q7IkYK3GAKW3pwto5lV
ldtwjFrMHUVAeBn9jBVe75JgXCSlfMo7FHYML0fEy4WIYBeDw2IedJ0AfFx5
O5yzNnQ/dm2gZdtdCr7NL60KbZVcUJ3GbmKjxLzgNqLGdluW8Egffnw0r1vb
hUjEmXWRPZ685VvBz0kKzBtvULdwHsdS9Pqlj6m2+dIhCyKPCHb8gZYGuuUJ
t5haxHRq3OIZH5iLZPufZkYItiiqj39mTY3qZPTOyUQFoxZAyM0ZQzvBAA/o
hNwhNye/Th+v1WFAkZ5yI2PzX6SpjycZcUfFKeWVfn3Jpfr2QJp+Y9R9mVe/
eVRfnwkr5Y79ii9E7zc42EmF09daFO/swe2r8GfSrE0gYXNgzyDrGTfU8Sta
dpXTT4p03Vg236pr0aSDY3xEYcuIWnfGxGeaD5Hw/pafTWF86wL4xQmTqLEg
DUfrMM6loPMjeHAPnTmg9ZErrmvTyk7ZH8MX/uKgsZjKglkZpEhHhaurD+0d
Sun8U+iKRSzUTk5pNK5PF7Dwm71bk9NX+owyryjvNZXX/QyoaHclBJ5MGLMq
fsfmkc25aRyqjg6i9C+vzkYILBNQEBDj2AHmFwYLNwPBDIuZlbbmtMnRQhZU
dxUgvF5vbF2HhK/wdNQlIkQzvwGmcs6HcGi70einVdvtAMLl7yWd4LPyGOES
wHDMBuAbmwG5B8usnMtSlZDoGuZYakTdeMd0pZwHK1nKPZjK9dVKKjGh0LrX
pyVswQnC+UQKMkK7PVv2mvABKjEmyR53Ya7/Jg6p94EwgL93ahZtpfHmwcyF
5+cqk52SrL4unfI3i5nO21kkwVhYfaqy8pbV05m6+5pV9VzWyQyWppLv3S7s
f91gQ5kCDAEeWeqwPIAMyvH45f/90AxTt+KGBZbaQh5LlzuiRKsiKJ4UYvHY
RGCN4ADlXnoM85Y9VHGLA9dio98RXVjLUKi0cqpoNRWcZ5o/514/Q7yVbdrk
fb0ex4WX0NKOWnMON214qeNLaARL4OgX1Ocids0h3vgtw/8EeQEFgvH5jAZt
HKwXyojku/hmFi1o3qD/OOEVcj4Vo0eFLrHPTux3MLNf91Qlm+CoZqm8uPj/
6CdfUfeRNbEp14bVn/IRFeTNQrNtYj3d9jGjVNKJUGOn6lZYAhovrTe22tax
mdjsh9virMbQGLYXVV++pZ9yJfSZH2tgaWFKKK8RVIVEmezEaSxrzHnm1BJg
szm9pOgwRxXi8Jh+Kl5p8apFGRlDNVrj2aAZaQLlZypSteJLGnwY+HpbYIf/
N43Rv6wAquAXDW2IM8wbEzO/Lu5Pr2//NHmJYBaU6j2JOrWafLccdQhbpBD6
VVbLLIejjCazOwDgNPuZ4DxFSeI0v6iuz7M7qU+2Y0rMY2izgO3bFmoFoktq
RvC4SowBp+2pLDUKPXoNkvbTXtFIq4tLQOJfVRqUvek95ee/TdcY/Q1LfBCy
rtkztiTSN4Jp2XPv07iKdwCvD0ZRkhXRcO+69o5S40TIVC33UuI+1fUUyk/x
6SBBVgfJGb1bWwhAAlh4AtNurm2x5JoAYOqIanzN93qWugI4bjz5Ijol7tFg
3+A9+4otBLCixAcUtmBJEzAw86dgdDhFOwnUrPZl8WoS73jH3z/xCJ008M2p
o1RzAjoqwDEwt4ZoSIeDT6C/28RkZxDDZ8CvQ42jfCwcYjhxz8gy/40oPBZV
6K6NrCudXIXKH8dNb9fCSoux9NwxSqGOKualc642m7t/rWSbNDS9WHsDrIQb
MJEFW59IB5vwL3HAIGeDzLCkxVEDUNqnwLaZzLtQYcEEgzlgYJblXwk19d/U
4thIIut/di5e1gE1yjfdQkoZk0kEWt6jFDgIv6nRPnhIui8h743u//mYc2jd
uXauyi9i5NwZNVKw0Sz3kLe6BNYbsGDa0YcLXsxceE6wOo0xbhIoUsE8u+TV
DYwX1dkrFVD2OpWozUeFZcd2zku2qWR4b/7vMQnj+m72l/i8gy8AwD4YSPHe
YIz4+Ez5kDy+vGlabA2yVraaeev4sX/JWjbUKxoIxUdCdGcrSvgHSsmCj4Tm
6/CtgDfWbM9eV5cl+sBP0ChA0ziKZzTzPxbp2lbo2t5IYe+oeybVeUceTVIq
uXPPnbfOgIbxsn3uhJB1IuT4aSc6VI3HUhHthcNFxnNc0zGE+hE/iK1dtx0F
9furfEpGbzH0eK6dzaNFqGHIo51QN7umAzgKLYDaPIZgm9Vbx9/8QK/56JBj
Q4U1dL9ZSAxLtbk68xsF2JvmonWmsCWGjV7/IzjeWFG7/N2aVtP6fV/AgDWT
vbImYPQ0+dm3YABf4wlU48wRyQ2kSDyuXZ1FitBY1MWzGplO0OkbR0raVEZO
VKOP+O+5HnoZBY1gud7hmvvKb9vE1FOwwJToDvVYFC2FI66LZnOORJszhnZG
6nuWXPJN+w5rJ1BCZCjeIG+I9haDreUCPrPSFx9LNgBA2myhIQbPcNDOPI6H
/8QxZkfqBTqLn+79ckby+7NRcDV9I+Sfy5qUQFRZ1ilC3iXXrw4x9Hltc7ag
PMxG1rynq3udWx9NBaZ9o1OEjP0Bn5iqlLdXBOsGqFITjDqowM8qOvC80Ljh
1Ptc5EbCClnppC4tg7wXd/RNRStEacBXL1Ll7C1xlggZHtlB9aJ1ipAPXaSU
UedbP1d66CwiBUBobv3sW3os7RH/KLydm02azXSSlPNpq3iRlKeHvYIOrfKH
4veXOC2c/mnBDAuQp3gGvGzBf5u91o8CbVmvppvgYHAZ3xS68iBmh+x9aK7J
V1s7LReFtjpFEixLZJxhk1zy+H/NaGFR6Z3Xnd+dXAWYTfM7yXenCAzmjeL2
3DVx2ExDjzCTLVhaCYVKBCfAbvPEqumW52clwAc+73SKDlUpwTvYvNgSvNf+
H9yOTpONCOTnKBQDpblzrUpPL9ZNMK4KgSQLdQIb8/KNmPH8OoZED+tUKeTv
tKFzpX3odKQS+xcQ6n3IrBFivVVhV1A2lRgtvj71yPNaXR4xXBxUrC0PqqqB
PeamaaKnBmLYPiVyyysjoxnCVAUE5Z/EP9yNF8V7Pt6NNhXb2/AY/V+MrqLb
h8U4MqVV6/w9DHiUFvP7e+Uq7LQltakw0S8VHJseD1D1SEqG/lZp0drcBtkL
SdIrTjUI4D7AbXu2n7OE5ENYQoaT2HIx5YA+ZgC8yWKnIJCRSrmpM9wU0QQ7
/XEH4MgAdZcpjVuwgXA76tUMgvs3kjN6Ax/aH8q/V74FQGQQ+/AfIALM8Gyb
8COHKF7WlAeCro/AUcXlZEdoocOD+nKd8miYXzMj2PDqdEcmB+2A4dw+eByX
XsCpcr4l1u+VSphyOPZrb6/Op/yyKo/kSuX1FsPj4sqF+lfkRQa3frBBOt6+
cKTIsuJ7+ZeazuzQYvCLHG/C2HXgeytlYTKgpc341NvisV9ZgiJl//dDPQXM
7fkEza13C2YfGYN1yLZZ433h1ogCclSamvMtXTGpkh1h19NlrCW3y/ckkIv8
dPMq72+0XegW7g16woW1gvpdv2pB0SIV+/4UfsV/EPe1CRR1gLa52s/MK20B
tT8fIYOY9njDznFAfScphKhQ4cyuU1WHFgFBIERCZHecrz7WRMW5tM/6Km0T
BFT7Y6cfUcP0nKJDw8k8I6kHcwC5GZ8IfziX5i0T9rOYX4o9sFPOtVp/Yh1w
8CJxeRSqhqgGl+IKp9PbX2wWuP35tUzXl3V+wa3LLcZ2af/GhUoxK3aoqt4O
NrH1CWZLuyr7oDyITWasm8Eh+xinMuzHkyIPjW0pZp134lFuVyZz46Ngvn3Q
RQgAOghckH5vM3Ggs4K9VU7u8FqIWb6qwc6v8qFnnid0d+nyGv75cgmAGEhF
A1wHzPKJfcBd4ze7r3Vcw/IPtxIvASLVf3pyEUZpfYvsCuiwRNVVegdXr1DT
hX65jCXFL9JqnoBYaA7bvjNUarH8XVO34Sp7HZ6v1sOuCAGzsFRGeydSKrqV
dm6WZMcOUD7Edh+G91g/47szDysVfiZuINposfriivipA4rXapnJ+3wk3dSd
3IAOqF3QzJaSwKDEyUN1++AlXkVK9De7yY4bOOf0xezuUhPjJ6fi+hl0rxTG
4KnBYCPuhdHDgoLUl0v6YA3o2WbcYndj7TXQ0f/McTbhW9EHD08lwWMsR68Y
7rIvM1Me27RVpx6E3m+nXFAzOdr2P7vN6LpwLWd4yn8gk8sIR848G7hBrJah
B2Qde6iOH/MzZfQvPuwkBn25llyqRUknkAEXpW+ZrBgfUTTwgQouVnPpieWS
7WNeDR7u5lyWMuBmns+/yU5SSNbGtE0m/NZw3exrKfwGPCeXqehB4crnXPMG
J0xI83X1Um5d0hlPVpuY7VOV4zckghLZxC8w0iujX2fEvXmQY0BXs7En+Kgy
+nWaP29QCLCT2yKbJMSqtseze+R3cG+t278bSEkBBe8jzagjrwuHyWqVkGYm
ZZqrVE++kVRAdZ06ffW0AdUxJXEuZzP/Y2T5hLz7YLo/5MfQ16fcZ7XkVlrr
NDJk4o1HHH8eWUQdCc3EDTHErwXWB54th51469pwYF8B9W3SuKig7AUKdHvZ
r3Ju30CJp4RaEbF770Dg5L2Spw2BrZEdQ8lW20Qr8B6x9lSIv9LXI8NgA8dE
uck3VuTNdZ3IyRO6aEQgPPuRSbxkM80OhAn7zUe7fUH3LM9sxamQ3t47C480
ynGGSMn0l1uPT7MJp7pu1S4EbNQIreoX9nL8dT2JQLS8fFi4vNWWYXpbSRIY
sTnNVmoGaEUE6sR/6l8SJbsmyaoKMl4gKSlyHOUJHy1tT+NHkOMSXlDbyiBC
AOeVGSNxW4s6dqbGFr8wvtXrHJ2aho4j2/m+jZEsfb/TAqYPuS0FoO3JmxV6
PTI5vDasTcBK1qF+twNFPICtDS7KBKaRe5FRtGfT4HF6B5eVVIDy0inRRL5C
GcKRRzXYiAsnoPEv/CpFtSwOg7a0jxqTpSJVNas1DM7qJNRCUU89DLDJF3bK
hKSgAXYqspFIQK+TNsZqX0YfL3qB6RIbcoemUOM0TKMdTMO8iwjdiLKMzbbF
9UCsnqVwMnbEqfuPHbd+RwbTm1p4PKIGE1oRzhQNm7AALPww7kcVELAPwTVG
q8LIxHmrCN0xtqFnJU34drA2rQVwnRlyrd0xxLxM9llPxev35+hWjj4cHT88
ybYgQ71b+epkXZ7spp4ItM4ryG6mbVGtciiPIzK4MWb1nckSIerMLD2Uu5Hn
5kgcyL01YfiomOr6SVV9Oh/ZZjLx6dGI+msTnMhI+srwwAUvSjIZj5s8QvQF
jaykv2NZgJvVIzV6w8c0H/tzlD+OKASKsyM3lAS9MjcA/hPz0tNCtlSCiOAC
BDZj/jS+LUaAZeUvWngsYhStbACt3zNxDciM4yaLbBF69rbZwu2o6iOn1oT2
tkMXLdfLoa4eVLgmLsqkOfLLSy6+mELfFFVWna3tEe1OdcOD6w6DRw4ugzKx
A6ts5RRXxGx4XpJd7QD0t4Os7WPfV23LEOZrSHnQoG7wriDtQ/2+GlPMHvJZ
n29GW/oeSPuWI8zHOa9n72LLnM9XnYRhMz84St/VwFWK7vNfGwSTHZowr3P3
F9gbR1P2n2mPKGqFkplXQOMhzpxMqD2XKve98eInlLFY72n//RWsEFmUBS1s
x7XOmCPUjmLt3j1wHsxD6YHp+9EP3YrqJ1KD6UKFNiUMYj6VQMkPpvEgHcmZ
Hmb5dPwiqBVUIigz6+lY8FDACrwjUwIhpTXW620a4c6ww/dfc0SIV55a5Yy9
PlvDjQI7asem1PVqU2FfzgJqr1Hkrw1Q1eWc22l/zhvdWPhJCFNlg4oFAAHq
SJAhtl5UF/t5pI0UFS/Rg/d4+gJzR7A09M4xRYPklxUeK1W2gdkRpvtwAHgb
DIcUrj/ap+tbNV6j7w2o/Dg5wVayeTkXcS5EMBgPI5EPLh7QQA8oGnneoi8I
IX/sEc0hgzAp3LNRSz/O+t0VqTt9z1aiZSr5Mcf9noZr+xdfm0FM0gsWclOD
roNCxM2ygDyOTYginRxGGVvy79pbSjk1sbviDr2UaLjomuPpV6k360a+y+sD
QK9h/CDIm1VgsOR8CSFOJeXMql84dLt+75wc5kToKR/ZoNb6/K9N0cseJacy
Tb2WKGq7rn0drNWJZutbGwNeSRMy5xq/3tQsRcN+/FdQfFA/3QZtkCBo0lPV
Fll/HMLugyg30Xogxp+5YQP1aXpPYKARpdt12J0c6g4gRTY4utUauBcRDNxR
/2ykqM13rdwqQrUbBOGPdEMqTxWYuRZz0oRGs6RXwFEcvKSKRlyLsb2+wOBp
iV8VzUBvkKO1FZrgr8VnfKh3EJDrfTcOCsNFemei83TcV9TnyCk3XqLqdH00
osTjdoDYDIwobdbWyAcvrDVasU7HBHDgeNBL0kVweetwmjFzuRCWWRnpe5xS
fZ3sCdMU4qvhwGC0Io1uy9VPawpYxuDprtMBVLA4PRPpyw2ksw7ul8NElXkm
uvf5VF5eQ0IWh0k2HRBVN3x/MtqDKipFEUcAs1lW0vNuz9DOdiDQHKy6I9uy
yp+hKyMRYI56tdgSIL4G1FZmYsHzGpIuwz9orU8ht1NUVY/GSWoOkCiGfuE7
JgnNtRki4gPpxZ9/CZls9w+DHhWRDvVoaOVRExYLbt/vGSinKIxTVGAMfE/8
nzgT0dpWJ1kE+/tN1WX76X9ulPVgra7YF3AqyxYEQuna+9pLKB2RI4hW7O/p
dWqqZsUQelylNPqEdV7WDLk4jvRJC3cgf/dxLLtlKlacNKfDTmzi9HE/16Cl
RHYY2rXubZ23wMFUv6NUSFJZ+/3dJeFdEdzbLWtYR/O21Fu/hPpZLoYuiW4r
AwL3oCnFP4Ll3CmCT0rMdxmRNbh0ZygJkLrLStO2YDkpiew+z9F4flyZceV9
ps0L9FGf7/PXxn5Bpy3BblHSLxeVFgwHlrycW7J2I5YjmWrrgIxIA7WRu3Wf
871nrSnPtONaIb1GW7hoaOrxiBXbafdn6a/taUT+uxqiG1zrWKTH5TFn6O/g
/Zhw24Jth6rK1tfAsnnynmKhGpsngHyI+TeMBHmQJckM01FX47H3P9xbhE7c
51BnXLHVvffmaErw6Di2MGbIcJ2P5G6VUgBzfNkXWwhja8F42K8T7VwG3wvQ
dtuLcs+CTRC1p8ip1UiWxHp8MjvLv3h3Ta0ZWjjrqdVbpdhwk5GJ/bOcHN4l
cUQcdOcRYcz486sEG6xK9Z9RwwOjDPTxhFwOPRB56NnTJcBXGJfxk4ZK7E8E
oKIpuq+r3kh++IeTEKZUlf6hDeN2UBDONC7A66mUPtN3gkFhIWvnz3gnJFbd
YLgYB5CCAf4OMbcDxIIoB7Z2Op3h/+zZUO9vTnPVS727ZtCIV2KwDGvPbS8c
UPUqzkfGcsmkzpnhCgOGlzwnpiqYxUOzmx9A0F9ENhj8SMgSwxtSbnx9/Pe5
pxy4O1TER2FsWPrSqnuajG0952ElKHj75oc+Kr/mggJbxTjN+CWi6kqwKxiG
mVbMi9MGurlbEP93oQFssQd1L0GofNgf9m+3SsaCOH1QDWE9EnLI8VD+OZ5J
Qix/k5kw7zaK6jFbWUEJpmNccRSHQ/08h4aoQuo3I7mwW1l1QjUaaAYAn0Ze
JlxRHdV1zUt5Nk9q6KOvbrRmjF9Vt9jLh23+st3ar6NK8ryb4G2Q10abNf4q
IRyXQ/KjT6fyZRucGyiaEioMQKqk+0/iNH4Ec09GiIIrdu+7NHmtp/YK4Lyf
IZ8uVReHhVusVxzu27nCQjI/MGk6nUgSbyLjwP1ucxcLWb8Ep5wvI3LDTzRe
xgwvyAI50eb3bPkBoGEN5n43nuY6fZd6puSVtQXeD60P24fOQM2VGjHFFMmL
qRZYO0gdH5cFDrJwYKeopdxD0bZ0Kmvbqd5X6kfxHMMSo+KoodA95bjJnzrx
Cz+IBrY4GHH2kw7+C4eF3yVYG4aGeCEvtR1y04wUqjsWGcOfJpHlax0fXMlP
Fx98olD0VhLV6SLMzPZGi7I6MGIk2uaMGvQgpItdBo8pCVIyRoKiR8C8R5b6
8llAzGCp0OBLDWN4RfV99wxEauSyogDcxTOEFtIawv6dSC5HOUYLeUzSNlqB
NFZIRkpAS6Za9k9u89+aABhxlcL8exShQJ5643uQjJ2WR6qKLarekcdIEEQg
+Z12ln8U8i6dh9e0Gb7w+t34xdd6EF6zZ/FOdPLCt3qV3bj4p7P0mt/biYgB
Azd1T8FsFn9jyNKVsoS/uw7ICwZpkynPlW/i2RklUKZG9x1u8B1STwrUBqs5
iqf8Kp4Setqrsc/h40tBUTqi49CAgwusXvXcYL/AIdlSYibMMg70MtUOsaz0
akn3mMaVjEpQlkkabs6zwYCFALoIhoSNV30Mraz99hDc8KGSghmgjBVFKdfc
4a1hikzdQv6C3TnqO0sfur7WODMSWAbREWNaucQJyu4/Zd5AC6YPLcMmYyM7
QF9IZGEyNDHft81jO0y3N+p6KwngDy1PeXWqvUxedjyvt8EPbprRZHLTHew+
WKYH9PkpigX09IIRU1jz+MfUl2//mQhTTVdycq6MO6deVad4WGOrJXY0ohfP
uFwQHB3XtbBhLg8NgjXpy8MAYnvJSvwrjQkQD+z8GiD1gxAOtVl41JV+lD77
PykSdb0srxiHCCRYQ8Dn5SqflO8WEgCm1knHqXRJgUKBsByZCLOdojnc5LFp
uPm56XZ2SwfGdLvSpVkAYKwUzByjaXKUXjzvbuYsNXKBoYV6qyWU+r79TXPq
b63Niw0tVMoF6QaAf8SEVWg5+IXkQkoF+8YuRXNdQcqjwVpk59vk8P63pQMB
0s3QzJAaeG+F5OCBJl+wTXbT9vVKjVNX4Wktv6xTyUYkITPPBJCpzmleRyZf
k26HpJJ44UqZbXVWI0GLYuVT+2anOztVqDTsWn/BurnpkM9E6noZf8b1kUzy
2C3zO2LP8kjGGxZ4GldyNaIgPv23sfhV9PoMT0xLSy1JjApeP1OSSwmK7kdM
SgsfnFJxteEg2cqoeFBCjf4ig1sopOJnaTpLeYimqOmZBcFHnSfRJJbPcrGV
k5gA2w0dqDAlC28eR0+22pqPPRXK+BhkUVkBhAp6kxcwzS4MxdXMXGiVdo3n
kGLmp981keASOAeJgWcnsVafaNgFcYauYF1LMkD5Dh9aPYTfdE/wmvs5+ylE
FqDxN2fu0KntlmQDhOWWNPvmTDMZOkxysSdbntU2l2QV8JGMIweeht+3e1x2
ajlg2Ys9xA+/jGkR3LJ+x6Z2anw/aGdjF75HEHa1b/+TL0ApbnkkNS5A2eK6
XKSCJcJ+KeFWXdiSk0FU6pM6pcOq3z1Ft+D8UNHX4cA6vqPLSgiKXQJwCiA7
A5wVuZt7E8rW7BCpGU1QxAqWvKTEhr99kAz2WV9b8w2DSUqo38izg1CjyQ94
s6YPsNheUQ+ynlTWDVdSiO9LkV009KfVHEkCnHowjg/DfG9U3E4+/W5yBldf
J3UFzXPFHZr9P9qHLfblqLn//K/T8NON7zvsRXEYVIJkTlX9pGNGRevzsz/q
dzWKi7VQq7KvvedBjo1MrEB+TnlbpXrdWQFG/mm0tMg4UCHabF+p5EGEudVi
xYIC9hdf/b8VJ0mNPHMPD7gwUOj4JhI0CDul20GfYoEaBiZMbgGdp/fGyX79
GbFgyOF0ezyx1uKtR2qVQnWLHXcz0kfcwgHDYLnriVwcaA7aB+4UWj0ty4it
I5MzDoOYZqRGDKUjkeHtA8Cr9B+zIi6PG5gjPgR8YanW99erKfwOewCUUfEj
JJKcyBF/fpMt1N3nORyi5ub8dgHPPNmajNYAT5ldzPZXCHB2HXPW/o8CXet1
82DEFa+1SZkhh4JIh3xHXD72aMtTsORjoGBXWYuyfHkWIHEje/EWHaZbAqTm
kw4yaCU++7TFdAdLLLGhmv37YUmMQP3kC9MsCaSEz4Ezz/rlellP8eVmh+dg
ErT7Qovk64gU0xUrOjTCTYlPk0ytpDjtSDSB63oQtvDZ6VijWpvgLIxQ/b09
cS+cvvEDqc76+3AVNJFoCOfJT0ZiafEqzoiuOjnJWuSA19Q4Thv9eNQgVlvd
2FaFhoAjKNbd9GkNwWoXHa6UFdMOCT/hSQ8Jxwvydl/cTjWrQCyQ7zyuBgrL
wUDJMAF88bCYlyoghn7+V4R80qJ3Od8K0pL45D97MEdpF9z1R7eno/QKqojU
7CmhgmF3exvAW2BEJ+ztEFW47lSmtMjZDC97b3dMiED7hb7BXn++ldw65Tlz
gKnZwEMSDo66ds2SX0zdA09OWti/0yeILrU0qfP3V39xwCVsbSKvprNEwgcN
jUqjzE+mfqdFr25Sh0+riaK0EHD5IPauATWfmnTPgpegHo+BxoHnmGL4U/Qf
fXtm406/1PtY+2HRLYIHm99PYyykJ7o7TfkOuZhOtpixjK312Z6fZe8hc1wy
5AGiq71rAuNR+1lLg62lBdYXAP1i3JHJTaZHWF4frEH/tNkFNEqV0ScTlzSW
W3Xdkbhhhv4c8WShY4SIcnfyZ+JJ7ZVjTJIV/bQNff5zenyizskgM/jvBl0I
Hv9Fcd80uZ/cPzKagmBEllNZqZhzgcuYJvNV2nvI+eArtblb0oQotgFpEAK2
rgh4oF2PKyXqWXz5tbp/hcMLiRHRKBLL+AOOWj32223YP5KwWNqjs0Zy5NrR
FU1Hse9JE0CzaZSlXnbeRt5cyQt7zK8lW1RnARhg7aTDLTqqUN/DJgVPHnGo
zuPfvuZN0k93u/w3x37dqnRCp/0FajHzB2sHXWLXdP3rWCm8MB5P0QQMUfa6
Gml1sFRZGCDm/h/DPRpvloDz+IWw23M5dzokacZDGUq+oD3Ud7qFrx4cQzdx
Qv4WKdr5x8dx38ofaPJqroZ+E/45jVJVWf92A/pRT1Y3tZFPXucuPR0JH2jU
R+bDQ3a7VN3tSHspAVJl09qodmufI414hcuBK1B6fnbN9+7/FPto0vCRBg/n
0jVXiW3XqVDLpZFCLtYxuxqS8POnajQe5pfTTI1fIzz+ToqB3CloWUezuBI6
Y1Ct3n8O57ZRVoi5CRMSElij/+9CK/H3arok5MWj42zlytlNDfbfUU7AI61/
LPcucKVxmWO4EREgV3DGEV48dpl1qIAvkSOX9qh4u59xUQwZwqefMjhIIGh7
6LfQfVjJ5M0qxnGauDg9Rozu7GL6OTgaom/YiN1+UFjsHWo8csa2XDXmkl6Y
fapxiQ2iVuF/gqqwn2LzbCs5AlGOwr9IIZjyWhEpiZO8Njr7TwQJsbwcaiVs
E9DFxtWwC/caYIrJE7yAh1kzcQcTZTp3NC7fBokhlnrFMKKcmkkZfnI5zq2s
6G1TwhDdKtq7ti/wjdsHbmiewwGmZW+5uB+5bLt8JbTauA68BpVoR48N1uv3
AIZgViz+82jO0DFE5liYfshX6ua68kF1PtQoPukfHFWpiU1hi4tNentm636I
jdNEGo3euw0QH80+hg8IE7YeHUvRHAwB1Sq04X+86UPsO36uT6QhY5BHgYG1
erM4jN0y5nkuCu0EURSCv4AKj3+KiJ2OH5g0pI37yPFi8/w+baCgp51hT/Ze
QJJWkFXiztv06lU6ePICsYjFVTCc+bs0Z6Ok3BsbzOJuP2HHivpph3SC5k+K
B1YGCkCQssrcgpBo5s4WPCwbQh340LEt2xSx2oZWpnNkSsgqTG94uelsYshL
qeA3YlKpSHkIGG0mm2wgdlotzQ4eOoX5ipIpQuk+LXjz+zogy148w3SmW4cz
YjjqIqpileaO7vzzMMJmauibj9CJQR2Zu0n9RogjmyfT0pY9TUCfIL3lMU+K
i4aFohN3ROTVaxeXzY/JuuZaajI4jTZEcEgnsvGBJ/b4jWCSd1PSf8rfUhei
LJ9HXaIMduVL8wsScCU16kqLZR0ZqgLonqmHUcIrCWX9eXKxJBm4NIqPjlv1
4mc+l/EqrhApA+PUwY3EwZFF94J97uWxC+MOU/1oUxBu8kOA5qFeZTDlKWsj
tHiYLX6VPBrDnA0ZZLQo6JO4YGz5GO/DJLBKv7bGeICDVCdZlc7A+SJF3yRY
GUFJgj/fVS4G1UfMcX8IARqLQbhLjepcXLKPcJht+EYhOPQ69jydHlOqT084
30EETjOktmLZgHOJh+S7NwOm1zJxElW1Izgj8HuJ1e4IsyxaCIm42emZAwzM
x4haEwOBOEceo5P2Hk552+4blyFCwls/LsfouUC3X4kg0cOw6w0x4ALl984t
Z1/qvCu9dvRCk+hJa0rXBnqIE2LJ5I6FxblXoGcKijcOhVqrtZKHQWjJ4957
imUkevCF3qWDPgLLSn+7APZLU2YrOS7wfLlCaOfoGdkGI25w4+owiPNASGVP
5Yf9chh8DNzsbEoFbiMNz7rkuLTFbcvoUhQXd/EYsjdDxwOY1i8j0Loleqkv
qbmMYfGSxnexarRKcnlsEwu+6M/PkA/ecilSuok8UY9drAIWEKAgAs8Y/Frk
R0TJG/NY4rprBArXqLslwPiqQUrKZ+HzNqrDNF1palatkLKkqBvI8Ocamxa5
kHoA4pAlnJAXjqjjMzh3/xN4ZCWLgleplakBJR4me4yQ1POkR30xQ+RO9g2Y
y+Gsf1Yu9O1Y1WHNmEueUwR2yQ231qrt1n1//ivT41EC9rifKNx7COFGgdxq
pI4NO5uJo5cNQ0fbHyOtmahZjWhWkL0LLzPGjQTzWueE6FHdmZsSBQ4iVm5u
zt50sNIPctcHTh7UF8/yOHcPXjkJKDacA9v6whyf8EZSfZk/S5WGT1ZT5Mac
C+t9oxqO/vUvVkdCCy41/zdDxi+4W8FVNW5uSGWtJmWt7uMvlaD/pYzqh30E
Z4LgLZ8qnmUbEi8mbpWDNX4a10Hs4CX5v8AuxEEO0KIpnL3Y5ELcZO9qx5RK
AAtp65LcUUSM0skLu28OG7DBPUtrCxcD2YqS7huDDwLYUwZjXU2l+19fcS6t
pRfGQYR1ebD0Gcr99nwn/V2At7P5dXUSlcYQLJdpp5fzIhxOx0QtNW8Uuxoo
G7k/P74zYaNj4bFp9ME5tMnKh6Svpuccw+BoZVvd2LO6Ofx8mItUSfRCA/EG
jOwDdJq+hICYE5xEG+LQe2OyxFcmxZ9XcI0AoXyFY5LHGEF8MJtk2JCjpJy9
3L2obelaZde8/qYfY9pdoFLvoaxUb1RYiZ3V/2TG5IbpYjoq9UFfJiQMoKxG
+TXCkgRleaDlZ6BsUU+MVLJZ8vFHIfrpUS0bK5beKPLYrUDAXPSgub6I9Fv1
HkoczARnNF5m3qLtEdO25aMfTxoIUgzi9vDv9KHTrB9PbxFEnFdOOWyv4C35
IGVgDRNG0KbpHj5NMIiWcHFFM7hBDbrWb46NNH/kHZeeqNHh1ba9q4eLe9Sa
t/fhrXMXYhgy+Emph+jVpr+PPgSG0Ev772jf5cNJklhoOWEf5EovSIbqLXmQ
vdAA/wFbDGYhKvG9GvHbUHTAa+wCKaxcHb9cTLVcsIrCV16k9vPKYUptDgAP
ptKAJCKNSsAfBWOzgV/RNn+vzqhrM0WY/86TlJTmZER4cxiRjzLvPAwhB9CR
QoseCfqBf5s4yuSnTifLu2r0UrzkHvYIC/niOtP0CsTQCbCKVnNwm8L6ZGxz
5KBGZTFhq/HsulY3D4MiW9lHFhO9LEh6mv+h3IWUxRnoFUSoNE2QcgK+yE+6
BnBxj7LzAhL4x9105JO/ae1LnhjRAOiOTIFskBD95lbHr4lzi5fRomoltntT
0HvwmYuGj16GArf0RMbqiU6UOuf1SwWqZEqpFTVOT3BbDV/rpIHKXTiJUmkx
niu85sNMWM+CQMUObRi8zxZEj9MQuhlnp8uacd71493WrQ/Z1NDoTqYm0NKR
jqRLE5CiTab60o6V4SvF6VVIWw62RdCMMDXlDfpFbVw4tXzE5k+3e3+kCDWp
FoT1llwGXn/lKz5K6NiJAzWAOVWR1Sbgz+EG26I0oucUH6efxTzJK9CEj1i0
hbP0FNm3Y+kbQ7YhlXuEg6Y+CxugxOw4pT99hI+jd3g6+DpsQ3zlCrEQdK1a
DNatIyEcFX1bCV8J731g4IYBkVX71qBGD+ZS2Si1U62tHk2aijmvGd0S/BJb
CCMxQmeJldGavXgxqQGCYOCvOLrg0KYPgVETe5DnWF+8gcXwBNgdHpOzmnOl
1VMtNlizcuBpW16Fru6a05564L/YMTIK/9ILZ1o6kkdag9N2R8zczEL4qebc
YJoeQkbgQxKz+8KXT+1ddMvUzdxSVibyfh+5+Kkd1+T2EhAsKYvVx9Qx3EeQ
t6tV4kbB8HV6GqWJc+ABokb3ImEwYzGXz+8zJGllNLrS1cnpPPdrS8wCpmw8
BeNJrtqb+AUESZB2V5HZKv2tDK73ypB/wWNJW7a2MKtlrO+dmo6lL+L8P90H
Pox2JPhwMdyQIWIOjkp+6oEddDIfVbx+kNpoCTQTe5wR14G2efe5pfr4+0qd
ZA2nj/6uoK7cr3uESGY7anyzrowWgjXMkqTgwxzb4plE+Zs24zoBy11wLMQj
Kyq9XbKKJTyOxXi/0ZVWyuu67IcosZl07rL6ZVBpjMifLh2gkh453a8IKGxE
rDfqumUwSPvuR4iCjMcZN1ksb7E+0DoiEDobQvukMYY7S/7Q/4MLoTdQoKKJ
+HSG53nH+ztwkoHI2sbPu4NudXjDw6lWJsIlUN9trRXjFotbKaNnQAY7mR68
7phF/sM8LD0zlVGo3LChMz26ZsUhUdY21DpwouTDLyRNwkexZSkMhmK6p3y/
1fopNewsj0qOCR1l8jowE12yH147W48nTmtiOmQ9D5cnhLdx98ZnrgvUMtru
rdcaZBC2KM102m2U/B5Xw0sVI6005T0hjGd3ArcE8lqkOh25AHIECcay8Ugj
7b8axmZg5R+JRhVPaHQuGg+Iz9PwBxex+TsSYX4cbzHjJJbivldO+5hoXIm1
9dbL9PEyVkdzDhS3AqLfFg4+OhRQgnmgD8QZ5JYiD1XzuXG2ztfDMT0Tpe+2
EmlxF5VgGETPje+9q/LisCBqN8ICQKBivIU6VZKWShXlFnm/VN/j9w7cdw/n
cEqVT8HL7oYH0g0EzopzOWL3i2BDyvRm11XuBslChSGt+YPMV/xUhXjssvN0
FehnNB0d2Mezne1RzfTWS9oRMnVvX2mqNRlXz/Zr6Nuv9q5ZjNxlgodmFy5B
NJlbnODIa0iOS2eQHo1R45fgi/Ef/oExZYVVpVtQCC8HkUbNKMiBcVnC4C1v
l+RIUXbnYADFdyByeRFTUDOFv8Y2PknkUn39fcG3cxETp5xbdoY2n68JpyB3
cxWsW/a15heTKcHriqpQ5sndr2tRSS9eTsPoN1uPP7mzAtt03RGsENJf8qo6
iwC/qeImZhAXYdc2uT/UVTBkdO8TEb22IMnb9LZ+dHOz8r0eyruiTdtxWY26
5pSqCu6vPI1r2vqfchWdIQ3VrW3GAMMZwmOC/XORuXLfw5jk4EV2s6Fsf7Q/
n89clCiYQqKCLPS/7vViXLIpKgpCM4Lq6Oldkd3OirFw64UYlo31RrJNxPf8
Jxxh8Ujy4w7fx8SEDJPElE2jIoaUc5Ml7msXvL0LAsG7yFkwyyasQzEGYY85
gG4nLKQtBeUyENkP8AreW5sWn/p5C7i5b9+BkiJZu2oF4xgXFSh9XYin558W
EXSdaCTOa9bwEh8kH/85AwwvU4JUPQqU70x6u3srewutV7p4nl4Z7FEDAkfQ
2GP7yaQQc8EkWjzJFXnIJgT4aqPgoOfh9ThVR84CBZMHXZf/VoyQvFPbUq2h
1AwXzCQRiG/jmN9h+j9xhIBYPxbThAt39vzNRt99+1n9a5X6eJ9hhyAgio9Y
NRSFctTbhf1OO4tTu59sTehnQCiA89dA1OSDHo4I0Yo4pvl9COIexGmgsL5k
EqWoE9SuKrDiX/+IrKA22HBfVxGJ9p/oy68UHCSwTpgbQFeTbrScHS4aK/9H
6SITGXzLbu4tJyzbL3qpGIIbRbOZCER5SquVuF8MAFloHPma5gpmZY19tGWx
4k3Wag2T04KcbcXoFCerK0lEPnb6XSdgpRzNavxWqFoSFYBAj6tg7h74xEH3
Vl9l+N+AR4gD7O64muEWDYi5f2zcfWjPMWxc0NtoRfrOXX/88ogBPBix/dWD
pJb75cEcvfLc+mXT2OaABOg28t25knjEEAbbni6O1gDzKNTjcuxCsamVyPUf
zsG6bMzlO9/01gIJpiQOJTVn6iceOIbDnrlzrlHFTyHQYu0HQ/Ft2H1nb7qk
xKU3ymuPxveBv8IIbXLa6HW8k8wCB8hPxSCIEBoa8yNmW2MHxoMm28j7TQp8
WQuu9DmiP8Qb7lJ4CoRTN8SEAc/Wf2sc1Fs5fgK41/QO0AF6byIC5UmZFo08
84+VOsOEZkR7Uo5qFcWC4GoKQlBecFVtVWEI1FU39jGJmuqScoYe0OkuRBi2
cXvtb3EQ4sUQhwLZ7i5W9qby7aJNkFK/2SECvpn9VLmisu7PQOvcmRlkHZAZ
5kiRgYMV0XVTWfhjORPleZyfQT60G7YLcD85rnCIsysp/DbmVpQdDoRPP/5E
h+pDMcOw2mkmc/yyU4JyNyHQCEG4EAgM07TvHemqpglpeYSUoQxZ08KAJTJN
ABMZCn9XZNv2b1W/Hleh38O+A000CtaIy/J/eEE8OHzRYBmdN2NWt1COgaq7
mgRwzALBcm9H/X0hkH5oX0dDKFDOdfapSULqd3wV+b0Dn3ePxD1rxnxRwmg0
OzYeSc418ozt75SfmWkP+3fI44V85Yde05kwETbVvRx1iCxe7gubWVgib4oK
PKIU+S/emtQqn7+paN1zr0ClQeI4aTp3FNw4QUSo+FTOaf0Bjl4clmAM0FUV
sExzN3gT8/1Aw8nLeHurGp1KkE468hPEHc/dmageoa98IHr1NZ3XXogl+ppm
CYw+2Hp9jvh0g/x4LvT2t6iEzhbRp1iq/U42LWTdWiDwYsK/pmB1ldLzOMbz
FgfJzxzlBZBWDcyKMbaMAtJlom0Mr84F/NTn6gp1I+aLPd112wXCt2cA3qb5
OKEtBKS61CcpVjyuyE4nuh7lSwU8FjKjdUwl2XfrVvE1+qqb8AZDkAWDNNXV
n+q1GhRqTgjMkXFcAfoeObv/hWO19TYyPYDonbB62ZXkniBrk72Sa38iCzi2
Qso8NGayibHKUcSQph29xJZAHLTyLppgJ7qsniIqeXJp2iDvDzlUgvTBw9/T
lHTIO6Ed+Wa3o2b+/2PFYkNqwvwchWd1qkR3YTh7vF6lse31IJ4XrM9BZAqd
Yuds6ch0JH6iNswqqcWKaT8OR3Iz4aMlxKS/zFgAivIFUUhUA8lBXkgf4i8X
kK52xpCMpfoSEpF3BjWKUDgQ4sDYL4OBL336IN9c+vPNV0F00mu6BCu0KzcA
0RuPCck+o8g3V6VeYhX/c2+2mazzqe/RdjjFB8TXj8Xc932InbsUmAPl5Ogn
03Arn+Kzb3FfVsMHMIX9G1eGl+jla4uMtubDZo9KhcUeRLvmdJDb/hCdJTAI
Q6dFvEbJZJdMiaTgefZbua30jnOAMpfWEZcwmRpFhggxIueW/pod1jV84YyX
Kd80MfhedbTI6pnjdjUGRD/TT7tQUb1Tf27NJTrCOfp37719bny/aAfRQuNz
KMn29UBqOkEWZ1t/skH1uhtLS48MtFfyjvURKcCl6DDizfIpyJQwjrnvrnBl
BJljeYwNvOWdqeL4G19ZQSrzHI6WsLfm/36zw9/22Ht8jrc4GYbXAsDFkKVS
lt35NebMNgWkNFG8ddX+JWV/dxThX3CKAsYDlNKrEXmzRc+9UjExqznONCJg
/PI3jiB1pocbBGDy2/3FH73Mexm6oem2NIYAQQvNUqet8vLIfGBn8U7fL3qy
jUV5/oRf0bNF4aTMHqLEfcBmgwpFuv7D35zFnlBRAOYJucbmNBfq5/PG0hna
dXPCPAs8XyWuJ1cY/UxqhXUKUx9ikUu674OqOq1kyz6iqkPh/2GiYEOzF+6U
fxg50VdEPq87TUOOqMJtcTaL+cAZFEgQUMvMtvUAjehkStsRhyuJ3MAMDO4T
gP/PLbLbFf03yMwjIsQ5cBFMreOCGFFMmHWCbeUz8a/ucrFQbWWhq+jfhZCn
seodSzjHghWP253+6PZ7RMj4Dq4oVKcgcpwgo5hfn0Cz5BNphcQb8xMCHSCg
2i+f/IpC4ILgcmmL+wRPe76TYWVaOWUsNS0Zy5j4LsebFEovG79A2KPLy5Zh
CwnbNlEV9lyeBjpugRNF50YCzdCwqG5HA4ITouEqd680BjbKVNpJewZq5ph+
8TsrMM5ALOMVaeFi8TMTbQaWNqHpiRAU2kOc+ko6PucypjuzBtUnsoz8H/4E
fpOskgDFzaSI1Glx6bga6HP8vT8gbAkCmNhjwvUmMDO7EcFzJft3j8i8ahEt
giOdwLcdwAyehPcgNA/jD7H/8tMUOf/kSOsM4pKFTLl4b1xP3mtXBs2AYzb3
vLhi53YhSBbNpuxgljPr3qrzvU2xTrWdD/F68WNsWL1y2gNIChOwcjSlTONF
dK/cSVP7NlFgXN2dxzwEqt+Y0Dy3gOtwP3UEpKS81P7qLie8MOYXa8khtajz
vvp2epnDthIy5tsNAKMV7DDjPAUw6Eq+WxjlwFNva6h+ODJqVSjm+9geUWOK
IcMD9xRRNu0hpxenzoMEqENczEnA0HpGQp7tzwCaLqmlCs4Qa9ES3H1CaBfs
KiVdWRy/6Cck25+bNGKBdYf+xDQ+UK1wBgQyMZ79gTDOPndcYbfyTOQa8naF
rB31trsqtWIFAKjoYvoHQ3fxQZjfgilEP6IrnZrvn+DNeBKTSzdykNLdak5I
jcO/7iingXI7UvF6+plsWRNTG2YX8AcAia98ChoG5wq9bVgteRauLaS2JWAs
a5HtMrlg3doCGE6BbrMLAGwNcezDqpDd8lQJwijRj5PCHX0cRKTEkmoqxRg9
/BmnQHxB94K//BZvFHHi9oZ5yl8s2zKRb4bBt6/MVbDfdUx9cARIaAWDpvlm
KgY+Gb/pRGdMNYRPB9Ui80M5lGQbX9x6rXkbbNfdXkdP9vFSqrKink2HWnux
bet7TJ1k0qkDw7UK4DMgxB0NG6w5tqlZSfGLVN2kVa8WZPJz2vuQIsLowpA6
7jJkFAz7dEe/oARL4WSVxxH9QuwujbF/maQIhVA+zl2o96AL5jpO/7CQzHN9
YEI49hftYaiRQWBoh5GAXZJW9NvFuXlbMUrXd9nazFaUtwOGFvj9EaY3Me19
LiG2o/KpFWfmngmzlsPXhwmG1sCBu8INcm2KDKlwNHY8OkU9JoHq3Cgi2+7k
8eQ+n+SGyNLl3hJSt255UynGtsrUlf/GKlyFTpXoRILVhK1I6Zf4eTQrFNSA
KUbnsBshPCw4pA3tP+Rp61qMWX1en0wZHD2JQnxkI3pa35Hd0iTvBWGQrv4E
aMG/3BxIVSr5SYyYhzvC+/SmdhN2ebZ0cUi6bYwfy0D4aMnaQaxcPxGZRKd+
sq9mqYV9mz/vfoKFUBA9sH/CzFFHmhhK6gvipSPqCOfsBfGpEaoOPyhWzDOy
QruHDMGZy4/d9HkFOQ4O5hp5GiyflqOzRs6lS+eIwrBYxzmiKzt/ZDKQnU1O
cS9sVgFixHtazhKBHZnNkwjSTQZfosULqAtBwPO8Jboa7hXZINj/8zK/3Zhk
XxyzNpDEVCfrfoAaxAJUpCwRQ9nVTIbCai/zmYkMp5XX6vW9pbFtVx/QekdY
Pqg9Zx526eoiLKxt+qj3nAOSROViLk7d4o041PzDjStSNma7bg10Ywuc7J5q
Fs3BAdVFYpxJm9Qr2E/CO8dcGN6+5sqbl1fXhCp7NeE8jrPFdwJ/tEZqpzQZ
QMuVDknG1HdCertGTv5YfPN6QRFShMqtwk2TfwrQ37eU9JQ40H69qmuZ9/xm
gOBWMA95dJUCeKJscmi5fen793mnKJ0Sv8n9AmxqzMle1EYBWRBL6+lfMV92
WEZuZETHKBxYqDjyI2clGZceUdBrWNnKjnojlGhkfpKQgZsSxbsfpKlm0pj4
s1KdF/ihzBL2MA2pXFFtMFLUvq8BeP0reVgLwNTX7IO3mbh3g6FTjmcJ1pai
RMZcr5AMpjykKeEiZTZQnzR++UNDoR5xVvVrqMW078jhR+d0f8n+bdcV3fcr
NNEhsmhFSpeDpqwl3BMlEQwDJpeW8TdcTAEFeT5c94XqOSgQfNEiXiIch/Km
uQ+kbfB8tUnjM0jfoD4n1RW+EsfbcLkgMgVFl4osksWTuqXSsq0/dPYE89so
WyAKPpAP4dS2hKhutVg8qGjb2d7EzLEg08aKF8WvTL4V30zgz+oKAdGADkxh
VSqYFyzILlZwBfT4n++JNON+KttZCkxFym0pgiYQUPLTnocluj5oYAiykVdd
ke2oTjUnoKQP4KHJA5ubRYbRd8F20YQ3JHdQqjDCV3wrh6e5SpCP58RGoR+Q
GQEgXLmvguaY3WDtV7lSj0WxkuVKu28KiQIKOsdZjpOfzwkTRnTkqtUpgNld
w2tfWJUHR0zNF5gGzoQw7VShhnZmMOkJvR6TOtBR+nJOp8PTNwC3FyW6+wnx
CSNqiuDpmxcV9X64faYciEiiw7xIrf4g3BXxTseruXhYGwWO1NaAJmk5Fs5h
4VFBHMH6mGSYlUQ2isDnR6v0AuGg6XtR36lO0vKrM+Xos24on9ZI/A4KrQSJ
OXQx+PUCvQexjB1gzLlZF63cpvNWENl68j+NAK7H/4mn642sMVpU02jw4cO+
xa2SnrSO86AL2/Y1f5+6MUtk1NHDMBcWbg7ZLGXZSCe+4d0XcK/tBlGa2j88
QRo985vZ7l1aFGG3/m85bVpIiyA+JvWpabQZw3qxwiotcEft3lkckNDjPL/I
PZpwX254aDOsrOd7eDVjvfnr4qfs6jn8ygak+skYYNzakd3pWelzxnXIQog+
U+85BHfhJ2YyzkfwQssL9kaPRjzXNzjynvgyGqzw03KPE1lKEWUHS1RD+FY9
JgHO+rPs953qxQS0Ln2NCALwETfA8X/cE89SlwUy1zOVlUyu0dFJKxhbXWsH
9cOI/RnUmdlu6pMhXUMpKSDTqh9Kg+wbEhjt4yhx17pFqNaCLJdkS/pQ+6pQ
Y7nFQFJjRFZ5mpz1l+isVPhg9ioXffSR+fhH1KkC9DpmuVgnszE+AG43q3At
nzVmq23KOhEMoe0iBKA4J9n+/P3YsUls4aTikRpr2t73F3U/Ga4K3RMmS/yF
yNFxEqUFTnVk9ekoWG+YGQA4MYfpLfybDiqsmgGjsBja4qGrp9xzeyGYt03e
1pGkZVnwaSX03Jl5wuF8UybFR61yR2ErFo9O2gyHwjb+QsMHlGycBEzAn1hY
pvjSCUtg8I68OnnhnenpOXdeGXOY6tNHKGIkDWVH1cfqxcYPw0yR2qSQvi/F
+FCCn5KfsJmXFMbRo0pH9zLH3hWPCt9YLRN6Qw4SGPdZI1MJQ2DrQiYzPrFv
QfICtl3V6mcUdcwMPtpIsZMmgFbnG2kU/Si+A+21pxAYwNrpgj0gZIRyG2bM
Mo+KkSAud4Z9cWpEMAeKM+NAFexBYEPUArsFzsTjTNYenDrgpjJKylwW44T3
ymy/FqU6Rb7CRGHgerDLFz64V9+pzT4a9loXYDakeCR+Fjm+ARY0iMwS3KL+
6Iky/9V7Zakl+fVBtSIrOA5Ik+iwvjEDuVXAsEKx5k+0wdStTrs+/vqNDLC8
K+X/ul0dwM94Q0DiwBxf/d/XF/3gYhufGdY30ah9eK4Qg42/QcIDsbUb447J
PEEvSclL7rE2jiH/xlD10m8e65EodBeSO1kR5V34KpilBG2myFcL1gwjI/2Q
NfRDPg5hFJibJe6rIIg4bJS3t5yDIFCoboNHH9j12bjLNFIXkuQeeTyRMrn9
Clzttu8GnIi1Ax84bMTtpietgxjDxHIeq3vBC+p8Roz9ZY9XidQuc2wIrsiR
Ap8pgPjkXRIKzuX9I31uKekVfd1EK7slAwHiDMEH7kP1SwOmU8o3fyRsy6G4
xk9fFOdYx41TSctirbxakPeecvm908SGkqpdsINv175BqURWW227gK1mG1Xt
Lj71M8tNXrtnPkD++CWdNCPExbKSaq/CwFN0XUFPh0spFhixvwb1eJT+aYL6
TB/0snNUlYPQRFvL7d1QXvYOl/60wMdm+MHghs3BaVoDuDm5WeDwBQIi2IyL
s46GDGktLxVkeivgXLUmqLEjauwCIBdJjYh/qFfBcKkY5zgZQ/cNdGaiiL36
UHrzqxfVpgCXv++JoaksKIuxryP3xkrMUoBODh7NQGqQO3zO9gsY+FGNrBdx
5k3lcy+I2CVug1+MJbgdGm/BqLq3OeyM/hbvgzFYbxzE5gcOkFp8efEBecms
KqQaXksxP9JkKTXRGgm2zZGnBKKEDVPzs0DIvEla7HeB1TF4LJ50RNQgFDWt
AKDF40hboVN7ZPDwXERQJsB+Q4Aq3L3SakpwyJkeTS8QPeyJQrnmofjadzkj
q3BwJHG5h5awZr/Tc0lnNeE7vkhE7n+dPV9g1/qEHsfSjAhlzgDRMeEc0gRL
QgfhbK30ZDtaCQF60i+r4pNto361PNRHY6WSgFVxi+pmIR96UGJfrkywOgCN
PyeJsrqc+QVlYmC/caE1fZvhSYjGgSTmuLFYeI/LNLiJOKUD3EG4HHfjPnK9
iWeKLvTqtjTQ8iPsGFdhBxMeORefJcg0J7wfyxLontwMMpFFo7O+MolE9ffC
TUf1pezb3Es9T84bglwTZiPC2OC7zjMk0KXdQRActJzoWKTJcVaVumfmNiiJ
kd6KunCvS2p0SSeXHgUQf07hUJcDQw6mE2222n4N9c9Jrok20U2Z7hvya3gY
Fwe6SMFusVCFwMtiGNZHrfv3+keStqTgK+8mdMYtdrt0N5JqRpz2zXULm6kB
MrkjUl33ae5Ey27/bLpn2Firw+iSzCgiDqq3gCokRvzebMA31zkdqGluXRRQ
2Qquf0BrAqSkslkg17wQCB6MTrm6LWt4V/R1aZHvPvrB8iOSxTFYi5iwQa3B
8ZuOfNDmk0eX/8EjFdXWizunnHaGKQcSFutCQQqO7PVLliR2GPWR/vkbHIOl
eBIHnU04ASHbL79o+TkghiXOZ5GJLwQt1cwqzOKP0bFMCEpOaiLDqhnUPqHE
UklJ6VwuksWvJT1tfZMDB0VXKDn4m3xOVky9Otj8W+vUr7n12d/jnBjcLCwp
2zqRGVauBdtxUhmh3ygdLLY2orSFSiCl6RtC0HoOsn7eQoWYAlt4UOibkQW2
L7+ZIJxD8XI/p/5uquwuNB/CmcbXJOj/pXw3FXVRvSvfJb31djgD1DBtDtLW
U6Sbq6dBpBz0IttTQy/o2aIf4mk2yZh1i8kg+4ovUe8EJr31Yw/tel+mKfco
1eLSDLwnb85ASNTay/hcL9074C/Qmof+4I938ph0rLLa3Wur3v888nt7Yd9X
QlJFbG2uEssUGC+qNHt6+fRAmRc5eLQuXsARIhfTOPlMQnwVAeD6ONryEVtU
Oj8hLkE/ipvM6Awv3+KI7XLzJd7DylY9xpKlaoIoYYRH9DxV96nsA8/LhQ4i
v/kpwWkiZDrCF2TocdUIkhv71PYQpxQuAwwidPGBC6cgLQu+A0Gn3MMU8758
IfnzGUm8YCu6SuSx6Nv44eAMIlPUTbB0oZa+XWNQhPOWC1QNu5wXG/Die+mU
9USjUyDTuUljrbdg85U29Vfew/rYtBz3BhQtgyJ+3nGw3+H0QFs2zlWQ8yUJ
+0Uvn/1p7p2EIQJwulie7xxAi8uwEPaAI2hBt2eDiFagfX1QdsIqImgVOR7o
/klZsvgqlb/R6FJ+czwwRLvFuui/+LCJ1WlnRMaWTlO0k+3m3uoU5ZjumZSX
nOk6KFTDslQ9nnD+H9atfYdo7vS4IXv+hpqb4i0EG6POXK3oWZrUcPnIr/Xj
so14L0pI7TRI7KxK4i67hp/SJQeiIaGtyCXzmC36aTVjLAi1BTri1MH+zlbv
XJEWQGCoDEsRZlWBl+cxjhpgfSyn1aqbBSrklMWDXKsjNS6kTb8GT7ErRkFO
gg3Xwv6N8DO0cdgGSv7K8yZ15YZmQ0+k6Vc+csF4gMTIS6s4SrjSMHXuRpKV
Hpc0oz1HkzHUNVVi1AwUGSY6xapAtXfUXcPKLhdR2gB60I43qzi2wQ8XkSNp
YARkS9wRHYOt5vuiWsDYvWaNoiLovAv/6oRXd+K8Zwuk/j+0fljOL4JU2sfY
TEp4dGN7j8U2ZorjNheUyjV+66DoVUXduIRugB5dVLp6Dl8hcrX7heThcGGj
DJM3ZOn8nJxtu86ZuujU5+pMzBeg0RqCZJfm9qQVqDs186FJ9Hwyegapa+TD
Kaegmt1PZ9q4NTmCKM9FgyZCJ9HxNR3QwtIgak6sVEGiykMvJEjtHeOXG8L0
35e08XI2rpOzTI3jQXiiV2kZT/H3gPG+CIWjcTRwJ2aj7DBND9D1zoQ4sCA5
SthChSObpd7QLecd/bfm/dEpOxdJm0M2VwF7GknEdZm9jrnIv5WhpTTE0wCO
YYZ666Knj4XFlE0juiv3UtFLbU+7v6jzD9bFYgpp+PnCIi5JZsLZgS9yDXVm
71zi9OJE46kh2AOwiIaoKQseNTjbAqiSi+RHJDqfSE8PL5jWfD7+98vWaFG9
/dpIL8PU97KyTF9BpvNOa2N3WSVk5iCGKEe8dkSZHo/iw8Sl0yzt4tJeR5Ym
3SkWbMb/anr02EvN/OM9+aPTwxGx0Rj+Q+anvRVtj6CuO6umb4dnWaSCatXP
f6GewZ+QU53nP9GCZw9qJHy3bweumd9EffExBZZ1VGffiFWYUUDaIA1zWodg
bOurz3QUefX9Pf1yiYW2TBUIAtj35daLOiO5lg5bfzTEHUv4Hpn4BF5xYnUJ
nH1JY2WL1Fj1jg/Fd7OVYeUFYvjJPlyNfVrGoVf2iGVZ5OZNoEWzgaVGiHLN
n5ShxcdC3ZpYy6MJPc5J1zRWO7PBqEOMMDfC4eS2po2QEWwEk2z1w7HOk2ts
mWKAcUidsOlUWlMgnJYiGcFvI1pl5UEqX7/H2x9ZWXtzrvv7VF+LeMxbSaj6
teaDso+mP5IriVcIQEIscuWJWk1Hltr80Zu+EjodVRFn2EOes0/SDOBa9AAi
FWVJEqZ5oSkgJrwI7i4n93RdRdvu9AXYH/te5CFEeKdNJ4KVH+1j6RJA0YFF
BXUDgQHDYwvNVaMjrSKCmW7fZupYnn81up4V3n0/g/EVGWECUhUhGsIVXXrD
HAK9FpFam3aWJAhkwnbD8QdBFGg6g9+rwF5GbYwhKbq9qGDO0eXFbILRiX3a
tGiZFXEmLsq4PCSjnUzXyDxoJCZWSu0LSeVAZL2mEsQxcikGQkcJcHPyp549
94saEB1pcJYXgnMY1pD99pDwrjcBy6R8vA0LwvmE4765r1rrWe99IhdC+Hue
+MmrwgIyWVZSV7bOJIQ5vqyfD1MV5x+CuYcdUHioFtpsUYdhXXm8tZBdDJMR
9sJ6yF7yeSGaaS0pmaI/SjgubI2Ah3XMoolGNtxdE/p6nPDii7tqZY8cHNVu
hudmw/QANTCeF8lDH2ibMmZ0qAdEtM2QwJp08YRsWVca+3axoY6kZWMbEfLT
gyz9MA5i2aR/1IRb0jjU9kJrOmzCdV6JZ1AhzrSOein+gNNxL4wpF1YbbWBd
PS6k0GgYJEXfI6/cYf0L9RR79Lfpc4Ouz48tQe3wVAL1Y0lcUS/nV2duRgZH
XAfh+IBTkFHFYFOqYrOAbebidIoV7ebU0/OJwTYp1SqNZwEF8UjjCGImVk0d
ul8THzNKnzZfLKH0sdZvDyr6FebiHrfTuJVavMcQYIRYLOjqRN4cNug4ZzQ6
0zsDbyQWr9grhqnw2PMNtKuiglbxVhk2+cn/CyIkLJs4nAOCouJ86UgEORdk
TdNgkiaB4Q3s/px9l6D66Wzg1Tbj2qMG4xQuHXLyuMSlrgLQKuxgmfie677R
49j5MHmogAJd7TFpZZPDf8TfMstVdCKJkOlHGgevfJMynDqgqqEtwhCeYD1y
UiPux76vwnkdKZv4G3InpH42DE0pmqGV0HI7JEWwmHx9OTKNnIfK329TxkQz
1DvSKN5XTpBNo/cvVpY+vDwwlpxv3YpfDx4RGZy3+yKs0wmgA1r0l5b3SqGB
X65XhMbcHVBsxqqOWjm4L76VFtvJrPaFOnO3e9998l6/Rd5kpYwzHcZsc5++
gI4LrtUYMMMNnED0JpDa9gk/UBvYIH2u+2A1Hc9peTnehcgajCJBOiEhZWzZ
QaExZ/FwWG9VAbXQN8+dLRHMtCUv2VAof4cAaZaQy4m94jAD36uI1KW81s0k
8VMyI1zij9fGjahsZ+ybeTX6piFgX7/wVgY1CjBlfuOGXXs54olSu0kNCqro
gcn3SDRMt1UYQnQlm1ILah4mFIW6BoiiDUhKtDrTcQkO8vrVzb9dSru5ieB6
sVSYI6OX5veB/tDaFf5xYzhCTkWRKVr2xVGBuf1ZCiwWi0K780jFfrxuzWpH
NQ2oowO3ICbnaUUNigbld0Dze/MPpnizIKapC4IT5Zv4HBtXi8XNVZlahhbT
MQb8pRmHhaOEsOKnN+cYcboPRRs7E0B+Gmpa/21iB3Llx7aYOOidRHO6uny8
IbyFWP/3sRe+3zDzIN87NGN48jxM6qEGtNMx5F1GSkrDnfLhAmie/SxDyeDT
5jkWeBbcwL8AcumFor1tKMJ8izJET1iA5ml3b071PsliLOBxL/u3kwIMRtTj
AiWTzsx+UGoJUlKxwQZ57L1IVUCv0ew5NXfTOSJuX/vMRrek1NdQAwvmWnX1
zRBjQMKVaHn8/KukjWGm8zKajAWDWY41qF5SZg+J7BDGlFzth9XRUU3hOaP0
NnUKWkbOa2OlvDJIMtuKqy3dEJXxywVKF0fTUSTIkF0n+J0coMZ0L0FJbjxy
Rp88EzZ/Z3N4GXeenm3l7PSXsDK+Ze/XtRLXm6D/d5R/ZJSx9jEZUBtc32yK
0bdr+h7G0N4hkEldthtE1D8XMMzcDgjvIJmjP+YzvYpFeAvLK9a5TzYZPVNE
83XcY8CxkjJL4RUOHv8tVhS3D28KP09c90JYG7wwqZVC+53iM1EG7H8PReqM
Y35tU7Idkw3m/gHtOX8MzO6xLYPliWnJvJQuUDkJay+1E8BetCapEvQ8xmDi
0KCTq/J8iN8bS7WzmfoP2BHTkAYYDueAnQRtz5kXbWMCzor6rYb14nvne0ro
LZW+z/Mc1WFuhRwtabr3aST53iShBcZZijW9rj+KguluNTkpeXyKM6xo/jNK
LTZzu6MnZkApK+oZU8KRze6SP2a4AS4xejeUE2zTKQEL5IUMsIbyExZ5NVDn
AT6uBP0w7WbKBBu4+0TqfsEXjxB6vzH1Sh2/PsWsjGCoRUNvy9L7jqwGf3eC
ELKghbfpm1q1IBliVxkPMaOD0dilS9kD7trpj+Bzhz2DMGK770xHjY15z+n9
LqBDBoxPy9dzb9TrETx0/0h4o5wn4pMECyG9Zupxs88KjeNgHuQfplIa2cQN
/dNHChBZgn/hZtfuD1Ri/PLzAGrdDoM/BwBv9M8hLd9i2S+KTdv0YMaFyVQ8
9LO0o8SGEZamJe3U6r1Yd28es71iTjuJWm8sddETYL2FfvEcU2qD+uWwyja+
EAHmlB2cTM9/i4EtwZUPYN6mzA6y8m5tGCEFUkjIPO0IgHx8s4SpJTLyd00d
zlagQrCeI3PzcdIVeHsYjOzSWjL1m3G6yqU89E/7MpzO/xvG0ktsg0S3ARPC
Vy6ga7lRbLgo5G/21QaHjDC1AtRQ47zXD6ja1+VGFt6uIs4VWFFaT4YKBDkl
ko9/dXht+yhFNgFkVihS7MTwNcpML7ZJBsirqvsqJy3Wqyk+qjXunRIk/Qsh
XUbW3c4kg6cwAyhoxh1cNDskv9F++TSqmcV+/OkF9G84WHggTNaO8gDxOzVj
7bIrEFwWaUBciKUWsT2r43VCfg2ehj1xV/dZMU+MlB3B7NRnrHdoLDg3Bpnm
PDWvBmxqIRQS8U8X2YyVAHtR6+JMKFfWSD2DVq/U+6I7WEzmWw/YK8zzOJFM
hSrDZNNa1j9Ygui9lSb2W28wEWdSoQYG4678Yw/mjfoxYS5+wkGevVtY+lt4
W7oMVyaWcYZntRpwaasaiJqxDkYW/PnkBE7br/pzxm5VQANWWvxWVAkli6i/
5mE1iY1/ronllj5LvrNcONNK20Kxek1H0L7zSkAQs8zeOEqWi43QR5eVvH6f
tsmUvCdql8EWwukrGqGfbFNoUM3j6bonPu5iaptxw8DqNphuili2hQ7/47KH
PAJlXBvzST7T97libDnnEmFbPwuOSiO80JNQrtQdNuixU5cEzLykkMYkf+5H
MfvkLuDiVNwSIql4k72gHd7BAhDxkrVSyGcvK1IpASrrXZ/Pv3dl6C2aKbK8
2QH0aNka2Vt7qUqBeWZpJigPvatHpuuXoCmOJkHbyZdxBerSOV6IEk7jLXjR
oj2iy612hTqSt1OenvCu+VuU34+3iEhqlT2MPpDB2KMN83dsEQqpZV7OsubG
kk/Vr7NmTraif4HN60kYbgyVRm8x72w7Xo9rcChsm58mpkGdfjEbTQ8rx8Y0
oZv4bdjsr3fOPg4UKK6XPVvgznsOEPGKJniSVSx6NptKT3C+0+agGa/0qhJv
ee7jN8/7VLBLmFgdNnB7JIViTvzD+8YC2uAWSSLy262uBd6WuZPAgYPFJlGe
enCu5KJOo2aPMuE/krFEjgPqIi/FTOa0vQLq6L+5xTNfsRWG/SIiFtRUMeaI
UvHaxZ+O+SAyT9ncQ+QXCx5YtZGYA1syuPMqEGKIgLLl5/rHwcLdD5Q46toA
1MgavB4yXtkTS9LRxByz+MbFijV+aE0rHg7dSwS91sS9nL3WTEbz7Pupv/Z3
zlBNawpn0kBXoJ7iDZR0THfn5ffyq2+sb14c6Gd2lHHArRmNh7QTZ+C+D8SX
ZSgPyHMjVSlWmhCtIoq2wfDrh9zTeIHAn5zDsITHZdwlXqEhDCxrv/chbUIF
eFICe773SwwL7wU2J9VKKKAFPfJorPsGvmjXBT6xVZtEm64xWbHDCZmGXxsy
fHc4CA1+IbtKrtXEO1+nJx64HtKX9lLkeYFiieTajEjHfRiaRxjJ48Fbuy67
Q2kM5ztY0lUTLOF+SqU67Wa0x1oVLo5SZkhhRNryfbXCtS7rOYsXxQQMzVcm
/ZnO8YGSU7d4ciEg7L4xthkJtAExkVpkOMdlG6Mosg0s8yxHWKEKuO20//dJ
LjUNt3Bf7+uCyvgmiydmNgeoRbevS2yoRKeHgBatUEaIjhBoTjjv1z4TdEWL
wQQvTQs6FYvAlk8AOrC/CXiYLbZk+Soxt4rOF1kj5Ipu/CPqQ6NKPnbemKrR
1cy9bxfZ0fw3UJwJJXpNJLj8HR5yxwZc2cR1S1DgiHbStX3HLmxeNLIf0L33
0OuCTWDf80oD8TLZnG0sPhBSb6yptXVylP9aQkg2C1YiBEQTJpAlsmmpej8v
6qhJOiS7p9kZaRlNSwcpGbFJKDDkpZClmEoQmf7wqQaTJo6SJKeZ/9NB8uio
gBO0BtIeBoCu4WH0y96dhLNftguk37AjWecUsq3kp707orXAz+kTGzC96TBM
G25rn+VZIgAWHgandLcQwPQ1LpYSzGzKnkXbxoOUqUYt+f3m6Yh5lJwxAz9n
2zsKCjHSfAN35+N2B8+bvuNgToRoFuMfmvbZSZXPSo6EI3l+yZntFM7mqXfg
0WXxu9CBZUzY6XXfBOg+9iqtl0dQKeqOh9MhlKW552MAQENRQLbEcDUicTpf
JKrIDtkhKc+ES/A0r1NB+gBYO32PZzSyGHv/NfqqGidi4qFkFAmw3k8BjZ+Y
yychGqxmnrbwqS6iW+oM2iopMm8di2tHHxrFiELv4NJzBjZbFOQm1xSWbgl/
Klv2j0ujosN1gDPD0bQE/F3knnVkHFZoRtuunqf7HMNkpBzpzZ8M1AE2vzZ0
zS6F9f75yWPGoOGw5tXpTeXP6C5APcX2wXu9X4BxFQkbpet51pGcYtWNc4/W
g1T1/e7L5VZ4NonVEGcjw/dihuoNsqcd3joiL2o2gIHBO6xILzczUCaZ8iff
DffL0/yd0WLXrH2Ld2OoBIveVLLHY6PAM/8nnTvW4eQssIKSUx8O8XpX/yL0
wmjSbUv+r26evhU8Bs2hWt2PxxSrn7DY+Y2zdDWfYN7NSK8Ve2/liyZ4aK4E
EveqgoNITysSv1gjehumjJYhFIKV3JjnapJMQ6eaiId0Sjp7QTzCYmg8Zx25
hXxQVWJeeiyx1at/JPnE7fxFkM/9W78QAnbrEiNWDtAvbeT0wiPT6IbCp0GX
7FGDqcxCPnplcY4xuvpka8pIVZcEiGM6elKkmYVTppNUO1g0QhItZInM4zfo
OGRmx+NNVbYBoPMg7F2rqduecrwJyh5kipgYKCwwCxPZ44WfJ1vOMZrW1Mc8
8GYpEaetF3b56FhmNyW0LTPgqF/K2OZnDbCTVtx5eZ6z/+cRjtMluDuVnTj+
jhJNIVBTWCrhJZLop07UO4D1uQvwRaze/vdmwQ0iBKZmiD9YEzNjyUTXUr4W
XUVyQOPPhigdkJouds2yRtAXw8dpBeLMVAWi42Cnc3sPMUAQLsbr7aIELlK1
HEgpCEM3USEOcs8gFOJ9bW7yvYlwSJFAhm8OytipA3QjcNay3U+yAa8LdlnM
r3Z00V3DftCzbxECiCFgc1Dm245s5PXsQTjYwjt/rLwvM7DmzcODEFQAxq1U
v4dy+ST2nT34y/8LHroxjl/+XqCIOgQ3U17C+HPEZUVnal9gqYPzdeByKQ2k
LGc8dKugfxP/hzUGa2PDY9/VTUY195rg8braWNA1EY0bCbv5FTVe2lwIoP9D
7hsK2og5jt3lzS8RbHhrDFhkMTV2PCQnauDvjl2BC5f907dqULvhfEyVCeIK
vn8PI+PHiAE/VktuVS+RTNkWOFqXJiLRC0IYKuGxy8cE1ZSZGdEMZY4juKkw
VBo71nolvl4yM31PDQMforiPZJxRw2YZ0sDHg4tD/2SgZ//efdnpn5rCQrEX
2HMFG6ZPh9y24kI19NxSDBYHhtWC9GTJxDj/Vl5ah++Z/fvdsoY9n0mtpZE1
FEM1e/GPKUAOnd5FpffUtU3/9k8sD/hXlYf5Ba1/YwHSGEGKa4JQ1WF2nJQv
tbNeMOLyMf7B5sjJGIvw5mK+Qh6JETe6mxIrejaJLFyXbpYFRsM+0zspBneK
wKlPuUC1yyDMdvoH11y3cZApFy0E5S+xoaqKEB9c6Viy+zcCa1C4QtZcvvWw
u/TRjfxlNhnvilzFUewrUtfHv+6mwc1Xf0qE+a9jXq5n58yBXrl0Oeymrc7o
NF0u2k3vp4BeeWsXQEYMcl+hUJafDDmw9htPcUxLAmFeCKxfvPDAGnooqE9c
6D+/ztGcocGy1zeExaGA6RQB/PMm7hGFWxG0A6QZEaht/QLrVxu3EbOg6qWC
cT7FAtL0sNFVNgoRwqgHIqBILa6/r4YdH0eljL8OC39zutXo981pRBK8MrNP
xuTySOgmhk8qF2ziYscpIZ21P14LGfGLGtLZu1iw1ClL2vyp2Jc2KrlSbcPX
8PVHWB2B5VjtR6yoADchST5P+OawPA7tBO+0GRe9Jq2hBdVs3n67omIv97Pg
pjsVm9f+FPG1o9fifkQY54ZCUo5wM8b8baRFl+yROx9axmsa+mlIXx0bO6Nt
hnvtVlGQ7QqLQLU6gkdD4GeX3K4E9L5e3wcxw7rGVFy/+980nzi3DxIK1ICz
6x/wPgLx/Q+cTWiRo9oCpN9h5fn1dOiH/GCrzp19cjYSYBely6eP5IkJLoP8
p6hlwSXYCz6Va21Cz32HVQ++F/zAIqQM8u3a3OKH7qwpwX1uEXpl/f0GCIGx
i929xO/ufU/6Qtvp3lmE94+wEbx74UmpLeU/Ftch8KxR7Hzjpjz8a71k0cs8
1MbNgV+EKD5Wg0j47W2gLa4Bfeu/m9tFVOyvvObuhpcjauuGq5sQ0M4CVR0i
qch6ArYRdEgZ1zRI159Y0D+nNBPUZ+nebM17io7YexFcddHViHPo1G3WCAKH
+m4kUioexJ67O9y8lwzIeXNsSC2XVcVjcylRSbAGuwY6o89Vz6lQ9Ae1z94u
/YXvvnxUW76NGa2K8WNRSK0vplntCmYeZY7zVSrEZXQwo/bStE6V4yKzyXS/
SDRHeb4F/TreyV3WZC1Qz/wz+QxiQfAangnwGpVx/YFPTTlHJMjtLBAykdC0
s/bQlClt0/aQrVltyIwyFuXqleG4Mh9eGPWk6HeZ7DZ6Wt72ar6fx2BvR0n/
K9d94gz0hBBVkFIe+M4jAA29TCBYyxpoFyqW6BhjswhwCf5u9CGuOT6ZFTLE
aKxhLP5zBVJx7dWJcbiTVgDMFBTxFmX29InQAoGGwCTZvkJeqx0r3xIVtuXB
TcWWajsiVju2mGQKiQY0u48ZCjHQF9NwEpedJNsrzUujOKyXC6vSEQ+vXZrB
0niyzNmx/7TeE8mPI+kpNzGdwgUJtNqAKbIF0pCVegiUgoxo6G+mQhQJ4GNt
/gRE79+EVGSCJUk2Z2VzH/UfIbbmWs8s051TDi4KD+MYxneQedT6ZlJjduKt
xbdqjY6JZDaPbXYubYp6QIkfbQYJP7KOBFluBybZ8HOTf2ZQFy9jy47xdIzq
YWqkAtyu0ZCaQw4nJMVY1jvTH69IdUn3V7oj6mATAgjoSZHKJqgHm0LN9aqD
eQUbQT/CALy21C+NWnvoS1XF4idWp25j252gs0Nm1xCU/YGHfB69ldUR4dAw
CmExJbY/SP0iXLqR3ZwWjw+NXXId5eGYznLx9bQjMLdRhqoqsQX/NqQtoS74
QKyCgafKNGZiYM0oDwNhMn8YdJ2cL7mQXFW4IGhWsLGXRoZbhpcGZjvtksky
LLBqk8iOV4HLoO3dyqAvnA2G7XTQFPZa3s+xpVRSRRxwb21FdXy89llGw3pm
M57UPOcM2ULPPGXWVP5KBKmGqBlfCi6lbnFuc7BEPOx96HhkGhMABinCsbXj
joIDoDSNkwf71VwJ9pxsEZQHFzi7pbTSkv0TUpf3FGuF8XBDRfII1V8qjmDW
IvR7wolHLiV4snfnPBDlZoa111LLtDzLU+6tRC8JnyO20pI+cj9RO2yXcTkA
o12S83+Vh5Q3VpLdvNf2gQZZUJMhpQCvuSpfVgdeKuO/6koUehMoGHeetkIV
uLk7gVe9Vd0+zXOW5f0Kbduy0SnCj/4qCfn11QG5M3jLN98WV4GK4kkSUf90
lPiEwzRJCUTdQ8gqyYFiDhvdW2F98cXVyBn9XV2cFJHDgZ7x2utyIx0UftcT
PXC21GJW6WzeUEHcNxf5mDYXtPLBESlsW9vJNpgOugIdF4MClnu2XwCS1fLa
xTL3bEqKbr6RhaN6NKvvt89iHQ+u0AmQlSmylt3V6SBacyz1QldfjRLzI2tb
JYVBfBKaqB0zo2sPosuH19zhT0aNqdPSgRo/r+O8XM3OppO8fZGkeUqNglXn
PsufHENsEjG+MjDVVJzKdj6olXuGRIRIayCsxP45D3Y9ME4T5kgeBkC+LdGQ
htN57rVMt7bLXfrY9j17LJDbAUxUcPivS0D3ZC8UCTXrr1exZHIKDkzLAYLY
czOqnBRUxyzK7KDoUFelwOIkaBStddvu0cu8ETtXek/+y0OWJ+Ch9nhIGSWn
s2ddkDmIHQktpaXpOacc8kEcvG+BvJplaDXfTxq+S9KXQkKkcQL8jA/yuFBJ
4Yaib7nlB/hm3IzPEhpSuX52AoE6uXrJ1dUnQZu8prnhZMlcL0vKf1nlS7LY
tVvG0L1m7wkdC1RnQGdOJI+fnCGD2K+VWZu1Hv6ZWXXMuTlAdvIZ35cn0mTo
Edzq3BRf/j6KVntLeRZ/LNazsB123B+f581Eb2sryNhFLx/3Pqv4QphtHCmg
BE3ogY4VTkRTsnJurH0jdGt0L/sl310f2hZEyZm0KEO2vWPIM6vzpJPn3pnH
jWUvN7jln9PapqZkE2uDrCtLiqJS7Gu6GI+mMDR1Cz6hXiu1zvkZOMWRt4mG
XcEfRWItvolrKGq4EEM7ARUrmAxLZs9C5ehrSijzJhfHUc/1fAH/jpbqEgMA
im1hpaGIpzz875xKXankagi5hFnkkMv7C9Yr3+LcPToZuPK8bs1UvfKonnib
E4SRdsu6fzw0RgrZdKkmop/PVLux4oBkJ48syck8kG7LEvN8/k6D/WYuwtQL
+b/llG21hi+6kWBcTmCwCssxOL3v7JKZi5yox2GzQ50XMrGlf03eDEc8ZgpY
yMdH7jCEwiZIZjrFKAwn4PE6vbDHS7GXONu/D45jCf/UQwyGw9IjiHDBf6F7
Uj+q6O0+X14//IQjKnrZ3QniQu9EesVBkrERiNxo1XmSznLXr7Frd4govkSj
xGKm7GGv86WuWDdBdtwrsHoqGoNJwBUFsTQsw67FhLoswSPbEvNUsOxVl09K
feBL2hW7Up/pkUdcI2IuJGeN6fWa95AVWiJ1Nj8zVaSTE71XIzkM1otfsuw7
sc99ThMrGXKW/+J/ysrKi9CJnRphW1vroWpUvNpJwuZb1ozz1RbgYqOWzQL+
8TbUu6OjylT1NuKItR34j1tTrzPnbPavn84CiA7VB8tsu8xm+5QvxNiWAksB
edjq69QSrBq3fT32TnlEpCAcyHRzsYbpLG8p2TfwxnYVKsE/lfN6LHIzycg2
4zXwfjuCPxWP976mnWW+huYkHxhOkTqBPxti7KkxmfBpUwNFuUaj2GjwxbSJ
1p/DWu2+EyZ/nCRWcOjAI4Wt1D3aaVsi6LLPe2CihcUN3Ii6mk31LUAZGo79
kQk+v0zJgfmB1M6VdLmskmo=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3GEU0LGMncVjw6v9BJUQdIeYX33fPTQS0lDEEkrj/v192Yhn1SKJj/Uwf1qL/Smp7wWuFQeocLIEVFqqkcvrJ3wLb4TZc+Qx0nxwz+otqmWTrcaoZcTGwliTRGIp7+3Rh790XJj8EBixBG/ndaoGqt9HSDuRHjPXL9eUybY9kLMAcZ8GMp12ZhWxZHJcdxQtjLitRb3ts1gsg2sE4LhVp3YYMQJ4gLPtNLHi6qr1b9M7NVHAG6qaqQxfZHQSCaeeuB4WxqoxcNr4GKk+rgx52hUhHf6ZDK/lkO5/093lqzaxAF5xdKqfGXgh1P38wyv1fgkCstoJtLHvL2WLt32I8BlMYkfTU1TefpKs4eatDVADt3YXcW60cvZd4II+ptydtqpu7m+ybSqq43/HqY3dkxautjPn/dlaHEQyq12U1efs8R43TL7zG5vXsZekzDodeCDPRtVJFy6PIBYSOnrfO2PzwWgNKfLFHwyY7ibsJqGBxqxstxGwLdgD5xkz/YJCA92pcxLR9y+0nzf5MejM6akVWEmxopXig/2LKdiRi9IaTLEL395beC+XkSTUaDmq1XHi27+x3Em1bnt3Fy+TqTsXoFf3Ul/haNk6F1c3Wk2UudfBINP+YQPAQufwZ9jCJPbA4RyuyvLbu1Re4bU9AaBgxJONhihITNSkg9iy3tpq+8YbA9wAGjJhFZQEuLF9WlRnqX1VAvlCUE5A2gHLFxpVsYdBIOhu9+n+KPv4iGMJ2BM+qmDHWpgNf4CWezOOYE1IDtpYQqG44rKhbVppVox"
`endif