// system_intel_srcss_gts_0.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_intel_srcss_gts_0 (
		output wire [0:0] o_pma_cu_clk  // o_pma_cu_clk.clk, PMA clock from PLL for proper calculation. For simulation only
	);

	system_intel_srcss_gts_0_intel_srcss_gts_200_bg3co7q #(
		.SRC_RS_DISABLE      (1),
		.NUM_LANES_SHORELINE (1),
		.NUM_BANKS_SHORELINE (1)
	) intel_srcss_gts_0 (
		.o_pma_cu_clk      (o_pma_cu_clk), //  output,  width = 1, o_pma_cu_clk.clk
		.o_src_rs_grant    (),             // (terminated),                          
		.i_src_rs_priority (1'b0),         // (terminated),                          
		.i_src_rs_req      (1'b0)          // (terminated),                          
	);

endmodule
