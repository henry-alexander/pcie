//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qXuujMIdDf1Y/tWzYNk3Gsb9xgvvnRkx9Si8/El1wnk68XPUOYpMvaeqBvII
sAXyLYftCf7A6+6p1xEdZ30yRhEMYypg8ghn1zYbjcps1t824Y3nOk3yhOm0
w8IeF/lE/msHFkLmpRocHCcq9jQq5KsFfesQo0MF/1QwF+ta/Pjo4QI+nPvm
621CFlxlsbYunRgRAI5wXJm36BpeqtKycEDzpq0uZAqG1S1oieE5Mqx9Sjt1
xBNNkMQVjyQiuP8/mfzyUoa+Gme5Z1hcSR8OvLaMgsS3RsHMq93jIPzu/szW
C+VNc43FW+N0h7cRb8Oii/IGj7cbnwLPGyVUZxNEmg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nfIZmFPF/6KoIsp15uHufbJAMI/12/zqB56mdMX5Zcvmo72CNkXKdxRaEBsA
6A38WgvXMCxR4R5Zu1QCI+ZNJUJRJiuTUo5T5gJ774nd86FQT9TeY+Wlczp1
wL3zC+JwoLUyDLSCZ2fvrdZfZSGmH9kociOo0IYKC10QNKq9xg9SZmeyEMm9
x81j5IENGbDvDBTROCmVCl1bDdpn9m5BolxeujYuKOh+vwi3+R8+8tBrESNN
qnQaR2HcLV3M5i6TzD0Lv2eHhqDX651/8OW577r8hYsAC21MThV7cqXQBxgm
dMzRpjGiEGUqoHg3xp40RKhSkF1ez+xG8296NivtKg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
i0YcoKW1zxW9urI+iKiqx1c9+jKyYC3xc/Sjnj8VMR1Cx8x1sHufiv5Gr5F/
lfZ02ea6n7CpUHvQBsWzfb1LIC2OJHfGCkKSFopZ/Q4sOJa4n8A4PWw3FTYT
lYQ72EMXpvd62+Xkch3wS3/TkOX+jXH48ScEy4R6kk00XDc8JwvVXk0P1oum
1MxYQ3CiPJIIJPfIA4wdjIx47bEiLjUMVFq0GHLh7vVZHGWYemeBcHIoKf2Y
+IvVeKUo2faVPGwxVsbYw/dE34Lkp+D8tehGTv8HDKKlmpXIAFJuKvaALZLF
mh5ShxccdumAQT6WL4Yae1cZx1vB4zqbN1asLclArA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qorUyba/g2bnlh8VmfuY7C0Oo2m/V3X5EVslcCuUboT52ysdZd9EICpGdSTu
GfXzdLm7eKbotF9oaN76cYQEKHq1Yrpq9rIJFVRptbVkBohrFZ2HSId91w6n
3OWfZIqDEMsTvUQ5njNhv9mVpGnT5emjgG3HNwXb4PaE9XgyCII=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
S8VU7A8aa5c/LokGbDCZ/mnk6qXCPJiFOMSSSSXiPAVnsX52LWsZRTdudLOj
8HGxAwDEtyl6ATqKPCTavqshPijU1Wi7MTbgDV/zBmQ/83e0OSG6jXi7mt44
4QhQ6gJu/k83mp08oM1xsqUn6ljVqng5rX+GXXlZb6NI9OlxaSZ/w6AUqxfk
GbvKlQQSS027RFKsxA9rogtl50GZZR5aXhtaq30ItG14ep+83XDDtrPTywgd
ncoekJJgvdKdfabAiMBJo0tPlkIlCCta5p8fjS4n6QaLa3eucg4mPRjjX9hH
oBw4S6GbfyKtf46UKjLPhOL2HFuh1IOzS6GbJ6tPV3ySIV44w1PHSfwG8DGA
Vd7a6iEm17PQ7GXtBZiUUv0TUC8NoX9ndkbTTgqYb/Yj/ajusmQev7n9v2rG
lRzzh9jMe4sUNMFRe0hpByAQHPCV06LGkg1bz94XkRlm02UI7TgSEpQQ7yyU
AvyGq08lp+y/O+BUD31oxyYMFd/WwD8j


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
cdUIyFQQ7ok/NvF0cL6Sv9cCcSkbY8xxOCPIC2o7MXNE3iUcTqM6doXQDnsI
MKnmHV2D2cTqqKiKIX+JRNxYikpX22Tz3mTOejTLmD2g4r75TO0O5iu5WirL
psXp7nEKhG3vzwF2gghCZVwHjCoCXUge6JwyhcyILdacyRrGHKo=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gRIrKFM/SdNitHM9G/cQXvyhQ+1SOZZZkESCGGEHUULFPZ+1bzUXvMjY9ip8
V1d81NwZFEUEUs6cOunwYjrampzOyzz1OR24MrWXD5rTP3UgRrvxTp/W/UTa
mkzMoWDZxYFAkogev0c7lZLdws9V/Rfcwfw2y55GUlg/WC7eTXs=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 106448)
`pragma protect data_block
tv9UxpiGJzsWB+S3ZVAWI7ce61X98Lfu50POk9KeaiKcd7zhLVmrJWdURKTY
6cPtU1aU33COikP+fdkvxp3Ti5TY4IKMNhV0T/5Vu6fZ33NEF8gl6e0otMj0
ZwHdDTSnBlV8Ktxs6SBlKLcIDp4cuiLaxIj9p+kIbHt1QQAhP4e5g0+9a8sO
/6bKuaRfDFLM2YTvW/qqn3pK0qc6cHnZTuSTp6XW+ADOAnVQfFOTP+vahtKv
YroNx2u6gZW1GwqXqDDmdXBL5CdAQzAFy5RV8Sjjc2B8K4cbHYY7PUoXup74
eEBx7vvqH38VnmTDggquKQAK68KX888k+rUVNz5sFh/Ogzh11JLeI4nOBuet
qw7Z5ruV11LIGi3UPjnn5JM8C4c2IySWY2+92ya2f2OVgPY9u0fdB4gI702f
Vlje7KNXR/cPhVOgrMzHrPNvgHQx2qcQBlz+TRBwkBdOiE84DbLVSJ2Mt7Ya
G6pspUltr6crcHqWDw7jwg1wtYsdrKpdXYhWESK9oBsYgSyu+p7C8NMlrS6S
dajs83ht7yg4p71L1X5n01HhploS/1QltMlTOareng6ke5sTwwdN8MuAwYnx
t+srD3YfAwXcVK1maT8puzC2l6e3ZiF7VDoRuMUZJg5aLAt6PosYfbg89Oy3
ehaVhT1J+hBfqAQm7K3JtfG3k4UZQrdk51eHYa9opTInsEbcYZ1E0iuLMLw2
Kfy94u9rvJQ5bdm6IdqAHbDIaVL9LTR292lncQHHTGvAkj19ykPxMWkERClE
qcmTSAyt9S+K48LLY2x6IUis1fWCrKqfaC+JhkmXhSYn8n4yL34NOyiIZX8I
02KlxC3q5quRrgMDO4YRUFoBwqZi4wks7GyeeOZdxpLXVgT4rfBAccUVFNDL
rU06qZDmRIjVE6AtsbocCY/My21mbOj2XSUWsYSHmuLhQgP0jgx7gjZ5Vx5/
izX46uVVIrMuh1CnL7k3j2J22KHOWX1PqlHVLX4qHjE1xlUx/uZ3tlPR/eyL
cM2hAmm8GxZFNllS2kzd+uGDvKHNivYjJO2j6lw4//9nmrxhxxMOdfL4GYur
sa12Npm3+3WUIZikHbkpVAtYzReC7NA6NidQeg0aqcjSsFzdFc++TrdUhsSX
Rx6ymhTpneOUJOBlsuMSrOTHD4tJgMxId9vxX8lVq9nOxdBqU6iKPHEi02r3
QrBAG3LbRc/x+AodP7kLSCNXqWzSCJilQiT7Hx0sRmBoMwDouZWoLj13K6Zm
4JFoa7FBjM/A1zmvA+Qd5EDW3LsBrlQPcItnvDqUsDyqXoBxPBw4EOBMqRO1
dYpSY2pkP3aauwKvVSHcKdtBkDlMRpIHftTzWMSrJINnRHXtI+8C2nm9N4vH
+d0QoPzUubZAwaG/kGku+5bszWMY0xMwiOTKJfseKV+AGy29nMhHJhL/4cBn
uFsyqvPpPwNKB11bT1BrfdKTrOgmVcMcCDHq2rrpb8PvetHNtT9EJObOj9aH
Xks1c7pE2hWw7CGMte/7TVuhNBwGcRh7T3PvcyUP+Et9Qb6kaJYzzZ1bOBa7
RnIgn+nLPy/qXJmnlZRkMo8+79uzb8W97HDzZCUeJXduawsWISOHyb5CynrO
BWTXMOStBPDe51d7qHjCY3S2TdOG8Tb9WpNOkAcBx680iDb6vL49WwZIxFCI
IaGJVXywxnbo9zy8qwqXjyiCJVfH6MGMESFyXSH2bpZ4QZe+CmOvgQEEGbNP
hpLb5D4HUDvm5pvDVAggjePFSf1aMqjAOosmlpQisBcNfHzgtvPBav+riQ0D
IDFib85ToC2Cge5l0erknQRv7LTS4YlD+U6+q7i/N5pGctFcSxyE1uFlmdqB
k8RPIoPUOCBSiFUpy7H/OF3HRO4luPaaCe8CJRAVL6sgpXRDQvr5nUXahWxS
CZrndlP/oDJnENIhqD9VyuT/f9et/L10pQoXBj8zu1Icw+M2FuXIQv/8pN1D
myoKJaNc+50GayC0eGgOXjM/LNnrph28IfyCtP/EXIRs/XaDdKaJ6yb+xrcB
oYcuHp0OptawuS+UB5LRHSPKLOBo92Z2WDp98R7aLQ/wVzH87zEaixlVdNiY
3Fegn9QXaO5PRvb0zaVr0lNtQHZmLUmWtbGegwUrfnNo+2fZt41V+QRlwVKz
DLaKsPVRhgVI3BWv/reuuOWBiNeof2VIVUoa+NgpzsV71EJBul8s7L/M3HKA
BIracsnbSN1CnXMP7tNZEBV3FUpUkj1Rb5HWuU+ezwV1qXC8mzPvByIAa3QY
4TOd7ZBsvdoGSaNlCwCD/Jtcncr4bTY6my88hHIUaDSMn5NU/+ptiJlK5Ghi
NQiBvMwUYOtT0LIL3iOy5JqN+h2Mq+oxEvNzxGDJsAMq22jhlpev32B6OKOY
KydNEzLWwIfJI3mI3KxZsFw4FRbePMz87ZDiG4wIDDZIy977wnnfUXhrRP1D
tyBrk2uzbohNcD1nNfiA1HtmKTBfF7AT66JawlGb49A4dwfUjX2bKqkIqIpq
WZQDoCh650swP9pBxULHu5LoqMdoKQKTM4BR5OG38/zGT847KByxxiYT9cNB
a/fzrzAINaXtECNjiTRAOIfNcfMRawV/3CuVg5AA4tArbhf6+YKDLyHqVXcn
T5FK7Sx5BRyY0C1+Anoay6UeIlJcaHJAYMGXTVJVE0ebiV1qGzhYMgnsGo9u
olWIYznP2amVOU/gvJCdPCogV4NlLtHVD7qTJ/vnm857jtYpXr55Len+YCnh
DeKzAxmPlDM8aoZNihnlMJ/VMGllJIHWOWjWA9W7pOdETpBckrcvciX68I0V
ktyrpA5uMQyGzb7cOYPbrew5pAbA2ZTBjVpOmH8Ie4OxN/LMYI8h/fTjCGBj
siLnnqN3/M11CIYa8K89rRL8d7ln5d/S2g0nT6d/dDZjpHR9gFxRH0EhxYl3
KonygozX/Sz4yCyV0kk78oyMreCin9ABqGWnIECpwgHC/T9YqMAHyE4HnPB1
lNQ7cKIwnt38g8YUGrIRQjSJmgXMjBVen18qUoYUqwtBGpK+mBhzqPZUIJOq
THAWbU6ueMC8KZinIpiFQopFZGJSz/o9QYGCQUO01jkfR10iZdXSxcJv15fw
JVOg6e1LoYeZQxMD7pNyZQapYdjt39m9s02QdHYGbhIUppt/6p9tmQaUPSuO
bUBf2fvMwAuY3mDrhTbLvxyxvsdBrLz/B/hR8jsRuJseERxhN31NP5AE2cWb
X3C/TzgcOj+RzVdAMIb72L3s0BXV+PPqtZoIAgt05C1aSlGC5NeGwf7dX3na
OKVwI7PSHUBZbw1+K9cu1qhrQDyRZ0Z+v6tX5T/XCorp8v1DIe2B+P4CVHxX
HDIyN3N7ywSLcbHDWF6oFk2bLTvDGw4BXwEVXiOLOozbWEoFSWQ6pY4SlzP6
W3d+roHHcX4TBmrB1fXc3pvaJbaOr36V2zZrb2qsriObbGuOS7aivFtv2NB9
jfoGtnUdZaNmHgl720jrD3g+Pth3Apb67TDXUdzWmydG40Lf9V0ihua6/B/B
vstdzODuae80XEtGUtgqENXeelxGgf4piozHb+vwIsIkp3Jes5jm096q+zLJ
D47ndI2VgsD6LNH4Zgcuk3PN4mtRL3Z3Oo1mltbtameTMNAKefV+3ZSWF0ZU
ZLAGd0c+uLhZ94YHADKhrhjen50wjuVxkJOBW6d+iO/N/fxQuhxoag35w0iI
5KnaEm3ZQjiC+88Qp/WIcNrIPW0LPv7gYg1u3X4tO68VpLKwvMvqcB0OSW6H
ALrdOaFioB58kWfLGGkOikcigUMLjADzzue2qPWx3zeLg/zmoIuVW3VRbE5S
0VOD8CRu1+EI/R8+hTDVEa6qFKUIxVmcJq3pi7H+3O1dhyiQiLuA+3nTbML2
SCRjPX9sHM9J2n+f3Zajm4ZYuGoSVtCZWoImO5Lkd50Nm9SixQjqaBlomCwZ
O2aG9SnCiB9yufHOs9APzVSwh8sMWpBZjWo/1jtzVFNZVsPtetj8qvFCKoyx
fj9ns1uBDOYO+pRIFUqJYtWdPmQEKyzUeMrzf5hDWN7pITHM3rTg8qWySuk5
UMiyIG8E2fg1IYmJCS2fuI9PouuFd9CvkW1nxTVfLKuUdtVY88a+ulR45eam
awFIBS0f/WNVfQbTEF42WF4dlg54GFSIHjzvwOpmx5PPCIDooXe5rkp5VXNz
uEk0jz+U8ouZ/KQceF1fXuuzFNnaCG8mijN/dvjAMitf1eAy96GEvUL27N4k
g6q/B+hIzUzEzxtlcHoYXCFFxVAQAbtFAI58w83tB9iuGOm7/ul7O8HP+Hjh
CXUrcyBdfeUvlnUu5A/nC83+hRUBS7mhW8A1RZ2DZ+SZvm5E6DdPnjxca1bU
Z8LOKHFg4sm+RUssxc//xlxowjaAxxu6RT9qlHeAVj9INWmBuA/nVC88yRXO
w0lqhp8sPv6FJyOVhciM2zNrvsOgepiUJGigONTQ3LRVa0gnlTY75bIAwe4o
t4xNeJ07Bx9N3lUqFyadNS9d0LbAiP2Bwr1zSDDQFpkR2yLr2pi+QzjXR98v
jQAHAoAwbLLCSnWFjBHBkmzrdIBW1xhLqxtsl7NiOMi1xnQ0O7s5Gop8wyPi
jCrbdJnOl21SeQkFnnnp8nZaDtRv5WVYwgAMuxM0gS8L4II4lG5RU78nVn0H
mN36xjPPKRnOxVU92aWlFUE189r5/yRBx7m7Jq8vB4/+HO4vf7QWyi0gKW9a
twJ19TBv74i63hV1LwyNXdsTc5TPN+YhxNWKZDWuk2ZMrM5FNJtrr/maVFSK
O8s7VZmduBOpkB1wtXhkujrMLOqMDk6eAtbBC6oELIVA+02TOqSbJW2WaphS
UgOW1uVRtGhnlRLq6IeH+Si7Nwi/9dHuKVUO2nAIrwghoteTqvQ+wjOWE0Rc
fRhoIVfO6RYKl9uD824itthyhRBY6VAT8sv/G700PXXmFWcHdxiOK29I8t3Z
UYdmRAN/eTDbgM7x3ecJ25VWEH8AkXlnUYqSoh2K6EMYPa1sqc8te94EgVzl
LtfhuYiQvPp6Smi9ixpTRveNQFTWFFr0f4mmehQITbGDvzi8WLd+FhdWYo3c
t2MamYNTTMpvHIWi9sz08KcBqZ9BCOHA4M0aav9b4t0231DW1LDNJ24aFaWI
vIpnD/TSpbpv6IEkixGwvW6XFSPdqfiFoXihMDJ9HCVwMPkevTGx3MAHxg+y
z/XI3zKV5qbsXHNpfokR0JzGhu0DciF2UGCaWP3kdObX2Ng4HNPdZT8zf36I
YFC/FB74MhETb0a/G/s6x5JU/0oOtZEs3qvGgFi0l49iOKE4mEQsgFRJId0U
fFYYO24hTFdmmUpY3b8z4p4udtiRupqyZ5pR9PL4QInHWBGhC+PGrD5VMUKi
jqDlesVRX2ErrsbLXIBqgfxE8LgyH7sG5lnjkzb/nUQkXv7LLtAk7IlOeA25
q/iY2tytEUGVrwsQsUePyUHe0nwzmU5UzHbZsCczK18A1DzAusFQUX5e2R5b
ZvcTW2GgebnjR46PbgyJXMzJM9NQ36i9KMqZikevylQkMlSjlLF8x+JRvNlO
Kt6n+LOHt+L9eS9yilgaviFIPE3JLr7WRxsZT2axWFQvwlZtaDQhtd0KJWwv
wpqAkWoBv5DB82WTlPRlJ/zuybmruG5WW6LhA73zdmkeqwTVvyBYohyiBYOQ
qcEZI6s8UxXhzokvXumkqUsaSOamxbRjWN6jmSOWDJrtrBEZZwP+8xprEkuz
BuqXI4ADF2mbNyMKbgQo8s0wTfYQSqLiDB1uPupw/XUQA7YhTeVtcnxWD+n2
dA7HFTWf8ZnKe/RHDfVf4pc/i9WNVRJZfrZBOXtOtZVPFN+3mMerKwKb+jLb
aT7BKO7Yd56PYqtqUhKC0PoglmW9ff0sJUBDcTkcLh2hnYwxi3CiPexLw094
qkXduydD4KssWa5Lwb5owaqfwA/k7HlNhd/5Q/Mc47phsu2jqa0vvUX19CzC
L9f2uFB5AS8s+ULTBNll/r4idj0uCiuaoow4Jgt1EVPrJljoYfksG89Y68xN
cWI8agxn5i7FtNzzo0c3M2LbVKUcucCrouQG5LWzwXkUZzDxII8NF/shpn58
+WXbJu9LKQW+S8LW+41jBNM5+STNLx/T3onHA4c/GK01l+VUrPpczeh5YR+1
YCMoaxifmCUkDbhkWPWyKN2ASy6TfheaaoMArIKDsMnUiLauTza7CY+cJBWN
BQUHMM5WdoW6JUl+otri7asXb5uvzG8sKeN/hGnJjbw+XzlfYztHB3c8ii8r
jOTATZYgFdjstDvVzmmexDqU75C4wmeEv28MVVLEsgJQetql58Bsi+vH4LcZ
kz7DihWIeuEVHFNrNYW/pF9NxEc7O7Azj3Cne7P3DJE7g81zhnlZTN79VgRg
/HBHVgOfQCmloVs1n8bJHTU4geccIZSgMgCzMcDu5U9VcxhLxBEjmobVFcB6
eA32s5rDz7ex3JMp7Nzs+MtiYiovB97FCdKJdkFkuJamwtMJqPq1Xe8UqSYo
2pyhy97RhdR+897LCydp3GblCliqOWJ2LzmhbXHobudHAhUuRwmyd4RJyZSD
KfwUgXECgvB447FI43P87we3onyu0pXUUGJbqFCzudePZO7cqzKj9wPAivRt
Kc/sPubpqOiXf+JRaXT9ZnHesk8I5zkCZExX64ASPd8E8KT8V+C5e4dsVm+P
JZEWLcIUpSvNnb+czG+v+0Kff52/aZgzwr2GDup9g5JBsNNmo7rinjTV5YBx
HXsdMMhtjDk4kuTUfs+t4FtMF6MkLfwgP3rZ/jAxn4FW3Tu2XQKPC5uYYOJk
Pby3tE9kqhoI0QczaGzdX2OrX7zj2bX4fo0xL6qV8EeOMkwu4QmGcGf2XRqV
h4BgjrKLhE3iGnlSN/KeE+myBANKSRBcg4g308xckcofRIbOGCepggsLRpb2
inSYeHwqzspUYDURth6p194vfuj5ioQPwX8PfWzRlNdAqPqvUvleP3ji7ifs
IywO+JSy5qQ24jCV0HuF/29ZaIwu0gephD1r7nRiv5Tg5RNtZeEpQ/6C3TFo
4KsL4SaPVqoy5lc40NIOmHswU8IzGrZt4G+Y02lZhU0/ItJMk16VQ8DZyFsf
m+fR67kJlCl5XA7tMmaLY0sxrS695QyGGkUplGhEin+vPLm88z5LWr8BCbF4
6GuF7upBsClVHsM1YYeV3VfTu+1pNCrI6GlmGAPU34c8cEGfpcilLebsCNfc
16tZerH9egEPp9m4Rz9fRhUUoiY4DiF20KrSgt0GZE9mENAUugmjAv4rssUR
HqZ5AVwGJK9ocmwG7Wun+mBw2jguTuNwbPem55lCHBJ0E/bdtiCH/YzNvNK4
dAfwgZA4FBhX1SeLoZoaNJOri9rni2AwAf/hTNqwHvBkrQjwRiy2WdxYvMWx
I6yd2Fgwjc4IGAzTXrK/N29KD+hnskb8BL+gYvfAQxgbjWokLaKRwRV5RLEk
+cxA1wsuCWVK8Y7RxOtWopARY5TKLXeZ9XCqHifKrSWx62lwdCZmDhBVqiB9
3H+0Pdwdvl1UVcjEaO2k2+nzc1bPvAlYRcc61sE8w/3DpOxdVfaJsWgXUTct
Nx/LjZfN2ft+SIBinYhtUb1eoyN7AVCGnZg5UPZQf4ttMrdC4ityBWwv2hjK
7T0lbJ9z10T4cw9tIpKz1gPa3gHgGKNHiuN583ibdalpNz3n6eQqvuB7Hpo6
0wrcBLh9pC52aB51lEArlXIUoR+wm6//GUxQMKtCPVA4tx2IiqOygrOlNdzr
jKJTH5PmlxgSZ7nV5ToSvIeTJe1kL3ADUbNaI5PStguKc03rYh3B+W0h7YsL
Gd/ThjspFKbkqh6t4R6dHhjoQrtoML8cGapw2MVlai1znSSH2VAg/8CGByS1
uZCCsdQM+EEZqanIrpjODzmGIHor5G6+L4IwNpRpdJsBfItqkVLAPA+48Vwk
NbvJYMwvvbh7X0Q2c7rK3MCH1IL82YX49DoiQsCpNC604n7IUGgSy7C7wC9E
CFdsygaA5BxB8VoNHP+hl9cUCbAF3x+YjN2Ql0p/fdcZoKBfKrOay9qxp83c
Mhthx0TU7N8VhUJ+eIHkBXRUKZRFLeaA4xj4ctkyeTZBEpa+f2EpNADYwnUS
Os9ET1jL45VEpW/fmdMjHJt254c9KKCCo5+ARrdfGI9l96xMYBuXObpaFJ0t
f+OxUhfkHSWKGiecUeiJvrn3ErgrKGZmPok2g401gYWkbc+yh5rU6KXvZ0ep
kXZIbuwgFyKCLPBq2Tv5ejG2gevl39+6oiXwx1M7DQt0S+sxDLNqYq82/Ebe
xqeMe+2CR5ErNDmTMS2LaFHt1S6WhQjWJHciD8jCLWQYRQsCkJR/0utmcr0I
CEZEpCY4KwNmBhLz4MyWY3JCrvBYG1DVdgYMRmhg4fN78Ouj3PINhpkiZ1a5
nzb8IquRLuBfxB7Jcslzhnh7lXl7/hTEjwQlMJldOD92ieLwoIxSd/GMrd8J
Udw6VoPrCeLVupAV9VFVzcQONXNzvcllx5LTK3YJqRRIRzVmirUdZMN3ESgS
04Xj67LS50gjCRlSBeJFH4jtL8jC+YJOlWXV9KJIIKMpzOMjSZ3uo4+JOIUt
yefosR0n+M4VAuA5fztW7s4/oqSleINlGs9FyD/QeF6j1nfXcaTtIYEMXGdL
X36j9M9XWjDYryNe3+/kpfam8W4Wnum3R78BkrhU0h0dJ++4t2MuOLrCZCjM
UGkknguIK55j6buz9B6dVYR1fflVNX4hN5VO6IR/w8LVC5SKIHFJvaYawb6d
YoYRhzHSmYjjDNDHW6u7sxPxOZ1rzv/qg3bhyAtxi2beJJAtV8bm2q36XHX5
dZCdp45vmgqfh/nmU29y1R50yIffqTPkkNKpteWH4ZZYxII2gEVQTkysxkGE
h9lcAZC1DZ7JqX1dnm8oMoW1skDXVHSW46PK04dZzsk+up9PLI/yBx1Jc0DW
rUVa3o/WMtNuzi13OL24mfEu2eOGVf+0gmxQ6O247CQew26rKtbH2S3z9N8o
pRTsUDDJFYv4hWq4C5KJey715ddGA5h1Nuov6CBL7N4zvfrWDCJfEBsSmAtH
eZ+bz0fNwUFGyXb2BfihWegcUcKSUC0fo2MdSqElEBKts2CqfWcISMUUsqFC
EShEV0ASfoSSYBG/YyI/Z7HATNCnHKbqtPeh4iIddGudFKrxfhGmVIWzBujG
D3t9VPTKrT4Esi+2VustyTHFk2FcfNmP8W+7uqme9oO8jb7YUKExHyKx30ja
iSLpKbxOFH0vQEi0ieE8IGxhBsLnTdp1XULEJJejCn/ay9vxUm6TNg23Xvdq
MCPPjimCCSCPDQl12bxWH81Z1WjaVff0wC6G0Ti8hA3WhGSZGMAPSgpzEyyx
J6vd/dyEIx86ln5MIousAyL8mLb7EFumpnW7/wRTjS4Tu2q1x5UjXcYe6jeT
pn2UHzhha+lNQHT3owbxw4OJMHiIYJM3qlm2SaFLdOYWYxRVQqNRNZyJuiEv
rXRRGT32rv54EoGo6dkRdD8V0rBOVhOBgtLe/RcaTj9KJye5xndWVrk5ldxf
T7XZt7YJz8DIwNZlcjwT864dOLdp7kdXVnOxf05uMBuuBqZBkHH90fFAwvVF
/HpNMKKEVQHC7orYjLxdbiedt0oghQKbOnikKJZ+sIJtrNI2AVBVkpZ1K2SO
RupNJ7PNYz7gfDgwITdW+eSmlbkiD1mSy/sDHuw8Rp6KghOQKSks2pxoEW+Y
+EGildsp756A2HoL+gb85i5K2xrPRKdNH79EaS8cC/ESzjEHj9pbnq9s1ENq
JOtSeOm7QlNC2plC70LBkKVKs2vAlyxfardVFxhPv38wfBPQ+FQxw/d0NSjd
g/smEJDMwrlJtnMe811M5DeDhZfgrpMf8pJqWzwffHBjBfm+Be6gNWnPI17M
Ul9zp+ZQrhryh/NbsInqDoSFLcHIUoKDXj1X5A4bwzX1H44WrZxPEtnsOArM
7i8p1miqpK2THgRFSFvl1lfx/ag7KPrEh+qMbw8HtSo3jVSAEjzZVrNv+3n6
c9k0R22vjyqvua/CXEucj2qMI0VEMxK9ZoUtMOIGJ+6mWv4m7n+dr07cuBZL
Za/NRDjTumfkt2I49NWc6k7q4SKrTISgcqTKPT/zmF2eA0PA0akzL1S7SH22
bvog4E8DJuh5JTg3UtFS5XyP9MNqzgFHANNNH8X6KQ6wydkWRymQx9WOIW9T
Ht+UuHu808le8dd7YkAa5uo7+IA3U6n2+DV0K97CBhxwKcvKtA3Qdj4g/zk9
JlRkUcosV7rjsDWu8S9kz4o9+/CT3OJeS7paS6NDVUot0sYL8VS0fGs4Seev
hqISAfEgiw0Dq8Dv2w1BqCl24kDXpz6Rn+PXuqDNE3wW4QTE4Rx4UUqcEIDQ
q6kmx7m4OrcQ/S4APi+z6kEoftjA7Y16FMSIiTysAM2jqD/PB5HzRNEU2jnr
zsxhzilMiwlcYAmOA+sTwVz/DN3lJLkKZQCtOEkbmtHByA2uoHtuOhYFZnAh
hoprFn9huyjAO2Xxp2eN54mKbdqdR13JLzUCjcTWJWlVDR35WvYl7FlebBSD
85nkxk59ZxJcVzPHMt3b0uN2MnltUmCX3JRPPEYwmgKkKv8eoH2+S8pkzn2H
l6bc90DuVbmtrcKp4yb1q9js7nTqq10JOc5/0g+msOb8A4yKuNof0ko/j7ip
4LRgP6S740Z8Ph7M1ji1OZTKoVkL2S+hpt1p3PQ8YPN2mt+hhQZO3t2dU5Po
Evh4RuN89dM9VXTAVEpsmFbc27gV4a5kNrV05elf60JTRdQJ+EM4Ysmh8fLL
x9tPkmeBGw1yWWl9k8JNgCga4xg3ikrvlAljtNrFQ/8xVYcRjZkGsGbCzNmA
TBAv3KX+DEzYkV+xWo9BgmYzqyWQO97e25LxlKjWBDpHQr5zZU7T2xB0bPSf
3kAh2NgPSuxDbwcDmG9c0fm923zxqh8iQNRruBaTtmDt6fATywzUkPY48K6E
TYu0Kj+3tw8gphp2lsfpXS/aTl7fyuvwgCpIsTDt+iBUFc/wGbe6w0UtR2Qp
HX2GFiZ6nVAfXOABf1ycjIOHRLF6zcz1JCwuDA3cQUYu4dy5rp6D/hIev4KY
wXcS6aAKY6Sm63Kcn25v5mwvtazU5eR6FZrithzbeHJtTxBvvGNkdB49naSV
x4Qm5IgR2WbI8dS2AzCvNmk3gZ8VUabBuBNDtiAzSN9DKiU/Ku0GGHQc4PJ3
K22l0W+7F/PczoqOglVS50UsA6kfMVlh3V4emxKS2O+3BGd65DVRt4VJVMNx
TfbiFcXcQxFyNHh+62VpGngH2uz0jlpOWmEeuoG+atrCk1czocF30p5NwqMr
SLDnPPTZVDxuC+Fv7HhJO7iq+jYnYP94mE4MG6c7b94GcvclGEr99t5OnUTx
if5mzGAQvmb9dGqmqNekHp+e6DaZH67AJFbIZ4S/FXW8kNd6l6i5XjSm+qtK
Cppzx8/vRNW54uXtq9bWADYEiDNYg1y0MgR0o+7wQuZ5wlxCkzwC/aFus+I4
ATopHP/hSq9cHnLcw9RAGBad5hyx4M27Nay404COA7bBHF6/HPBvzNQ+UOWb
jUzdpNQilkwu9l3Sa5+Alc54zY1B+haHRYkGtwnc2rOuotxYQxoBsYZjZvEh
IhNqxLlb9tawbvcOYT2VFvdDWktnE5ka8x9qkIyiivtB+ePJ08gPIDACzhax
RXnI3ZAoXJa8aIrB2ScWHDRTssZ0rEsQZfTB20JROxwrk5a+resP/PCHup69
V0aG/iQvI9IOw6Xp4mUSJHk3aqgeLusySdlUc/c3c/FHQ9pHdEDbLOeaa8Sr
VN/u8eefsr6GBb2DOhs8oEUpFOdpWxxGlbLqq1kNOOJ5N8KXgzjc+Xt10jPm
gScc+qDvlpM8naMnJAXxAGFS9+SOudt73Jr5CGjSbyIbo5CdMUiFBRDLBYKo
3RZMyBPd1KRPUoaUsQ1NDrzqVn5r0gmbo8vpefYOIsmJ3B4dOaMiqTgz3iyw
TAdGbA2+bcR1CDvr83OkVNIoMo3ob1XHQg6A/BI/59LuZ8JOPH2XDLY1GVr+
uEj6t3qJd2HrZA6k2ji2BezUHx+AWR53WM5bXvbJOF0Rj4+ig15O+9dNOOKz
jQlvVD4GIaE/9m71QS8jCBRWZ8nsoAaiXUOnBwGrQ3RC63rSVI5mQS3Hj88e
e3U8ap5J/TVdSTn2jWi7u97lzbZ8nA+QfrvMvzPWL3fIi15HHP7Ds485U8dA
pKA51pzP0GWVXZqaxv7177QVx6Fo7mAQOJotpdhjO/E02PGx/1ISkBK6db5K
YD5+OmS0FU7zuhqlwJof9oWCiW959g+Rjc7fzU0H/HZLw0nFTH9flG4etVq0
nlglnrLPXH+UMgUofQSXOc6+MAkFlMtqltxc2tDihS9mH58eO2bX7aXz+oTq
OO7youKiOmKtWKf9L57QcONqGdzTQ3eKGX+5oSi2TRpV66+b5p1DkwRyq1wZ
XehukkHuEL1kk+BXe2rNeH6cES+QNf3xdehU6eAM6mx6jR6MKa5KmZ13lHiF
ITrJJy7sKejLOfis/JwjvkpYF9rE3esqoYm4YQMJtHU3dagIJQYwVeQt1rYw
qthsYmy8C4dLOZ9SiowE1uOFCvz6xBq5Qy1d1FuHw7UFwbp4dIy063g7DmvU
6/Fj+LhRW0N15EVRxEYUVlhbrYeWFeBHf6IsrXXpq/lqiEs1GffkbVB9XzCd
6kLHB6BUO3O3/J3vFNN8p5jyIfKVXbG/xw8kwtfCN/A2TMi/nsxzubfnKuIW
XBhkmPRZJYw8ZGWjEXtteKLy1vEOwH2IljqzEicnfOWTnEhVze51MrL/fSeo
sxNhcsIMIPTdP4BaKGCblfXevorTwReI9qCWeZzA/TJDtOZ/JNC+pjopYx/F
oTXaoYG9hOjmP7qvz4EweUJ9rKO8M/dPpSC75DSgGF2pf68eipquWas66EZO
mnyHddu+ZYUaYGOtsn/ZkXZeIpvc8M2oFraEvLkde1zVzwZ4XGeZwyZbbfpH
y7mfAmYw+ANllpLQgpVJlSKb031Kg4mbx0dcaHYJLfLX9p31QLSHRkZwqSe4
w3GL8egfvlTYykqIH0BBgjYSbhrDlnbDZO7ao214dZw5r36k+IkYQmhPlyXJ
o8iRwHgao+Z5FZ7yHy3uSOStvYUCkUNCGFPNy+PB17QsxA3zcWDHOqKEqmuu
3bRjUnavqqSuVddfAHmUvWZauTDLWqVie8neegRJqSqzn64uyTDIHauZtnCv
mtj+3apOA7UhIPjWnD/kSlR2fLubnXwTBilHzrc0og47KCq9C6ucdjK7o5As
qJhiiNw8LNdAoBaL7tXbDPo7QCIfXUzXWzoiWT39yBNmrJbbrcyTwQsQHtTd
G6o0rBtb8fYXQLsk0r1x8FB5Y3UCRO2deXz11gHtdu1sPj2IxgrDPnSJx9cA
qyqB2rOdGE0zY0IxYGiKjun84WacT+Mr8H/Zz15dcBwSjowqKDRJiPEMrQCc
b8JEMXMED/OsjY1nE8hb2Gdvfm4BlvRQLpzRgYYrMbWhmhZlc+o3bPUcuUVl
RtfW6R6lo9N173c7a8STzvlI3wC2Qs8LShSs4jQMSUN6b5c+nERNpe70JS5d
8BLlaMUyK3wPtC+XD3JGaivo9JMcpHOyKHUiWb4H3Zw6cQfai/0MnsuH6hv1
8wz1b5UAv7WBxe0sDnS3lg6CsE+0vQWdxXfdKhddnjY1a/OLRYyIZgDpEJd3
Zxmtqjl5du1KXcQAeY6MQ6s8FM2d1HQKFfvb4EXelcyhLc5cBY775mBmNhmG
oX0w20w9rA7PiAK43tn/AYvq9JM6rvAsMpGHSkeVIgiNTIMu4GGsMd+6kjcG
dfKJqHrPlhH2Dz620Wy0xo4u2eS+YhUgq/gEtKf6wcwtKK26PP/5oXBIqVYw
cT2DlfW1blsUaUOAJH2d8wELD4wd1COnPa+JXq6AtMECGfZxjAdGPp+lASvn
NHUPt59AhqsBxfyEtIbuHvRpUjQ4h+H4+nCmC+v1Zj3mMGk3Wq2dYc3oheUG
oJoSDHsmAX0KJN/BjeUWVNVycxUnPb2Y2pax+b7t3NO7vBkFkuZFON6j10kn
IDiviqQq7+E2DfQpah0NO6MIykimzFjWgVTvuLUhXbarqai/P/wBdNPzCQfT
pcQksqn+6Dksvc8e5dImbaEgvJqdirVtnZUku1vqvk6ARQz9haCdKDgPsWLY
JW/IwrD9rU801xkXKM4q8RtneVkx8C00Mlk2zIh25wunb3N0kRHz9ouFgpfZ
UJcILrk+y+5mztbLO1c+lnWty+3qPWOsj8+nWWVDZuYRB/weI7K24b6j8IOH
Vp2Wn/IAD8xPrkTyYCqERAq42vz5kXEY1gkt29tIvf3U/5kRwnpbsiV+aiMe
ArmBtVaFGsC04dxnHO3HwYC7QvWmK1b7LgWYuPgA8xeE6Q26fX6klIdLRtL2
Hno/c/WdY4YZ/FFqce/v2dVCnL0Wi8Ic0E9w+KtVfo4uCcQZkQAYpQxuheyn
/XSLqSZF5k7/2Y4WTUkwSfL8NOkXnSwA5hw6pCHQWbl2MfjtviJESl2xdwD5
cKUXioD1BwZP4z2n0cjw43aX8Iqj+KpVTk+GAX7+q55uFQFXd9C5mNEdson2
JuVcMWhsevXmtpUXxLHl/4gFAWAXOcxUYRNNxj5HV9W8vsBHDy3kOLjjnrsz
I05/4OUGbgeFRa0qMCraOZOhoW2m8dVNJGIWs36E7fIr2dsqPYENw0SNjIyD
38glAg+xIhHheAG8n5xxgQL3nHHFrTU+aT/1IjS9hSuiQngjomB/algKVf6F
Vsx3TSG0d4ZUmZwG25U+v43saWrDCcBXSfhjbq+HXK60ePsWLzmDAwfH5t8l
2RJ8Pw2RHj18t51BLasOiGr7raq92/aDkWHc5PY9+2R+JX8yeHr4XZP9zwFI
oqkzUBCCmhJMKVoMO1/BzY/TbgGcQxMpnVyXNc8yrHRjkW9Xed3apxiOv/+s
dVHZzUDPxsGyeamMo80GsnVviRBtVM05nN79iCgJTCXbtEq8IHyLC0EMop7z
9kS+zyfLb28utYWKh82HqlrTMC6vFQR4Xzae8f1iC7lDDm2NJYn2j72O26U6
1LS3EMu2tjUZYmMSN7tzcES0wmsURump4naKQnSXMTpK6tYH4TdwshH84i+v
SXoe0OHfQi8fQqlhueP2s+r6Ah5ETICVCnHVv4s1FmJU2ALmOPP9SWy5oecA
Ns1Qq2MTpRRaal7wp6zw96KppwLp3pNc5nH+9x1a3jkhoJZztnVush01cOLf
uyoJJ0Z+fpKHhqGcRVdEk+brAj1v+dtVgVvSYsXdrf4fwXFqJBZ8dtdbNtmo
bY9+92zs9WfPIVsOALvYfi2RORxoXFTqzJ89FC1bIVGMf3BC4O1tMqCPlROv
VCtz7pdZ+CHvFxXBo05YY7UO7i61h0TWq1G7jQM9qSKeOVLIzeUrdOiXnQqz
SJBMinjzPVDTOoZraIip5t3LXaIQf/zDYFiWb3fwX6cSWiK6yhZrV+kzS0iX
zCj9P41aCXP16eUVfqPC6/srYO2QgDhGH6bkSi2BJWUGiXpvR96wsb5+uXVG
ZP9oqY9v4M6c8fm9fj6Me1hwEMQD2DrGSUbacsHVoP3BEwE3900VqD/GCWYC
o+yRn4WB4Q/TSW4DIcWP94/gR9bkpeNKWEWbkCjqUCe6CR/sL/N3l+06tlKJ
uam23AIGG7CIBLjq1OtBiG5i9UhxCYYaDZM/zlQMZ9HrRmzL9O11z6TIxMov
Ntf6msq9/BjxXcqKIBDX9YiVqFhBas+tI4OOSffFpdgB1hdUFbX06a+cqor5
NoBCGEQJJOXO9X5tu0qNvZvINqH+1xEHHxLRbf8hDB+TdFm4dzkEDsghqu3q
oW60qaXABhZS98PJH0d3E4Y83CRZR7CoCz/cs6ptcu97XU4GUUAoZae0itVH
1cXKFtTsBSAQ6rZt3lw4ssb2Uwe/f7m8XiWweqPpI4SE1R9HoDnRaSDvL2ux
Ugj/VJimQ0yWWjyuKY0CDXCE/CxgD8htnkGr76NAAMFF4JsfoMM4yDFyu/PM
Enhpdl9SYbGuGquItuVT/PtqFK4lM0guOqc4kn2KD1NkgIDPXi5m2FMMhZGt
DGbJXWiUk0YAd3jwxswKIkuhFffwl2DgIk1ybohqwidXWzoo/zeFKbT5m79M
ZWCDMOvM+I2xOFZGak4C7bnrcAhOxYto0fD5wSwSFnd1tcjCb/Vy7mYUTQcC
taH57tQLJ1cNUqbEopJYCgw9Qeq/fnBQ9uDXZhkI7LkSuuLL6rKC9facwEFu
TWEe2Y9ctEFVq2PVHmK/wqvMZQNcGvwfyfr2mSlqFto6ejJoYPvVzwQNYCO9
sa0iqBxb/SyPxqzywhicInQnm33Z4WK+W9CgCqSU9Cl2d/m2D4YdU8skumBt
Dv13V2sildpqVVXoX1yE9ppQ+rueHWFjAWKon4l/izfO1HyN7KiUreCE/APM
z3/dAGQtN9RL7FDaHIiFqMumvqJ98SATWFSHVMofRjGG6dL9ORCsQEw4SnxX
OqYPac6gAdce44QV02Glbvgswfvx0b6Pz/2jpRn+xkWV+fFTQVJ8LHgRP0q6
4MR+aLjHZlpY3JQOGn2zyYCODpxxYZaORyI7KoaslcXtUxHtuOs+M0q5d9i3
0tHy0idmWqVhzaON9/RSrnXTqSFvNQ2UEv/aUS+dtLhtovwyEZIyoI8+/lcx
ZCG6OeIo+O6T7nyirLX/KEFiOeVU7WryMq2KlCwBqidvylF+VjO3h6leu0hE
johDoSjU2YXfbmn4SsaDz7qyLP3LUKGZNBF6yfRz2Wv5Vfkz9CScMa5ssE0u
JWYHgXDSXKKjCVFJvcAlr+AtKrsRYXaeW5KajN4zEhLduKBkBJ4fBJRuy//P
muFhAirhOhkiCX7wqj+V3F6sL5/oTL8ct/ImdeMV3Wg7b+EWHMYVkb5ihJHd
uyA1Z15Dhg8MUDnIpIldyYB0O2B+8Y6uquWKh1EdFZe27c9w05Ldbxwdslvu
N41zKPdc0pqK1bbBrU3JyCxdo4sRNaqip7CISuSZDEKDAc4K3Ck27CXw/Yli
2AwzblF8PyrPLob8ws/UoMDFKmDAPS4PUhVt0DVRDcimX26++kjdlHYY4ixC
VUKMg7SW/F6Tn1iPw2xYQgms/Ht3ZsAlu+5QPP470gpIolzlSCfaIHeOhhok
RPt0+7V4uP908lgsNkjz9kpwo9/WmG8+KeBw69661LYGiXRR1mrWyV7VXKti
IU/7rMchpZ9DkYfZbt48+dRfFxEYqyhF+DcA1dcOClxEm/h4r1A92C3g2G3o
CXCLSpi/Za3uUd3TP1deEzmEl25qEsJSvj2+jNpXQqvFn3SElOz9cUIBGMCt
NNhMjIRrlquhnldszUTPrU9bsYBu20JkfyXyXgxVvXbMCcT3n7mnCTn16bQF
2c1BXVPYcdqFoynz+KSHTg/Qr51XAI4ChieUPwiI7UsDtlP7qqsRxGHF6OXB
x8BM+2oYufq3usI0tJSDSaRQ/ufKIo6ra7lyXY5uzK4kQz6Nc3e0bq//Xq/w
GxeAJOHMZRVG02mtxVsVi9CUMZsYMKS/SHNWqN2ery/k1bgoSQalp75DUwLS
wg2wmw/dnAxOK8iFvtJobs+Z2T78LXVEb6n1UrpFJrsmqsOEw2oTRD3bP5Pf
Ux08C2SI+/kFw9dSotkWfKp39sJssRgipX5BIURr4gwLJqyRnWXl+2RGKK9J
Cvs+0wT39sNphaGceH9sfC4lyRJwVpcL7W9sufZJx/jmQgwkND/0wLjFgkVv
OGVzwx0ya327NMT5onXT1rzgnVdOY43XU6CfGTl69Gv15leVA3Zj/gLrXytm
PiCoNIUBcun1gkB5MNHPltcvcCWG4dz5o/mzwXJZ4jxVPi91yulM7WoxbrSs
XHXHKV8PF/006hrAnaYIR+IxcgFYqQiMhAeMWJsXUPaB9+O0t2TBR7hX9ER4
KG1O/5mEVCm4QXxg8DvMU6hvPo5HW0OaqJ3DMCr64AP2abkS5dkNRXWTcOO/
TpV93ljIvhelq34Ow6psWkvSBrtDmBjAGyWyVWffKTl9oFCaR0eLkzeNZVCG
liyTObj4Nq/yjFdm+OKyG+w1l5TYqW+unNHLmRROHih6JGVWpZu1W5u58sDV
FZC9+wBU2pLaa2eDiM+jVVbLVVyM7AmuQWa4YlspIkQfHwE2sKx1iqHkNRbJ
y0L1H1wJSdref8nZp+zTu2t5bASP8EQEHXeC9pTP5ssEB1WEBFvU/XvPRnzB
VWtSjXm4r0RHWQdxWMfUknaKP4qJPOV95HvvDC5+FshbSqL8D7EnIYIuLNSo
+je3WOrI7zHQtzIgy4HBoMDRC6gAhtPG6VYGVnkmzXJQZq1uTDuVroktyL5K
SjhEoQJ58GtTVHpmBNgWNr6O17tEfX6XMdQ+wtJ6AEX8db4EG29K6sgLT4Dt
qQR1IjnV15H+bgnpjOapMrWHp5Xm/n6Am57zQqDkbgDqfrNV27xCJUIUSuuw
vHxIopC0wP/7CG6AuXor0zgvf7t3NWqX+xYqyrNzdwtXerogdI/3fgXUpoq+
upypDwsTfLFtAojE33o2Xehg9JvIeqz+hstXs6TUE3J8JeoKSh+s8xBbEzow
hEuekYPf0YnVWsEcp3/0JZ4F2SgvZvCh4cH+/MQEZKtL7DQAhvcmQX7R+Ntn
dMT2fXm0fYA110Qitekqx2TLYXDl197Zp4MLkSbfrsJsrYQUb98kn53q+rds
r/lum3EuEzfORTeHw6kPZmnLE129fORJu/cYSdyTzbbLCxOFWd39rN2U/tFF
YjL9c5gt8BdqyARUK2rBiFBojDnkQB21ybYwO7bo+CxgNRSS5aRvSOUwuRUt
3+yhNBDH6orMVUloVOMES4f4owvLW05qcBBG4NV1ZIRuY/tW3rdYWpW5Xz7c
/78lyR1JxP2cEl7sHsOBgitxZlH9mMu1WPwmFKsAdmbciXUn13UjfbhDFeae
L4xchk/u1ebYKZl5bsSlNtEn8XMnICDM3G4iz7KEPVCTxjYpu+3BueXAjI/u
SMrka9Zl5QpzAA51QcC85gc9pWMlx5/8+E0qEzN+k5Ntmgw2f7Gw7RVXB9+o
FCUINABZuKy9h9tprk2HnK6Dtg58vSl0Nt0h9paAGZvfpatnCpw9mmgHEUV+
YMcDQdfMCRXFA63EVDaHMGF4DS3zJiH/3fDKdrSiW4PoiS7PWDZ6stoKFMUn
YZ83PJo3nfPhC9j34lqIe8Orn6DbJYBFx78mmGx8P7ncu6k4HjFtGW/8B5AC
fuolwxYPTQZo1I1t4gi71va5GZ/PXxyPLL5UVxz2GJvQf/ZvOgTa7o1i8TC9
crN2R4ZreUt4haPhHNs0olm9L/OJlp27S5C5q4yiMIkoWEQQLu+S3waj9e/b
I0LQQnSjUyU07K0OzK219zIosM1PMNZ5t78eJQfnPMEBg+ShjEVP5At0w7Uo
IcbTivw72bzG4x63/Vjd3lSYT6NZGvmCbjtikwCkouNqU4JPIF3n4GtGJVBX
KBqoPDamvBIkXBpPajLBKhDL2Kj6Gh0moFFJ9NZdJ6suWJAy2tFWOkr8qmtV
q9AQX75wd9D+c1ou40GstAAUEiNcJddkC5HAfPueFhq8bolgyAiiBQSE8xtS
+o1x76E1VZFc7Nl8aiCt7rG55km5L3u2f+rXXAVaKkmBnwvLf+d8pzqrJRfr
MqWdpLgfCO2EYGATtCLTD3OZKXlzzYZPiC9T6cZGaZzesLdvFnih9w+x2IXt
pUMZT6nODNKSxtFmFIXT2gDoPfwhTvgnTyxLXRKLeJuaufYm9pq20Eymsjq9
3Hobtw+f2tCa6iy9jA/PRGrGO74/JWC73PmubXiDJEJBb/HWYXl0dagF1Jbm
JXzyU1D7LtfV4pl/i+15oKCK83Rb8BZsjV6DKW9tLoiQIPjDu9if+MwAN0M/
fq8MU/Ykng7reGyLjKtvJWyu/j/GgCaUQaNwmqzBiPJ3y6IcvcAVp7UMJqHg
nmpqbQO4Mfa5GFMwgGTRE0CCK6vLhYs/3+b092oS1x6IAzTzS/aD1IsZ1iGm
Pfohj0CBRXBFUeb1QmTpr+tkZXQFMTQN5QDoJ1sUQPiljEQPngiQMLPOefAf
Ergia86is7IBE5aq5M89cmrIikfxwVQElwkHThymG4G6w3H4agasFDMnAODe
GmW6DWGl+OKp8Yp9SWsWlFAgpXtPodpSngQmhFUOR1aFrYwTRaFkmXAXo1SM
JXTT2UvwFNxJpMZr16NLF/ZY/AGXYv5Z8QKN2tSRLdAyuaBnIUXe/JpKykjB
cqwkBJNTDs5410b0QIUWucxpO0hYZV3wajuzq5ryGulTBvYHoJBhLPPmaXZC
7G0R7UE4VrOxHni4xSiWJ5fCSq8SaYB8gvbYOHO1yCyPVsaVimmx5I9XVshB
oMqOF0sHAkuD4xgDFpeZaue285lCbE5H2z6AurlFEyFcvMcfOhrcxo5Ve3Qw
fyW97fBDgl466gBd1fE1Nq06gN4PvbTVH7KcDcFemwitWTmXEaDAJxbRE67f
i+a8gNbsMMXmI7zaXWqkN22toXQPU9ys9xIW9s5G4EYDjhPjbbZeQHgFdxCV
v87IkHkPC3f+wCJfVtcPIzmKc4LItl+WbjOfUbiZI/35iDwLNyoIk67qnwOo
xJsg8zmmtLACBVGdScW5E703T1GN6o1UPZmNA3wLpIa8prbZgs0Wzt6gEofh
HtcNrc9NW0wtTe8ZQVvOE5OcK7Fs3tp8DOU65kriDmlWw57cpTsTEOUwZ2xs
Xoz6qQ/cjE98qiF/6jac3ojYTIQ5lmhOcWw8BQ8gnRguiaQqYifZ1M4HfxOr
5WXXbW79RQYq8GkUZ9PtuE6bvMNHt0DsCdo6AIvEcPXoj9pMrLhZLElMkdE7
c3XLSFr8HWsUvfw3hjCXkNAD9BHHXZhVB0yrKBwymX7gUzDOezzPI+7LBO+F
zlmXVlwB4TUlqFY5gUdiFeHko20kEPyMgHlZ0Rzb6jIn/QiWjevnWeDBdf79
sT1C9Fp85epcrR+s6rmAP1KvWzmpcOx3BCx68ugFM3rKcr2gXjbVssFjHF2P
x6QiXnXftCXxtGY6uXF+Z2ZV5STOWCGWliAuRJK6GZk7FfcHRRZUVv932CVw
EYlRxApoKzZQa95DkQb3j6I58iHKfzYp1ATOiM0Hc9hSZjyOVKsGPJot3uUA
dOBO9f5Wn7RAN1sRHvoYhI79G6V0c50NpqyXemSCMEf7lwPYAzuJMBqWhxGy
bHo4ndgllFYA8agF6+fepbEOXGABxLOKxo3Y99bSYLkH/efL8cDyaEcPaGjS
MDnfpevMJvQ0+JetBsa+DPd/obqlzIKwBXPcwN+6Tk7GsEQ1fAn9rj8c7e7I
EAWsAZzU10xWEUS8VFng8LaOrHGkZtyU541XbrXze8dwagBsCuAP5dr5JPxb
zPjSp4ThqCPaUtinQ5tuVhd0Wwg2EzxFK7wE+8ZVzHqiTni0opMxKg8VVXHa
PkZl1cGnEpIgoQH6RrNBWYJpUPcHt6JDpCe/GsfjgeUjrN8UchpZQQIbRwkn
8qhyffBL/LdTL17uCyq4CDGaWW8xzc2+sUdB88iFraF7MutsoklQG42aQk1h
0ZTUPzIQKQTDh3La8VkKuXmx7XDeNT8pnqv5dP50Y1t3lUJBtIjy4jRQ64C1
W9A3/e/p1QqXBkrCcQL845rD2OG3rzmnVH1Wdz3oNAmUTZ9BJV3XMYFnW3Az
W2uE11jqvOGp+IhWp0sXsNAYG64EAsMPe/dovyyjXCMzvtC7zWClmlguarSb
PhkAVOwkM7Agzv7nsKXMlgoIYaFK730yvpAepPKCdPw1JMHX2h6MdrnEOWev
nquG8ORyzA2eOo42MaqQouOa90wkD3pql4QjfOvZLp1Z7bSat2At0RgR2/kX
LuBYuKok9jwdaCkl3YhIo/1cjz6XuuR/DVLvstu6r0QeJcO1bmV6SICUD4Hm
e3kgj0gfsS7d85HJ9l/9VgOnis70s/J/IvYoRS+gnF/UL0zYUZH+KRUCdOGS
24+2LZNNJlPDu2VjnHMqH2+NSORxBJ9EzgMbSIY56Fun3IUdQOkRdYof68GV
7BeMF2cRrlpqz0liOcIl2Cgpfvc5O88EJWChiaVuuRNTAyKSTYHktj6er0d0
RIeB2Hra+7ilGTsmZz0CQQPWv/sGCubdGwUf3v3Q/upBNVo4s/0dR9T2wETi
p90lm4EnSHbXwzAwLdr7YNUKjwWM9fAU9WqnFy9qiIMGaruKaWSv2XfnKE2M
LaShcnEplPHL+3eA3iwEK6aFzybmcw/99Eq3QYpThNUhZUnjBWF4taryA2Xc
0LzYim9CLULGrmru0XoZsJI6tQtO0w6OByhBmNjoHhhT9Fduet2GoNa1idQ7
e7871P2EP3hklEpY2oYIObgZIYui+Gc+ne63rDD3+RjjvBK0IBC7Y7hWI7sT
PLra1MIk2WGL02v0kREm/12wShA62Lxtoe+rID1JYULM2ydmVkub5ZDQT3oh
7ntba+tUBxetYKfqbkCeTVFKuFj37GdpeSFysfGA0ktz7H2w//gTFegLp8Uw
Yd06qhyTrfCUpx8L3wxdiAH78KzrX3atA0Qy+EClrk3RjntjwrJrK1nUrF3w
7XmMWVL3AVSxUnfvFVBqKKhchuCehsHqgP/NYhNJZWlG3hl0ENGUPgCaCNC4
T4ISI2ierpk3BWIgaH7Okk5yC+k4XdgfRXLOxd/ok3+zefKk8oyqIY73zw5b
boKlMhbZZ2HWPRYH1JL1lJOLHs9F6PS4S5REUxwszl5xvnfp/NkbV71ysG2s
ZNBqMOssJWM/YSBAIwazzjhA5qSB0bX5cc3aG3tpMGqI0msa0WC1Fp+pc6Mb
o2GVKwwGxDTsQZkNDDOCfHnGoRefynSRNJRVUxa39OYf7+27y95i0Pjx6gyb
IpOyJN8WEOniuDSKHQRPLaNCQvbchX1ZXjYoJIXokuq6UK3wjc9WSs6pLS2E
yEWp6qXCaBC/h8trhpXN7etGtepTA5xwJ5a+LGXuPh5oPW7fC2VtDht/PFf3
3PXAGEVUnEJS3UkrkTSndqh/gzk+jA4lThYplXJ230+2WLyXC/kjHiP6bvTo
+YtyAeVD4LIWpjH3FNoiJFPoVxcA/1GgaZd1FVvl/p9vBvxd8b/y2yLtOxyb
ImL76UW8OzFMV0az24YK3bMChL7wb7ND/RdSYrp7bMjactTmHjIuztVbWuez
IXEb7xdXwlEestLh1qQSD+4jIQFPQ5T6oy4d4GcM6QNwpsNJQDX8ve5enjG0
Vl5LweWPEa6Lm9596h2ecrYgIA5QAfYfOsHSdwHh1EAm3DJyIR76bP3AAgzz
LmrQod/KVjXzWUWsGNtWlbwMXueAqQrkpRtN5Cp22JayurR0dgWfCllVg4nm
XxD4HB+3lkVuparvmTeds9aLT/ow77f/Y/iF/8CnsmNdFyudbd+QBFz6Shpv
5oUH7wmEeU+BWmYuSRc2f61YWlVqmd5LkdRC2+vD4+0WhxQfIzBbjXS6ArTZ
ZsfQ7SAFvgB8OVfM6Y/+BvKZc38FaBMkHKsl4h23hQHkpw0evIQQu30W0vQh
u1HDaTX7R96TMbDYekY0BEocogrNe7iJ3xLobzTYPdiKCfnm8hdNFY8ciA3H
iCJxXijJHxPFyhNWxzLe8VfsYCaqaVE6X2nKWI9id0C/82cRtHfC86F/SwPN
b+A5b67TeBRpBUI5t3pPdkXaRrtG5Qjs5o2aiQpc0Nqk8otUaf8Ra2TdH6ZC
XI+B9c0dvOFB06OBRU4n3/6xmrbTmAdDZ7B3R6ce1d+COKK1fAlk6ekpXj7w
Rao2qXPpOVUBCOYB61KNSKeieHrWXGdtFip4WjevEO1ehSlchMwK1rnMl+RZ
1948FdgtkAgbDYxCdouWBmIOWHl0yb4Bc+NK6eTGz3YJT1+CY6zru2AF6/vl
YliS4vJaxzMn8v83+694g9EK7NCYpuNiUZUnoD97n2A73C+X6CuOcfgj5Rcq
z5sd9Cwp471xpYLOAyBhPxKmE/FmVKhSo7/rZ0TCbgynd4f5vwxc2Ou4wa3Y
9yEZxOjy2uOQZahbabFQlPmngMDk1WH7a04jI4n/DcilBNO3saF7tE89P8Pw
uM6Bt0V+t2LjCBkUyhd2/jcIRRGfS4oK0IyeEwmCGTgbopIAjJHMWTpqQgDp
dg498TY0tj73JXWEy/7z2lQL5c/7VNYUVTsrW9jrw3qejKB5wrzvlAZB0+hX
Fj05QyPFYNnqqWCWez5bYGADo3D4uQW4jdd5ndUKXCf4oHlUOJqIR4KgJmaP
38pT9hDtVPncrrEYuTPMFfL3Wa/U1SQ+iRpjqzluCuoHAlBeA53LMqqZtxh0
I22lj17Zvgye7y0tzY8ucJj7h11iyhUqgvpWQDsW9/XpWwzGxsUN0VrHp1kG
XCKDLYl1mJj1u/keASsxm/5XDHvExngfmhkx1vglwri9PTkZu2RNuoc0gXeJ
bLEgOvtLvJbvVLxGEGGBgTYM+YsJvbD658yCUsKRssa60xVtFwbfLlVTCmlA
7n9HFaPDwSRvAAcaC0KC295hzzEDr5nsJ3tLMFxG+eTDL0NEr/6DSXziowbx
jImr3wzVdFIrbP+qwTFPpqJHrJ+U9VO5l1rrDrOri497XqEf+bMHfs2AthM6
jmFNZ5s+/ZAQxI506V8DskunN9VIwKjwRgHPwmPYf7ZY/KnYRv0WA/I0t0jj
VG+pF5ubdrStWNogBt63CwSwgYQm5Orgo36DGBr2pU6bq0/0wQzmhYKXVEhP
2ukh81LK+V7PhKvoq7L9K7Zmxff2CuhXbzrxORZy+neIJ995y0H6nJxWW5Dm
vnXL31XXD2BZ56KOl0NseFrc6hCOzEbQ8MIXXhODmIgqz6p/88bC/Q/z5WFX
RfzqO8Z+wmStM4FEWl9OOpB2PkNvBHRuOBxA8TUHDSO+I44pZx7k4UXb5dYG
ZAogm+igdpkiisFK6FY2V98oS7gJ7Gt8op2BDI25iqJnxxII0t4vYJFACRAM
Y2DSdZaYYl9RkWTX8RW9iyFxmQHVNakF8Z5Wap2fnTFxC3yVELefL0J2YP9G
6vKiN3zhlpflqwkvOKIOGAHq4m/swOl2CTv0SQk4b9LvV9K3M3CYbA1en52L
KtoTi/Nz9C8Jlme0xagAG/KSD+Dysphxjmd+W38ZCf4n5sGQS/c66WR2Dg3x
aDCU+OYx7BDeI5xpiD4W0bd8S0vW8LRsnsvnEswwt3l3NJJ9m/gGv8A0v+kq
01b2w6tZoQba0HVVeACl+Pn0tqCK+7sS8EXBCR3oV7liD79yy6/MJo8QAIVa
sI3OIU1f/dltWUvMN47RTNhibxfA2bODqW/+IhlHCMJ4QnZcI5xs8XI0/Lrl
HXhDFLOv4YOIzVbZBSmzcsVIy8Xh8Y428k5+QcF+U9gogCH3j5rCd5DuWrD2
NGGJrQ82Ml7xwLcLkblc7b1Pyoi3Nu4XeGR1QIXHD/2nkBzc1OKz5Yn2k45t
ZZK4HR8uVPaJEa0unVGxxTj5F9uZpPup/2/YSwa2hq0QSVOOunU4Zgp6lzFy
IEDEDbAfFO0dFJPp6h4dxt9jgCgEKLn3qbIHcG4RhOAVuKIBS+Fr0/LhWiSE
GUMmZDhwkYEe2wYuV4Qkmt9S46dlYDHchJwJjoLHZAIpe+STgbJsg1TGUYWn
bGkH8IXb2vfTP17o6npkczOKc9oasU3X7Fnrx/XL5b/oTpvJejE9XuXy6LqB
Qtf62WSZb9GeidvkFDpbH913Zx8tiWkfH6MvJqhB+aNrDb+X1ZsPu8QMP7F6
dK/OpsU7IElCmLTQTbWNs4a1IOpMc3cxAMEJSE/E/6yp3ZZSjCbAPnOcjCAB
pVaG8VPg22uQa1Hraikbg2tg8I9xs13jC0nf5X1fM2Drw7CKHm8e52WJ3G7r
vMDAtPgRmWiK6GAPgu1tui1FTmwElodEpu4zKjraE4VkN9NZ+pVaDw/W1m2k
0E45L4PoY85d3vXwetjF7hu3KacB7wuBrIMet5+7fagHzbQENVUqYPr88iZE
S0j9DIYvKDiVjxzzrouCWSAB0D6npUi3i+f7AdQdh0i+ojBXj1YX/+ieIaEc
sRYoVlpqcNp3AsXi4s7931btirQhU/pSSwRAH+2ej3RPy8Ciy7QWUL7057Va
aGvgmYMv/ZKt9QPFxSusiuGAFE4i9oh6KUC4DSoRwbtx6MaY72GsFmyP+GtG
ialbO3Evx8oszdV2d2gQx9CCx77gi/P30jXM4AszF3PiDXZ/VZYafmX9TIeu
drcAZT/EipusIfI1IPrcN2yHbweVFoR/Kqvqdr7sSowpJ7hY1S2DTF7Pfti3
2+aI43vf6VmsHGJzcYLAyqAjtMwMVluDeaFZsGLLpicOs5Vu6j+7qCvDF3Ty
75qVqohHeGet6rr5l1KHOw274bWshVelSiLgabgU4XbN3yFZeq4n4kO0lSvW
KHsDSZXGoBddB+t8yT4X64S2hrSWRgy03cZVggMSl1lcmzRAqYkeAt4rvo2Q
71lYVIphxWEdn6/9uYJapKqhc3U3doddhD1qvx7eJvodMMobMEFT9Bn2gXKL
dNypIg1YYIRVr/l5BV17Dz4ZUGBR71hlCf2RjMfLV6hzvQhlw93fz4le0tDr
H3VNsBrfKPgR4CiAlNQ6LrFMRNvyNnN2a4NReNEWOBZttl6v3Fh8WIz9JpEQ
yRGyN+0wIREhgNIim6c7wCS8ampxPeYD3HfVxTQZbOXaJs+K/0oxqyORW2V7
2Yqswczb6dl5Xdk5ctOUOv1bjgjsXlqSgaRy4IHZU2YTaI3uAcnxXoOBz54z
m13JjomZYMdKylOFJkSazldqKqreT1Y+5TS4MSOFrngrSM6f7Fk4HqVE+gcQ
YJMaYqLTaPr4PYFSuxOrJBK2/K2SMfOo0m/GJT8fLoLNrhlny7u6lb/mgtsQ
blh2cIXn5bKc/DopeIToU23pyxK4cirWjGtP2JtF8UYrPlNGJv1aSKOABJwD
QZQoOQc1vsh6g4VyMyo8q+LK7A68+SpKofmkSUM3WHDoeSRQRIASOuAX4AJh
UbbhSQCUEpLwNuoUX9kK9ZpOXrgYIOb5au7EpI0S0GWEVjm78zuqy3Vj6zjp
+/kyQ9/acnsFSFLip2SAH0oJwplde4QocTBZu1JqX0MGlY1Qf/yGurSuFdsd
kB2l6gNh/lHBZrU7E3hzbke1IcpRiMZ06Q9Zv6j6eUL14WHNbP+B2nmWGQTE
dVXN2bDbJIOB1bl3SadziD2tUX7O/ecNQQ7samxw6hgvbYSgz3aLDiGcclkx
cu4x9z6Ta/DdxONTyGwnZXffmk4bsIsh+t77ne0jxmJaS9TJ4Wt2MwXIzCz8
q59VMZVgkRbgm5O/yFRJRwe2tH5UA/dTKdf5uCiCLtWPk1zXgvRq4ar8mu0o
q+WTEih3TPSNQLfw49jzF+wv5OCrmEqNVsEuXKJtfdF8pkT2qxSOlfDqnnkU
wX7Gq9OrkbD/9qyEVwWQ2PrNDbgDNulzg5WhjJWjlnOlMLdPn7obRb6B0FDe
FDfHZ0GgCNpu7zJsZhQYz61J0mddtaYOO6HIGW3jDLZplhsukhH5HEUkPlRA
KA/NrQ/MfQsGTcTHVdlbg3Qj1scXHf0rwA+oImACW6eLDMtKlj0CEvHEG+6c
KvoUbmK4wKGHJJztEX7i64yNxnNXxeGeuSVO/xG0RF+jERrpCI2+PRbMnJWO
7QunXwIQeRkyOT8POKWdM5udpjEUric4SaodHXgaWG9J3jxODRhNUA7iigQH
Z4Ou2FCJdpO0oscGfu17Z2MYjyX+RicjSK/wptRhF2vFTYi20+ucSp2J9MRL
iByrYsV/KzVcrFerCA3XT673OTfFaYN0fex7NBdNeU3cKMna56gyoDN0gOkP
AAYD4gZbwFbyTtJMAZzc6aTaKpsDwXyqA2dvNJzPrukpN6aLyInfc6CszwOi
5g/gPvHoxjSq8KuSvwZ5iR8zMaVjd7LgcKOX3cvqJEF6aK4S9ovF6D2/Igsh
7N+cocL4m6jNWzkVouvRafCTO6L+PTBF2qgKbAuXGlz2z3kvuzxU+GrBF3Ws
p1e6NUAN1xyVlQXFUBQUTsNMZynFCeeo9sz/p6kX4/aWX67+S6tTgt827BWY
vQYg7+WuBxz8mjNQxgFFq/bUfz16+KIc8V5Tc3WIggecF9ZADYq/1wm4o3Py
7In1ny6IOn0zKwLh1PVQBVmFjvTPZDKCN6sK0cF8QaNkfva41s+Pmmk5akqY
cHX/0Hz619oENFsbCXTz8SHmWuhOJgC8S4q2XmJg7p64YSifjTEIeggbdcsM
tUCoUvv/O7fbApxDYgYuCd9GzL8gXSd6OnhFLkJPYtnbJhppSrVtJm6hnNbw
bvDI8JBjcDVzZpm/e+hXaexnBQJKqEvqhm0j4FzuRYjWXVIRjvmrkyHPqQt+
/xxTrRElaXmO/LnOfQ63hP4mGDBQh9mtvZee2nO4jWq/+7wrmk82BfFPwnJW
UxZ0B7e6sIUabpg50NHA3yqDi0dOm8wDQw6DSNr9s5kfwrgrQpl3sMK4InFi
pMrdsdgKUaI12LSpGCOOGjsNoCirGzXuoZ1MoMisFLP2WWYEAZrUA0P2ctG+
yZqlEhyQ2arQ3wzhvTXj1t4ygeqc6wwtKYNbm7DAzFiATlPCYFJFPvsyCy/5
xWt7IhOswa8M7yx2vlfbOrh2fsRul46o2GGq5YtKp5RIzlbp1aPGPx6XJqgr
UJ1yh6jlTBD0YZFS5oJKZwI+8MTVKFxVUlfHR07IVWniqU2Jt3BItZWv2V88
wenPNmwPl2IfciaQS0YKhdO8QtwrozhjAF3Lu64KeoeXPOMp4R5yyP82Y4O+
FVW/+iYXDcRvdLKnBU1e1ltXFRhd3hMkMT0MFKGzXkYMZxVZNiSQZG9lFdy3
Yi8usceVttIr+gyLTx6afro3M6K585+aMsSR4kxo5PvQC4kmtC5XonJqS7Fb
Obh0GVk9nkX5QSpevvx/mX9zdgf0UkT+MTC5A3VHbVvxxHEgwjipHO/zEjm+
0v4hLpB69lkI6GT38FYU51q+ecuWs1PqX+DOMsFR3MC7msVA+V637NhPP/aQ
NLztQgbHklAJXe0r1wg24CbNu/Q5GCpbwkVhPaHzqG7ZQYbgIw0Nc9ceK7gb
Cou2bPmva+1t3JBvZlLZ4+5x0X3nlO8nUaj00+2djRbHJsuWEc2l9aV+DkR2
/BGXWpHN3o4XkkM5pNa4kYtViUaPOhcZpEQ7DSHrONE+SLb1zzZPO0qPQ3Pi
Of2dq0aDnJDzcJM9GNUbKQw0LYnwEW0833OzMrzXx7vFQgx/feTQfHTeskAI
llMx8idZGrBJM6MFdjdq+23fenkJMqLimK1akubnf221vyD96ZC7a5C3jEXM
sWwJTCd6L4gm71DI2JBwawKgyAgk+7Tx57KbzMvJkGunzQB+1fjUUq+qGWnK
dBz1BVHt15yRt/743Vh+Y7E1RTJjsnXXEdEhefV4kVN2j/XXhy9Dcc53emb8
f8c+Nwe36QE2VpKVBEKmYaL8UujObDJ9Qf1S7eFRSm4njsx7/JaMGabHdHj3
kT4EyGFgQjlSgGg5mLCX1Vo+kyyIg+VnBK8uFmdAfDqJWe4dvrwhlfzNWC3Z
TYyqDJDjh9EpRSQtcFVuphL8OGUdx1FE/FEmKnPaSOF0Hy1R5VesqKaeAk0t
jD5QOFLidqZI8xgDFjwkP+IPlmhMcOp0acDx6yGxn64wfF3orJ3Wb+vvbrIl
e1y4OlDtj0ouUyo9jmlNokBWof5TklN1fomayFLCG8lK/GQPS1rafcEmEZwB
Idk/VESnw3cuWzqtuGRq7Evwd1xKtqC2dGg+Xa7ev/0dxoL3JrBoBzy3880o
ZEdkue20aAlqIJ3QaConCZdr1bwphAowWxHwULniSSqIjjw6B8KoNxI/1/Q1
W4hQ6O8IESnZHRGoOa2GKR4o5pSfmnksxxhEjmxS5dw296/H0mAh9UFBu+XV
lFOzvXKAv4fCUbqMQ8Yip+sjbc1ITPnuPkygf2rn3N/7yvXi04sN9vw5tNAj
QPJ606ET+uegziK93zhrY3yXxMEGCSQqBLyREDlc6hmmi1jsUzuBiT3j/ti+
UqfPwYUnr/lOjupa1KgjaHJRYZCHhzZiHChSGRapgyzmCZm1qzfaDhfYBs/I
+mqoSZm7llC2ZqkmYkxD2T7MjQitU5DOYzUGxVWNT9mGsqMnT081HCsVZDbM
ivhaR7qmEgBoQUN5d2vZ7FAK/NN6An1DizhO/Vg3Dhai/3M9g2+QvJd/URNk
WGSVQ6lTEbjEXVwtZMxN6h6wQ3Kr06FKm2IUeY0BIgonKaPJsX+0XUwzZA6V
L3zjGGQHNmt8kLDq/zA1sA2iteEEIk90YA4fCBA2Rb4E6eK81cWxoelkrxuI
HY2RhkqbaxzyjApGzvZwFsWkQfuiV2Vi5GAEJ3kQYIqXPaDyhJBT7ZQWflac
hpnq7GdeLawcieocf5+28X0twuDK1RM4+rQe2iDWea/8IL9PfwgSq4qxeaul
PItCliQIaZMQWzlSzR/OasNPZ+JOG87VDRdbS3KmjMIrjNweKn5cBC/3VdXI
37tpgl7YhzUIaVg9JOHUFpSAnOTHiUCae/b18P8ZBmbcCy4JvW81unMJ/L1a
TSN4mrY9eWHPMa6uXrRLwp5+NRyU+g20H5sk0dtmnNUXQJ7swiQ168vhXVKe
Dea+NnjVyx4Op8fSkagUdqFP+2lcwLEILGGyACIQOzVgcB1KS/R4478T4P9f
zqC/+l3OnpYaqDeI8/f4EeR59MAp4KkJsZ+WLYWJ4JbUflaXkOEe0njyP14+
zRFkcMVyQwOct5g2dUJr2p44cHrK5p51cZ0w6pgPRWHHgiNLkx6hR3uZluK2
c6OSPzAl74l64Tx6cAE5R5c6CatUh6E7rLdqovIobTSFEckFFtASPhH0HvTE
KEeWx4QjVuhnJSAW+3R2jmNBxx1/5jVItnqSHIvLmiPrv7X3RuLjPGhz2Q89
SQjmYlmSaL9tbKtkWZ8HY0nhtgleCjT5GNELJqGOEZH8ogDMSkkSQimQ/AxI
oQnzH38nfurQvBXYTgvIg/8NfBZgtg8XQvJOHANESMQiVh2ELqSi57X1V+rG
KVzBwARvezJNSFTrH9UxD96Wc3Y35hhXm+docH+nFJIV0fYY20ddm9clxGY2
Kx85AKR13ap8fD7Vxglg1eYFJi2xOEa37HaU389xsVmConcS/MZmA7ASkk7l
DsrW/9mTpn8jVxBrp8sGFNmKY+nseECnOPaArJz7x+Y2RZtfTUdxYstkhEjN
UmMZ2k2dtiTh9i30yWXlvz1HlBJXaAb36hr6T4fVDfJi7e72jVhPywSdlR2b
enes9jgqRKvegm3b/NdHvN6fVRtZfRsONrRFw6/9NYgHHTk2OWSIZhTmo6lg
TaTGkpfbEFd+cR4QrqUV4qcakxgAKuhopp1HNXAu489o7CsbXD2w9maY92Y3
gqKUGdAUi8Xfeos1jp8A6D3duQvb1kojOCztusbHMs1F/cElWdysV067wsQN
1UOKUhA17Lz9UxYDzwAXxpGJ862+OI/VHSG33S1HLnHqcTP+ywVGvoUhcFJU
LUkUWuyobltK49xb2xivJHctzISiPDvwruXliBX+Bn2inMkLGDzhg3eTeYpk
GIysOOCS84pbsmAzUO8ezr741aP8+4LE8NUkLPGfI9XUn9e5YcAi/uBnUHPl
DTgVO4gqiT6nKgBApe5wdc5WSroD+/Yd8Qddkutye0UmZnpJeTp0uOO0jgXv
tn6jTvCSuQ05ykRn1AxPbICt5UrMVgyCOF4/D//UNjnbcyzpWykjT1/sSV3W
4CP+U9u/QjgvaG+lNU6SPYhPsBEJNjgNgrHpPE57R+Ul9NWT95xuGV1wG8dB
WucWPqU7xDYlfoO069S1ql0VAFCIMVT2rA+FneH9jX8Vzp82aAdEZbf4zx3j
ncJlzHyyWFLAI2uxQHg/mX+iI0jpF23GaJDpnTGm5qyaPRZrhzGhD8h9+zAa
sInVZKKJshJrsf23Zp03kKxk6PCGYCLZzXr2ymeSrZhTTlraAce+HeNBvgGf
lXCEHg3pKQBcAkTWE6dAbCjztQuDjTv0sMAySx1e/uLQMnKdjqLKkZwtlwD8
keY/ck++mytxREcmNyN6c9XxQPH8WdtIGqBnvhPqabhAMzYQ7R49x/baoiZ8
f6Jr95Jh6f+bvpr+OhW8rMpNf2P7EOa9aaUOso/jBxa2ojE03OgPPxPLaw+2
LV9StRlNBl3M6BwOSnilsW0UTNz/q4wQnKC+uB5vwIFM/t07syHPzvu3BBmQ
Oni2F4Y4eUop+lVWTjgm2N5Dk6iOiil4t1Ysi7Fvqi/S/mJ7SMjLevXv1h12
qCnedqENF6G6o9svkpCp5HZ/KgjirdjyvYQaE7mC4SOaNtkuTKjfKRc39P2m
mhJp2vME+skeY1TKDF0hA3sBrUhRAqg3JdTic5C78gz80h8q7552OkwvaoBC
oe/mjV/78lD3ntcT+ndu7DA6I2465MXt5T3nWBrJGjxCumblPEQRVdmwaf7v
CNtFKdIy5CETzT+ByM0VzQW1Z9UN3wtRcQb91v8eQDJNrybGjiNxNvNbUCbI
7Rgbjk371qKUz713xrXNowCXbPtDiO8OlWM31J9dmp7S4iUq5jqJYwvhBUwl
qDkpGNYMxdpAyeGDd1lTA2vs4dktwWSy2TOlM79GW7xa/gYZWZ8Y+8ISoQM+
g6tV0mAS5PRRDVkg4HLI+rnwNgavTtc9l8MGdp6pZOo22N6yW5MBRbzVekvN
Po/oSzizJMWhn0I/2boc592KFQk49PbNib/nr22RuSUllT4kwzO12LtD011G
EE2g0b567mh/G9pPRJE1UEOBQ+H7HjNmrJNHjDSe1IuS6QGUSxtHs5iKIjKI
/cTg3HhlJKauPwXOXdPyC3DnAAvpz/jfpqIOrK6tpPXcXtZ7QjDAHw02YOSf
lZu5d5wPZxGtJkN5YiGdQ83FrN1kRNapzpW0W4geDyo+k4ADeBVRxPGZmASj
qoGwcnRwB3BOzRedFN0FlRIhw5KaRXoXMmPpx+5JehUYsJkdNpZyp3iYVn9w
ed+zwdjGDZyPFsgzBbZPWFKLOeNTwLcEhddVFuLG78+D6qAPbJi6UPyNH/Hj
MSVceCRvbQLLEqLb6QN6YjzszvhM4kDOI1U4xk54oB/+MyyVlShkRzybOUbS
Ld9wcTcozkZL8OnQ67rYLGeQ203uZLNPM4tdbddO2F58QkCDBchUzMdLNAnR
und680QrlcLcWIn7y8wGI+DYu6Khs+vmZRp1z1poZtjFLVDkAGvsIYzdk6Kh
Rh0tIuzBJwkEDxL+qhltlgbbv2XDvED3QRJdurKl3ZG57uO0UismTBoi7WVB
CmvrVQ7ssW6boiBHJSc+JrsvsUuOFu+GjynOChOsG7E2wL5+wmY4UNDhu3LB
QDn1BdvSfOEo8QZX02/PLg7pEjZwtWWTE1Au5HnuF2B2BAGUnmBZzm7ZUW3Y
NF02U65MaGnwRtQVAlHwAjkCc2yefetHF/94urPoS67881egVbAng1+N5X36
n8btUv1dYmfM0m+MNeWAzKujxzNc/RYbbhhfZXydAurwvy6I8KK8ZoF0F4Rh
UcJlYcvW72UC0z2Gwmj8wj4x6PDxyK7mqpTNeY2qQNadN6ks54JcXUL7r6zO
bmsWVLzyHi7tFeuzp1veNNRPD4pbuFMQLV+/Ic//wk24RWX3St9WXb4cqbEU
3pHVbtX9lqGfDfj7RUxnWqU/K2cxlkSsuPi1pay3imIaHHs8VpogfJwvWcYA
4xeSXKiPrmOEnYGMXVDPPeUYc0nxCDdThCS7NVzxXZ6CZhuYww/Ay497ix7O
MupgCx0mVobtxpMT+NzG4BWPw+AsIBStOrXLneMWZU6PgFVp2B3HDbT3Nlt+
KxhlltI1aSd1RKlV030bQnk6FNi/QqCh5T0CBV5om/Uup47NcK41h06OGEb0
gPKdgoCyqaIi04+oYZhNTp8eC5OhnYYDzWE+LylHjTXGms3Ec0/ehLNiiFL7
8TOg03Wqt3kuci4WfmstOPE43LOvqkfeAyACeyTWOCWCwXbtLvR5u5ETugpL
FVWh9wIzkbxY8nNahHluyeTTZPie25p2GntYGlsD2Rzc+OBmvaQFmhgwg6Sg
TR794g46mCgk3c32kXEVrTb9O7exYl0+E1XHoFGOr1oyRyElTFoFQobrpl8N
QMV0l7+BJgLGco3kbQB5IkhX2JDFuxv3N+fKZcHbAFwJ6PYRMwPLsxdly/Uk
DQFwHfQdPIQReXzYUGDgQv6FQDIdcIu+mI0e9uObwBES96q4SRah0Qoq5tz7
Bxwn55X8IVMm3ZM0vo6YFnDfaQ65j0IaIbk2nHNRgrTtsr/DWM714ISZ78QN
lbqch7thRXi7YvSY8B/cR/FuZz+d2d2Or4xn7sPK9QenmI2H7MYcgH8q+UvJ
xPVFj9TIAOGDxkDO+mPdEIAomRdgeprWBH+j1kejoVCtl5L9hZdrvl+MXHso
jCs/yr0hIXirnQrQy0G1gZjpATy0CpqLUxExtehokw3FQV72XM3H1VKcD9VF
Z5SB9z8LuYbcHlscKa/7ZTtTJ2ByXis7EF/2fO/2yBKjj6OL7gWZu0B+kb4r
GY/KFKL60KhnKZUAhZ9YCXSEIGGOw5fEMbWzpThaluFgVPSVyHrvbDKjInpH
+RVdXAbjgFOF/wG9Zo0zBFR1dDMyEckGi/mJwd5J9OUjRNeKp2FLmiJW7dpP
5292RvA6bKGmpjZJmzvuJ23cfWzQ3Wv4QXyx8al6bCME/Do7B+y0FD0U54Gl
0AqE3rdOdm1XmKmpEjjUaj0KUzkxBkUocKtEIEyRWUjDd4kF2uZq5KQd0ObZ
ahuuq2VnnGIJ34r3EP4+K7HoKIRdjySi3b8gMzWXPNMuVYy960xgHooFFGj7
eB8tN3pX973dhet/p+A3hq0+OUt0Oqb+fxUqHga5OGPYWi/lbM6HLEaNrQGM
IMCwCtdFzKZ+8yn7jhpQYCMqX/aMuC8ew/1RdsT3bLWkWnLlu6GiLqknTRYP
xgvu0DwopcGZiAZ+g74h7pMRbGIev4KjEuTwtqJu2jNSGhW95qVA9MuChT/E
V2Fh2fhYQDhHnmTXmkK+pAA5GrjjvJ2aGlbTwBdru6ZhgZ5ZcGFAlcVLczOc
jkDI809PJ75127nj2O7B8hknG8vyMXnEa9/XDKAqxuGYCMp8YyVjHMpLz822
07dcNbS78FzVsTrlYdAE+8B5f3FDBQ5wwUMjY+VJum5WlLyJYcykHxgS/8EY
+IoEx8NPurM2lbH/sOdP3TJFyl26Vwa6Hd3K4Z+gPThHt2FauQnJKnvvs2x/
b4Qlpt+PzmrsdQnkscQhRxZO6Whfsph2iVhgdmUaTY4vXLzs2ha6tUJ10VFN
tQh7uLYTamVEzaAq9Pb2+n2ZIMbVXUIa3B3pzhVUG0sM1/XaQr5vxtN7NLqi
AATZ24koZhreKNBoU78cS6vyJ4fvQf80WAdb/9DLey3D07uEwndgPriNttQg
Sq6FhSjoHVOKj+ZJzmPNWoaAkjT2VEGOYLwjI3N+yJpLZHRokTDe/aFhOeuA
IMvymvZStdYM21VYgwl3yyaj6ksfggqVCXbs2P7C9Sdn2/JAL2QDmMY9uPXK
GIkv6qM7zAUlMDvZahQJt41VseVU5uZkrb8G4oLStMr7XvO2kauzn4NEhgFc
dZYGy6rAP58opNFElqwLsmVjvMEABr3nw4wNAC406zVjZHDjbMn+1nBFJFSz
QS8sE24ChoSGu9MxJmmBWSgxvlz/SygubgcbZRdi1FoImZQAmy+zEvau30Bw
c0wKJXVnAPV9LhfMDJT7HPJq5fOr9b/AAzI9PFXenUma9u531Z/qg4GUT/N1
w5rodqPsqJqbK6S1rOSaGS1AyovSQhdAzRJ9y0s0wJYm2Xe0iuD/xTMXzWxL
k/e+gFowtb97PI+Pp+vghmUfjZCL5RsneoS5aseEvz1XQqo6isUcDAnQV5fs
QF7oWDoPztTHF6AC3ec9pSdPsbuneWZzauNAg0gmYhxQO/hMttF+BJTXzWzY
2g09xKp8d8vJuBcy1yhHLaC8ozYjSVhwf1KkpXWvLTMX89dnuM25Y09MawtX
+aPuU1kWtdiPXE+StyuJ488wyT+dhjmzH5rfr6rnB3Q3xmjOFXeQOelqvAmH
c1lctTgYe8Ky+oPeacUO5bNSsB1AufUuqWtLTZ+eQTwNGY97QZRia9KblhdM
DzvRRU7/Invi2ndKOIqjGkpIWeqNIhoSPHwblb+4o/xmo3N4z7mrLspYxKY0
F5Rjfi09aTsulFmXiT6oBV+Z+X/D0te7yoe9z48xe4tov7QhuShiAU8Fj9JG
eAtst3+ec+eRNvesb2caV6B2mGmfJJUrKmQb7ZEqIBrZTBjGBhbwkiYzHDnA
x9lPGqqvDgRKRCmHt3XM5QKsHNhjsap8UeIwjBLGXQ6qmqW4nDlJSjZiqcZW
NiTbs6EEik+jw2lisxhpw1rcyp0iVy8nNfZvTIWe/J9p4O6e78wJbm8+do0d
xU2GT+Ei10HSWVgtoQrIyUTbHESmVJTH2KPyp21/rElZyXnRY1h32mK8UijD
45E/QIB7a3BDuoCHPZ6YmC4bvx6b7Gch4u+9Qwwx/+LUiQSjtzcYdN9wuMON
RmmKucRNxdLlRuD9X0N8h9oSmvX3jJTHFHImURnMkxoHz5BSoFD/XuEnKM1v
MTVTAZmQub0j39HoGg6RUL3SVMvDhQ3wN2pg0i0xZIVh/xH17ClkEcCe+/65
EHbJKooIUVlqpHQyzW1tz2Xxc03DefC2N6eRBEgB7ViaQlwHTiXD1gxbHBqX
JOkaYZ4QdPqN097KnObapvYOn90uBTU4qEMO9tHiLD4Qqatqr0ZxYdobaNag
4dmkJQRUvgaHLsaHNKRS1SbBhncUILXqJjVZekEbWL808BnfJa3icO5LrGn4
2b5MXZCDnHrX9NLMUQ8Fzq6zehSrlJgBTJfisvylG79pl0Adf4+tLM3/+4sY
bf+3dV4nsDNnOYkCTjy+3yFTwl3ZuZs3i8zvg9ZVbEis7vdx0V6msCo+P0eW
VcdW1Gp1F6ZPFf+1Xq1RxmDSysncsYYB4yVvu2b7g7aFZyN5pIc8Sq8PNL+y
OTbfjQb3qUa/baJ1Ij7OSxQsdDLBIDobXzhIMjVarCkgMRlQg7nGp2ump97W
NWOYeV6lOS6uyezgHJuPNn+LBAYZB894lQGcUES7KFt/qzArYIaQI3Twbfor
W5k80BssX15ocsEIlvQN4Hy54d42BWuh0Tmy32j2Edn9eTb48T1CJOXnHzOa
oxu5629+LnHOtvT5syV5fxEIX11kOxzT3qGCIQ3t5il1Yxzaf3V5eWNgg3O+
EYRkhwifZ8Ps5SIOqTdj+oT6wsllGLFFOGhs/tw9h1PKoLRg3vvYSni3AhXP
IsGIcL7VYDllDM1Q0nhjrgOokSQOzU/at+ylSuD9cdHShgVXWo56Vi+1Hgh2
9vp6L+M/VSNF7N/5hdwJyLl+zvkeCMU697bGSbmptXPv7+LEjgs78pqYJnoL
maDriTCuYiYGLdcjDNAkVKyxZewnbov5wyo6YtlLEB5TBIMsOAvCQXosCD0N
cmdr4hMxpr6L/bjGpJ6aUZ8UbrEABL7zrHWZJbtNrgCCTqjQDTiRJqRMZAVA
BiDApxmiufT+noVWdoF6zvYVKboOt3jKjHb97SGQW9uq84mIHlvbaN5kkLXI
IdVDziyGmpxZjxfYJgc5r75F7IVbfc3PUGGGUl1y8NMkmbPUXY5tkk9rD3K9
oo04LXWDu83R7ZAyHhu8uvq1qXXtwTBcC/Q9TQxYtsqFePQItt160VaXEwdd
OvsHqSfShLyf0QTvKJaHpXTrvnhPblDRav4icGPMtnNyo0rIYPpCtj+xgDZ7
SysX9h0ied5KvDmSqnIJezMZBLt97xL7bZT+y13XGaEQuvqxC88VcLsReqam
ozkx1XpIYlYywNN24Kzp3bDLXjMvWEgNA6RD8Vyo+K0cqxhTKXaaT8aZVUlY
dgrKRkRzBXSnftFLtqtVLvHL9hokvj//7u8JzI3bat/iRdT1Q8IVxNDFZkIY
3bFOKGac7x1RaAwpF/wsMHpQR4qk0tlAyZja1WtLQpFmsqeMZX4Lu+tsHM7S
n27Pcws2N5piNdekwaLyw+myKFZvTisPj56wqicuElfdsJEtrhd2S1Kbti0j
capOcdOwHfTht5MVR2AJy90ZPdtuUbz3QUbnTXlTVExRaQ7Zxa4n1zYbGQyW
M5sU7yUoMHuzAebD8xl2w92UOA3bAxXKjqdA55S9zZaErJ1D/uWqBcfv+3FU
PZcOWC7k7F98SDjbJhOKBsY2t2E+7Z29LK/rOvXIeKWQt3VSQ06RGZan/QVh
5XdpsnLVEQEGDoqzkKVB3XEqKdHkM/ZcEziot1VcAPuR+Zz7SH1NgNwNQVs7
Eq+LCGJkB8TdGB0QzxAFg6RCTM19D70rJrQNWOtFHdQDDYdTXzzkkH1qR+gb
ZIFQiRoPg4JKCAhwVNTH1UA9V8WxuNK35K81cf2NVU2+TvHF6/Im0EHW3qnm
r6mqPaF/l1S/oqzzMLDdte7UrO7XT9swJoKfranLl+Y/XkJWZSAnK4mo9v5Z
sjFD8d5noG4j9UmwTPcRad0IYXW1gtU0G9Cd/P0fNIP1VVTv5YXZCRI352j4
tPh3Q2NHtBgHF/uxA9a9v9GOp0HOo5tMX9gpUJ98te3cY6iRUfO9oCw3gjaw
QChXRgt61A7wqURYa7iCEvI+m8woOAu8Y++oZFj0wUPc4MVtIzp3AwCmbqn6
TpTBmPy377cbydb2dIg66xqGlvlMLYMTs2P66wcOlt++zEfSyQpc+WxKj3hA
fTza0Hxt27m9Vt/ZVHH5uFkseshtkQDylR13l17BdsiVLrCDU16Wz2qavNvl
Zsh/Ks4r+ZYkQBUhXzGwTnQ7hoiiIM0A+PYnxCUqi3hQg2WHKgkg1APQ6vTz
tb/NoPLVney1yl3VstfLxXBd4hHN9EvTe6inygwJ0WXJCaNmNza2R5qVXY4B
JefcONzg/ofUwy/kOCImmBKTV5xtvlOR2ewzJ1Th7UwZOBgc7M2sWIRwBoHw
fXcXTSKKIWOKo0C80mPU8O9bS6UEwvVa1DVbqQBPK/t32Wg4duxxFU+fWecz
sdmRtqaRDT0vmlC1rt6qoldF6UO44V51yUCo6ktB2fmZi5KpyByyEMUXNpIF
AmRysJ+vDD1buhiJByMYuY72foFlWKJk9FJuJN5xBdFsFhymHw3b+gAg17DQ
ME6H3GOEdR0tRBk34WVJ91FHSW5zsE0toONUs/QZxkb8d3PBxw3ImSgpW09l
LOxo9kiON6lApt7nW3JVaZqMLDDQDTEd7DAPNdiAQDgAxWPRAb9uCgf3D2Nt
lz7ALhG0qJSRf4wcfebvhrhuNlO+paHeJ28YZoECoWfE+amm3slNjFFKQ0W9
yM9lvaUM4/YS0iG6SlUT4CrSqJyiNbAQNX4G+7MgbgL5++NvvFjFH19ckNpv
LF2tb3DLpB9oCjf0sgikNEfGle3oxneJXFJHM2WQHXEZDP5fw5sbjkeUy2Yy
uaDXkpFw709jnvn8k7HJBHvZaglClx2Bur5wK1PkTbB5H0oqhG3I3m4bUaOo
jAyOrMqxOdYC7OaKfpBJBtgODhv3JDp7iGW8O/MealFQUys97WqKneLNtZjY
piADPKdCk772hrwYKC/pEWcTVYLqfbQIEbTR01Mw9/T4jnFQ4OYPBc7VuwFk
fo0X0qQMUdsy9mSeti2jmlPq3QTJW2PR47GBP64Qcl+AGD16k72BUkGsiOsz
XMLrLb25eLc9yIpiU1BNwRd73IJfwY2bro0qcc1Zp/r9xPgLb3r9ZsmXSwHu
RKdcN0TSs7so6b/DU30edfNT2rnDl94mPjTkF7PheDN7ZssFM51HRmIhw20b
tf+f6RK0TKt5ojSfqXLWOyhowAiihqBRyEQe5QejwH0B8Wx+Hf0AE9e7zxzO
Rmga9tNXBkrfn4bM6T3IqONu9eD2W9X7FNhcAuPGxsL7TIjYZ9mJfpFIW3/F
kJ97movNRf8oR9KuVyDMk1il5LO/0fhE7wKeG80WnZq4tasPlU9XTTw+n2gB
dQnvNVFLYrFPB+BC5ZH5nKEduA42ATgFFymU2ulYssqnquE4I+hEEdhdxr1r
8EQIHb+dxoU7Hdoo+jF9fcpPxXm7AlB0lDgcDphTa407dNSH1YZ0UXdlY2pg
8pubWD8xkSUMSKjKbK0laUmziZZFKmL/xTyQ2n6ckYmrKTzBa8ga/o2aWwTo
5vqbmuAqdwxcEE6qan1zVv4BrO+CbDvISiCu4wpMzWxwwLGenrRL2GudGpTA
7/Mg8iRC+vie5PgqOaFWB3Iug2H36Dya0PMtlO6pfHp3jQKsS3gMEbbpwyQN
LeqMGD9djRNrytnebXUBbFbY2O9CtMbwVCg0eSxQQwkBfbmhGVygRKUlPl1W
RIP3ctRexMTbEcygJSV8afsNKeLEBDEgHZZaCqpqD4uSDu5x2PNOi9tVNzdo
Ut/lVq79XkGryd+bjGOi83bvha2KGM8MSobnbD4OJ02bT2vDIyVLiGv9oaww
LyiWtiPlZDKeDkWlJqn6BTbFdf9c5RIc7HP//4t09MEZq5vjMxt9m5hN4DI3
4dhLaAXKdbhas4rlnl7mjPqkkyej7dlJ2lZYnKJnHwTY18Em9HQbI7RS8lRT
wUGRdbq1O+xi0y63+EEJrqoukWwO2KxjKTyPChkD272g0MTpAYAwJLfrAL7p
AUd0+xxQXj2q6NdvGnCK2kRRRUdEP74OnqllSPYdSZaF1HDmH/9XdvZ2N/NW
ig1XQopm9yFcqaQiD0L7mSShA8EUvFc8rtaHfcJY9qAGn4G4GOeqykoIbhSU
4M/mP+rEnyWE71xkHaxQemDvGM+tp9F2dUM4tPep1cFQWeusA0r+dysIHs8d
F0Wkv9R/L/tFc8CpPpyuPn+28r69uLXK258JRj0q5YJMBKogf0aroMgmIZ1U
/eQRxch8VqmOvJHSHbNWBZodLazXzPhhJlMrnYWEkr7GibaUhWR/IA76NtQx
XMJMlfvD4pSFN8RW8BhPkMacdO5VIbYv41YCudioyh1W5PxkpKyM2dqJRun2
OKpwkdX6C+o0EEEyvq7tjhuydaBKrvSzG0hhB1eut1pclGSbtDN3goy9eXWz
Txd/xLLOgOzeEgTzE6PVtAfff8L5DGb7ou9W2VGsmloPq03kQ2VPkPp7zEkt
P2cLET18Lx1VwId6GE6a4pgxQTwrfQuOI6a1ZaNcnAsdS+GmpZdcxlvyWYQu
W/n+CM5lFgjd/RZFN1bSaznXGyd8osidLKzxZk9ubX95uAowMf1rWWvtLJwd
kUKhy4X8FeL/N06syaZQHKE5t+bfGzOL9bUm4sYcHJQXLPFLJ4IoDNezk91Y
QSg2GOdyqW443tMk1semZg4xjQh+5NdD+eqRyA15E20YxtTWqx6OKKwWl9ln
Vsvffdyt1w19AJ0U+L/z4WjOq7RHp9A2ysnP5/Sy4tmlYuMTGOqNP+2pKLZk
iGggkDkKd35qjQ9mDdwpSeaQG3NQ4iCKN4Sdih9MXAxyrjiatIBtZ7vdMeqq
a7T1gNYvW2esWu5UVWm4EICADQ5U1LO2KBvaqflq8zWjAiuv3UkV3BYYAed2
52UjQS7uNyTFRbsR4zVN16qPk9azBDRIoRPs7lqGx4UPWO6TbJbC21/MN7VG
GaLJO4JcbkyoHOTChISKCYfmGytZ1qguv54e+Z/FGhvi+glVwigkAFoUUxUP
Nreo/i8yR3yVjDCDgOSN8RsB3KM68BpmaL5UgN4evgh03+h0gGAhXEvfY0E9
/aqFpMGQwPaLhMDA97gE0njg8SWr12IiD+4Y6nqCOBNxx3U0RtNo+T8IDGdB
1KtzKJdmcZPaTnzWh5qNyVKfah54cYl60dPzR4PqhldxsVNaOmvbB5W47VmA
fohorbKLc1LXHBy6x1fszJ4lWZfUst71lSWHfUdANEoZWJKrOnMG4ZeuiHd1
OGQgYabZhv4AwDgZ5gcd7MnUrpJfkRdJLvOJx38ed7XqZ45P5jVNRfQMsXh2
PRfyyl8YP0V+eCuKI1NHqdRJAbRXohxSR7ILK6M4bBp7QfnHZB3gRRynzygF
+B9kFMrZ9JrdAMGQjtvov7adhS1kfDh75AreHvbRNSChug8+c2EgYY9ulWCR
thNV2h3wYnYHUP8LNrhmB7Rmt+WWIzLGHTYBfjaV7z4VmrHmflQ0KmynM1oB
iU0MbY7veMCDqv7cXy531nvNAu2Agd1oBxM/+asDuVqXCneKsgC5Ciq3tzZD
Cw/9fQqxRH3/2gpdC0ck9tfxLj7iETjTw151Z2X8aQY5fPOkHcZf6ezlKpkV
vMqRVC3FrQ1nQErTMWwg0OLT8yyweV4zlNFf6J+E05Dj5PHZyQZc9E+uu0d0
YVG/g+L52njE/mzcCioK6EDm4bKRDJbL0CY5XqshLHAvFG4Q7PXt55PesmPH
DLQgoinxpUoVe3Q9KvQzrQ2CPn2wi7mwOlepnzU4Neld/HPFLlm/ezxmWcbZ
v3sZd5R+vwWhKlEReYQevs7jBxnn5vP98Cjehtd0UQLOlMNC1+inr7OJLFts
eGRecmephbCtaAi9bc+Kvvart7XFA8oOGzOkr1gbl5aaxMAdcioiKz42TX3J
m4XUq1/zrKk93OiNGIzksm5boPj1inj2JRcxRncR6sFxo6OMgSASkfccP+uN
XHR0qKxVhxBmsXvq4TupF+zzrBFNwkWubsv4W6hPlwP6ywsnEXZAZPdSfepC
ZeMwJiZlIsyUbme606wPjlIl8Wt3JmyKH7IYm2f0oUShkZBwJCc9YbnI8AUo
pmD6+nzekGCO7UKCtQfJjnHr+iQVdaOu5VQ0xKM66+aC2T41e6Ed/HFAemwa
fr30wfr3NtBQUS3w/qftM598U1gOSl3XFxpKG1qkuyXTNU/dyZQcuFxgFFaC
G7QbVujYkRY9fena2FX94WQXo8ia0dqVLtJ3mjMGQDW5XiBWn7BxVEsyD0iD
20EBkGXMysECr09p15zxLvfo8xHnd129Am63NZKtne3597ExrMcAcvMb6Xzg
VnUS1kD4nWeAJIpdXYFtfoOSG3mPazqLfNAM4AhuO3USlH8efWduh5LtgntF
RUu13uK/YJw9+piUkhg0w6WfcypGlcUzrgWY4I9MvJfD4YYj8MxHpP1yifgu
HyhOGz6T3OOf/6fXd+Kx40rbGfaJg4HCWcifBk5Ur1tmaQHnlBcV3sBTAYW4
8iXvDHbVPSjlSf7XDk1EkGq7cXa8ZOJp9Yf7dvv+oZIy6zR5Mt4Y/e4v9Slw
2CUGLMeWh11A35E3MV2gyNOUJKBYFyh52TIsSM0K4ieWF7iArYtQGvfupVAb
rRYDl2jVSXSUGTI6vIx7KTPfC+OikNqvF4WgD/SHm9XgrpTEQgngUBWO+JmW
dJVxdOUI+0DYxblalpGFIXLRtXG8BxAlPefkSF3tt5Abpr1emio9ZlJtLPTB
g+M7Q87Bmw0qRpaIuGFsJ4rM6UYQucfBFifP5yl/ALCn+YA16zxB8uMRS0Lr
8S48owpKoB01pwoKqEFTlUk7pJCdv2+a574VRzW9AdvKtVQNw1s4TrAKmNfj
J7bepQPAs7cfrHWkQClk4Qf7/5sGpGvi1MTs8FzN8rYYEImyf9Y35310bZvQ
VzlbMPqGe9HXfgz6i6s1iRdDorU4y2yGOmiizi1VkNuZZhrqYdk/d1IoTvov
OvPEZGq+QJwykbO20vNtVOX3F9/TBZAIcPiXAyvsFGKV8EtwtjU9IsdrTBvt
/HEIYiikQU9nodB9st1mWuzfundNDwd81CozRPezE+FT6BKJojt3oKE8B5h+
r461FsRKqll3ufaquY6FaIyY55Rnpj6PKjjAW/xRJXq1C2vhwHtI7LsnuUcI
0tTSd6h1Ep79VJhgp1hEYvNPhNBh++yZxaapJQX7GG6a/S3aztxrdkiPk4F7
Dst8Bl3HEUdVBKCk/UFaYz6IF3VxCDlTZi6Pn+YF9h0gfkHTH/vQqBjPU+8t
Kjaa30eduOdvnVwXhswo6phnAidSLUIGuaZnaDs4tYvsqvZbzcwb23oXyMYZ
p6Hps8LeC8kQcWYUZEyhrpNDl3KGYLaicOFYhZ/mWnxgLxq9x440KCJrQpnT
T4EvN7bodqpHlcifN8EwJUCAhoiOQBm3u+Rtiu+H3XYOM/eT5J39TTRW3Cx6
qfEa/tTmoebWSvZb646ZQWDnq5IofEUwTeqJmqK9KA5kt/L9JYyk/PqxO6yi
rEs2YsEFg6Ul21gVDd5RsTJ06pUBXiQ4zyJSz4dOa1JCET4zHt+zZogr2a1v
9tdZZtDy7TRpAEHToYMg+TaEe+V54SMiGJFFsHQBhiUrnLSSOaBhwc5uCAAA
FzNq1FrnpwvkHvFRxa4n7Fc5Wp2Kizj51IPvItEgl5prZeHy7okLmuD0Xi91
ysb4FlJWRAXcRh5H+2LHlc/BwpCngroC9TOoAijsLYXRPqm0UNmzKGNK7chU
c2miIDrb8OK3UoT0B4iX00VSSGbdGUnZZERu6fL8qBa2OEUpmd12WqxSE1bO
aPTD2pGNI7oul+76ZwHTNB7Uu0hTjc/Eo5DdrAlAC4QbX/P4/UkntQ/tMooL
LY9FBE7lfSZw0gzjYX7unSdarrMHOoHWkLS6RZhLcyjrXzBApJaBeo01f9UP
eTcYeRt1vnSbPi7TiJ65eD4ffjcn8vdopnJBZqZA+n0i3HIgOniNkxj4ZvTp
kPdm8drLEdFl0DIin/bPvpZbep5jx9/C8sERNHLlYwDjEo0UCXjIDQJISJdf
q+5iTmHg97p74YozzwuLlVU/Px98LJ8UIyVtyWSsD48N4HVvu3IvO/Zu/PFG
vVgo6ZmfHCJusN5m4c0mk6s4FSZ+y5yywYg2Uzqv/fcKXtpkv4bUwZ3KIFKW
BxcbElVWxd2v4qQllIa02lR/PjIRtdOLTK1ybscxaR/N9MFg/2nNP44i1TGs
rzJzcRg9BbqNLQLWpwqBo4ebHi6MPz/eWFkxD/T34v0fcCBs1rdSnjbsP5f7
zQygztbh3q5YTHsKugyYUFA9zNltHOyutuU1ve6nukKpIgt7qIflCF8bOnF7
3l/Hc47XSB9Ex81MfpVhX0SNzt2KJ+N3/kDgi3kZjLM+ayJenzi3NQoxeCwX
4kR5JEXEHbYWEGruf73d8/0DdrWFBfGwKPoYMuWMEerBXPFEC8K0oh8jyhw6
/yhERhyglARQv3jcfjMHT1yRTlY0LU7ZGSvSQwIPJDobZzy8xdpM8svGcJxi
J4qIxDTrvSX980r0/HH/Y7ly7ipESZu9FRAri2rPUYWKq+Ijvd8PZK5cqnc5
z3No8Lzt/UfwrRg6Fg2tSu/F4OXsefOsh2G5hcovjklV3bYXvW796B7wNU+p
VsxeUHUFa2+/xC5ztzzdYecCbBpngeAGg1jjG3Ulm4aedCmQXrJF2xxOjbgr
G4rXn1lA+fNctLyE6OPcfkD7mrKm6Rg6EpA6pSRF54dgVuOinF74O53fQs5m
hl3MtYDIqAumxr6rODwbjr63YOPcj+tjMiICrjr/3ixST7D0wjX6+K0yJ4xu
5MsRKWoHWrKge+YLmKDGMRMUWv7aGmxGEr8lxhxn2VLi21HyGjeYopgbDqZm
PPJjyzcET1uXH82Hw60QQU+LJcZhYgKPV04jRpBLGMbNslBz5RV6+C1kp7LQ
ZPju2+3KeAcEkBWDmWJmKwekjYpCulgS1WpyTnuqG949AP9UXslWykRGCawQ
IOkA5bmXLVBGpbE9uWUl2HQ79T34otU3SHWhXRovAMCLORwvVrAk3jaSPs7U
Km4dXJPgf7RyizFc8/a09PsBW1C0kz//dFkPKEA2+it/y8dgXOLbIedkQKKu
lslODOXoF7WCOx/OD41jGm4T7bJQNTWzEoIKDlIlXGCv+nmJJz+a/4/KLLry
S4sf6ehFQiyqV1eybovTsGaeI5XQZ5lmSmPVRcPl/ycO3F+DHwb7bJeO15V5
EWW1h7noiT49r1PKanqPbZ+tUSVJharvyt8f2LTd4KEiGCmMqi67JtqRs9Ak
6GjVzY86wBZUixfpz8/ngJKWqybcptT6CCi1gw3tFL16Rd2cz3r8rzlejlq4
cnosQvE8Qlx+4JD58Qu38W5mVEfBDfbx5y59iipf9OFz/LhrluR3oAqEPSZP
4dVh5t8U3yWXTL/P9/Vh5cw+uwTJsNGPF2DUfJ+M/1dkIJFtTslkGZSv6TH3
N6Z/34j44rlyjD429IGAXG5beDIqrpwgLfJjgpfw5MItR4FAYOXXEdZLGhwO
Zu+wd9UhUmtoJZaaZb9E6Qp3ajK5UbD4P0GI9UB6DBQ2bt3kOMf4hsx+Phco
1aMqAVw+aUQX9deHf/2o94oQamWk4TXINZPzgFkaTGCwvlEcJhv9ntAbgBjG
tsvn8D6DILNnaMRBehahWPehPSnAloT53a8QbCmd7J4YvOH2TLrUCM80Po1c
jTyi8o1ZbxHI+D89rLQxNdLxVVd3XIv9eFyX9qbnzZdkPMWsnhgeMrziUHZW
Tk72NpKOcsJQMLJHDqE4uqp1DnMTW6RcdNGsEgosCKvU8CpjlMSVafQwbSKm
lPgVaAI5HiwZFarWvoiqsTZSdv9xIzpX3mAnzQMO7nesBa69UAglJhKpdodh
M0Gaumah9rEpd3LCNTcICqW6y1jDZBaCUURYLH6kul2Acx/YM8MBJ73dbfzk
LAraRR6C/kJKKWbpAafcrXNVOsob+wnF2jSjFPJZUe6QTOexGugDXK6huBaJ
nyN5BJWPocRg94zzuID0thOXvAdJoXVKVsUVElYAqeL99IX7Za0rULtObghN
jkt/PbVbw3Og/CAMpubJD7aF70G4IphIdhXtwnqMLhkoAZS/tM/2I8haBALB
8DORu7jxwzQ6PgCXo/iFjbaPrzaaTZ1OmYcYdd3Izg3+BFpqJgCVNX4df/zw
V5Q1ECLfzKC0yW0RwcpT3zZKfO43YU70KeWs1uT6s0/XFXnFPWWwmK9rxxMp
CJ6z79SKfJVGT4sSCaTEn8uZTMJIbj3Ijv2sCO5dO9zpdl4s2XJBBCK5JsPU
hOs6b65QZJcnvUGr75O1ZzGQy/d+9qTdNvQGmmi4y49+6eJVi1R7jBLF6Ne0
XkP53f9XibxyKyfm0VmrZzxgwmIifyajW3UJyx/Bvu4lDIwtoCS3g+DuNo15
m7anpNoTCilB2RNUCdK5CUyQEvztW6Tuws/xlAxIBoTU3nM6weIsp35uWT8s
xoBIvntRZUh6HyX2PcZ7baMCAF2Ur9hOwdFk1YhbnaG2m+kiUF97TzRmYUQj
H4ts7/diG/aTNmVCkTLORQk2XTXGmABLRMD95tCR1mFrUmpSy/LS9UEsVUc6
p9I5Su8hpt2BGuliOb4Wupbd7R2J6O5Upepgy04WogXxVC0efK+QTw0UKhEk
ZFmjiTaAywO4Y8A9k5fg/3LZ1IL7KimMFGFCvyPK8CXBvZ1+TSXj3mKAxdup
T/wofMxOwgB3w//7Q2iyzXlIZaCpiyqPPM5xg/uZETkrH6PJOjzpjttM9kXG
rkwHpGvp4VwAdygOXW6qETFyikcITcWkJHZzRtwOLPS/8dgowdPX1gZWX8Qg
CuU4rPz3Ov0JxAg+XhjDm1APRvVLCYuRjhce3WJFB3/npJR2zbORWQludilu
57yXiruHxNa+pTd45CRh0I9M4ksq0gcLpNYKcQluDzxrbd1PqBcT3mpQsJFs
NFGFmsyxd9m624//BWTzGzfPF7hjuNaExuoPObTzyP2buyfB58MQWYQNeNfs
4Bi9DELo7qCcdAdg0Ty52XZwIPC+fknZ779d7WgVVDNBK7YWZkWLCyLJ+GHs
c8gIQOBpjIdreZYuuQxjE+zGyAY0yjVcWpSHzTT/KS4YU3ve1RadWeAK6o5v
v3mUSSGE7ofleDmz9ZSBGthz6XGcFOR/9nUlIP7u1KgfzMYKyIbiDeMI/Kjn
zkfL+Fy1WAztGjUDkuaV+YkhD4sJM3ap0bPWN9MBOZOse6dQtvZX6psma7Id
mtg2qmOQGLtepQEOEoM1S0ELNd7WJ6cdcKRzKkFLDy2ZjBDm1gHKTJvkh0VW
sErTlu1AFJF0FC9MxpleII+jjqy4uC+6Pe8RMH9SR1A5XIZQkyvYXTKy/kmA
zBdKAAkROKPm+kRXiE4vCIIl5qxMPJMU6KlwmDt1Ky6ghc4Rasuop6kjFwBU
VdShaRQzTnw62U1y6UVplS3ssJ/8KrYjan+1IgTq14IL0obfDtca2IpMJohU
QS6tt1CyWSWg+d2zCyNWbAIioFDXdVEptsNja+5/Dc+thnjDwZnY4C1yoxc3
HccTUOi/7fDMqjuPN1/6tkOJ7J4Sy1Gdh/4dAe5ScDDJI56w2K+R1TBejvf8
H6ka9rixzeUu8qls0wyAsldQaPPWByxOgxjGx6L0kA+CHKmoboecKW9qT0M/
KEKtUKnjxFM0AuNxWJSH7FSoU3l3RtFI3YG5jE0e4JK8rxR/tsxEhOa6GS0S
ip5PY26WXvyIAHIfg8DGL5xTYs43oHSiwNyvltz6C/+ek14Teoi1dzDwMV3Y
thkxingZkpa1XPNrAGe52LBWsHJq+pPAJV/nqcwOHtjphodRN+I3zSO0Ds4B
j6fFZ/y/lF+rAXaR8k+ECJL6L6il7Bz15yI0p+9/kM/aVDm+tHEXPoPy4Fah
/yTbHuHMTpe14xE8cfp+e2jjiAxoNCr7aKtMWp0K51uXsihWAMKiuWhux+XH
n2/AglB6+NjrolOuBoAZcgJ3Y5/Hrp2u1WEUdBO8BdMhR3z11tyefTBvgKUM
IKdVxcgtFP3ekJJpdVScIijrUNvvdqGBVDVTkC5o413BNFD6mZDCnPoOOBgJ
y41qSdeOhev79PAoyfgmFvBKykd48rhuv6+u1nw3yMVqO8UablWx+gSxtlV7
Vv15Gmc5n5iTOhrWPNGhjD33Z5x88e87Rqy+1zQiIpAj94YPgpk/HK3OMy0O
kc1dGAJyeMqX65goBmVab0MqtdkHDubJyQ3AWoOeHkXVCp8yqEltgvtwymc6
Fl8XEEfmu8S5RjaDW3eTsDNYepVFvZzy2djXlCgiJJDiuA6UhrMnUn+O/+yB
Y/kdsMvobgLau6VTj19dmwggU5IsdfxGcAK8zu5pDzyYN7FxzmP1ZxA/SWzW
fsudlop3VDdkZunLPx0WdigVxdAkDqrNatzhBYFF0FzM3158g75gmBtb563H
Odfhp5P0q+n5Q70JhXZfWdRqByRAHwz4uilwtYNhhZM7bCc1MbooRYSoEQyr
FHt1Z0SWJnicsv4bZ9JvafOKtt7DH62t6lCM7UfVWx5cHUnSAP3JOHMojyRk
+d06148vbvTQ7rNnj0LXPRu81HRQMgNPlUoTEsPM0iaH528BDIOu4qZsWTLA
/9W8gOI8+2N4yBbhkRLL2wKDSp/xQscHFC5cNrZfgo4bAw1XIPMj0bFWLbSo
6F3/RsEJrLqx2CUzXQbSgphqCKWONwf/O2tuQaOn35HCveAxb1xkMtVKjChq
6HmYnmapUio5dnsnDHw0pBQEE7rmxxAt4TRX/5ZvN1sTHyddeKZdw+pFZpj0
5PYtbC0O7EMd1UYnpFFpL8kB7Kubkp6vZZnGfwp/42VAtcK+gu8/RrjbE3gb
qecxhY5lH0FD9qJNp3I9i7MMmSYbGwV+jy35eZ/i/9gsv+q31OvAhrpBBSr7
tEuriKO1b5ZayytFAdeBZm5UgZEAxJtFchy0roTA8EOQX+VG5OFD9QUAp31n
EfjQ96Uc4+wHqnr9ZSy/3A0YYxNcXNYoWMEiqTGj8Dri/FLRaY2Tvi9poq5y
ywEPUcTMBiTv03MVWTVJH6avfKybZfVSglcE7Q1bVvnW94o9wrxdUo2NpxE2
p6rdxeRO0hpDD47lLdhx5RXutf8TyTDomL+/Tv+bRSwRJz3cnYCflt5Dz3eA
Vc3ULzckkxcMGXIOxJmdyBgGDjU6lt+jEq7bo43nvaXqqFPk4aTs7ffdKjAr
D8p+Yw+qJ932dVSVNixoCYnHlDk9IFsJ8NW8fa+w0d3g9+XDNJzuA+uz1y7Q
A7fmqwxa+4Dbh9PT2qa9E3SAytcbguEWj8WFs0unKon3G7hT3x/f1ojKIUgH
pfSTxKohqW70vGwACI/WStzThLjPCEay6a7LaO03qV8iIUnSLZjux/CZQ0rt
iOYiqrcPMzt5fGFp6zDjKwjY1NsRIQxkEy4j417pVs8X8nZ8BNeKXzGENTaF
Tk4rIQA2SnX9NqmlezgPZ3KCp28w4yrx+wTBARm+kMwJEcRAeyr2rKx5m/Wd
dAKy02E9dfpGSw/TUWySpnMoN0vsKAIOxMfJ8feefPKhtyUL+AG3KCUvVygL
/btXEODjvxveTuFyh6ogkmcSafwFzouX2ZZF9u6WRDB+yojCX61K0HR74TOm
OzrX7GrwBVj440UHi/UWoMfysqgTjixxTJmPWAVfpnnnSqDu3dmddfMAAkzZ
mpNyHIN58kcHwG8eVi4JXIjOISDe348xDm+6SpTwxqiztzTRsqgk24zm3oLu
xuobRE4i4lI5urUdzQTkd2fe0BzrDLL7AAxvi61nzjVQp/8EfOFYZz1SxUjS
998Q5ZpxER4OB892BCqs76cYmPoLEA1oBwi3oT0ZL8dp/hjv8jPfb5o3eJpL
zoxHVZw9+tUqlyujuCjzUqeUBz7Z1egakKb9RuGxcLgzPFUmS7iBlNk/3mQ5
tltrDqnXGlUiapr8l3DYIkIeuhzFuyJmJCYh/+65kbgAf9lfs8sm8DhFq+PB
3w+q6jnXTdNN2rVlr9O1/FnMCitMjVcIkR8wcc+ML5mJKEJixSrze+mezni5
y61ITlzwcPspXswrlMAOhAVmHH3sQA0iaCEk3w0Jc/kmf+z9Dvg0wxRWXeCU
VLDV+GfcOEUu6rQ99tudUnKR5n8C4bBcdQ7FjKWeChhXGpN6vJXq1caec0Kp
OVCCvJD7U2F+DrgGjD0dMyO5lsADfHfYa9YwXOJTBhv+o1pCB8g+qaQA6HVG
v4uXXHy5DBHEAY8Zroehgcl1zAmtNR15Ic2NGebrC6utpCFqUPy/FhYYnOZV
hXkwT77/i9OEOqJb8Hv05TN3jyQoBM5Ryay9ZRrPH13e2QP4TOv9QdsJnamD
GQHvP0wOpzPAiV+5j0tQp7+Lc0N17IIatQHFoxJrowHQyPY10IltPanAXdBA
P5fGAz4kO0+al6xZhkwAJmfbU2YrpYcQ88l26+m0jLT9vvUokDVSw8asqDJV
4FwA92JlFiedJovNFvsqFvQtFU8yzsnTHVbbxKV9ALMgdEdDvtQNI4DacDM6
c5+0VsEubIeUskprtQnjyOsDgq87Bhiu0jQXvu/mriEdJ8D77f5E/Bgm/iwT
Y8C2POFy+nFZlIyMH5SIInAFH6Rh7fSxAPBI4VpO3frEOFq/oVG/ntzMZz28
EfrTvsYdLAPFl3HDRphytqlkcg8R5UsesB1HSKkrVGogt+USYtj8Qcg5MqrB
1RZPr/6ZLc/2TH2PChgA3nNaHf1eT6gFQPvT73b+MKGzeiw9zw8BXQObadUo
4A13rdkhcuoL5bz6N/fanifBCq38ymcH/GWZP/vn/wyok6JBxO9xKcTonDcf
qOQOUK6kPnDDr3k7tC4VOELEFQO4nYZBvUf6nD8zgGgAfSRfsu/8Wz8XxgM1
Q7/oBYzDH1F2SyQ8q/hE1MODsqYWthVMMk8vHIvU9GGt4zMksCMdhGyztD4b
IDMRqDnfI+U8SACepNztaQHgzKWpyxNWC9MJfe6FrbdLPlf3Hm/jAOoM2xox
ji4jPxC2C3eo0In1JKb6JfQ9Ghr/Q0DtpsbQ78Ll4nXJulIh6DFCaZwt7svm
tQ+sRIxDIWTnrSRN1A2J4UtyB2qAMbwewoLasLLlp/YGNSiASiNm2XqCh/tk
w0ptvDuB/BQ39AmG214qLdKqm0lZ0O2cfTRCrNOtpgvKyyO+8VYVFtwTiO4G
1kBfff+fe1RHH+cCe13s7FnEFmNWG/yyu8VXFY5MwouCdTwOGAqwwxUjtGM/
8VY59JnDRGJ42QEn4MyqVLloT7azB1fuLRL9/tcde1NH+S2+ZnJyzX2RvREP
cGb6DcmbVujaF4P0NpjupDTrz32jdzSJQByCHOAcF6bUIF9+k6KQaPhZT+QS
7GOV/xfe4LpfQmEfzOsJ5Ppnndqm43qtr7fMzy0BCAyFXo0pfvhc9gUC0uoF
5hnPjLaim+5k5b9aRR0I12OghXv4/sWraChUYwRztMhfHjZpb5N+h31jii1R
9SFCUHJV8j3+8cgohHDriLpCMXfgR7gIyJOnSz7JfzU4fiz1X/gUXPky6o7d
cQGmvdnd6H8g2fP7pHijgUeKKu3umeUj8ADBXJ2tBAYoEmUay1TIuD4RlzXn
AZc7qw0GZomV6hCd4SiDGYarY33EIXGib50hSxzEZ7aX25vzMTkJ1afuJcQN
x5blFl+rDZ8lp/Srbk3kAMolqYoBqYIMMaMVniLdNV+DK8F3YfnPDtMik2Ue
OZ+x0YuoR8t/hh6yoW+HgHhGq3MMgKk/Bmb0H1qR+qgPcNgbihvJmwJgvicZ
S1m1orjGMM4GqV5wn4lYQgxqxAPWninCPzNFjL2uu7+bx8xoldmlSaNMEJPI
+imonpKCpSq0NMynkR5XXjjIwqQfQQLWuEg1dwq5Y5pEDtWHFSqGDjwcQW4i
q8gf3kmfniXkXHLlqwORqz5hhLgccacGBV0XX6OKU/gIhBz+mD5ZTdnuLlXW
fOHyfSLOXBC+QA7iAHUlJRSSqcQGiOgwiWHmvN6Aw4HeTCjO1fTxoxDfrvOf
zmOwHCAwKQsVljwbcEL8w6mykzBmTK0n7IUf/m1lC58svuW9NSQkTmThFWgP
D7AbjRyYZXRwvlQOXm6+9R2ndIoLusHnuwXVZWq8L9dnFpFToVl2xcPbYXOS
mjXdK9uvVXKb6btMaHjqkHL0hQY/5Q/7c619B5KHawq4EIIil3td80v6J0Qc
A0k6cr6a9TzOywmyHa8TToMDtQNwrEL9s9ZHB2hL1tlzIugqRNCzEA66CjTB
hon2o2GWEj05NIRgIj68P2cRu3BM7Foz3CNZfpMONLsDg17RxwAGVt0s4KcT
FBxDkOHFGUmc4L+Xzdlq938PWayDF7XKEfGiDJmt9oSecdAVzqNz8Va6218F
saFdYMYs1j746jG4QqL5ud/Gg98EU3/qY88RyM1oxchI1O93cwQg6xLjweUF
MQCP5LTIy+dK0FJqf8m6s7j7UL6STq60YXCPjC7XzcDqwpk3jY2B/pnE9jjt
ICDW03AzvJjJkwj4s9vKE0GclxH3Cs/PpcN4KrLQbVIxHzpjgvSPLt/ajVGJ
eZMV31z10CwdfOj623x84/4877IdA3U2Wtau/kodejfLigscGKIIb6dCxJF4
OCikfKViS/DBte8m20RPEvEUVuJweZwrULxFoSNrblU2J7k3o5SwFO8Y+rAs
RvC4O0vG+gcEGp2Ehovz3luCSMa6dC/3jDp0FdYYjTNDUGlv4xfubQ9qPhE8
qk4rgsw9TZMrNt8EVfs1UgTw/oBZlHjoc6e3DusrAax7ZLvLdWtWM7So5YTe
okR/27jFgWZlV15SqdPkkQI6lyt9P0iQAcbT+lGaqjpSuHRkqxhdkMX3A5Kx
va75THkMY9Jvy9rjrn5Hv0ha0CO6Ayt5RRWGRAtxTZUUP4czVYZs08umCjMx
Kma4ljZYVpmIQujoepnNs5tKQ12KSV9plYCit5Kdo22ltBSVTEeEyKJt6H4c
2kJy2V5WHA5msrM3ZCvfHShKfpjWXt7ivDBotgEZfqXde4cBzdD63i0CEFWR
Uqf8uZ70jkOXPHt8w/ic6EVtFdFKHk+RNcm6HJcVqFIaQoy2UWB9DcBGx6Q2
LLPRDOLXb8LVa6acOSMdO9pXWBZ+RGFYF8CsA7Fcot/66yYOtZ7F7CFV2Qb2
ylnXQtcYjL5ZCSx7K+JiH6YvD7P2XVLVhwrcqnhln0rR/OAYQtcsJc7g54G3
U8ZwJUvprw+UuCu730EV+KagW1m3ccCAbBNX0v6RY9qScYDa4hDcqfkvnByx
wMELzKUWcwLmHjJPJO6zqt4XGodxBugZCvZ51+QVhMZwRduWXOAUFR4HA7CX
l4R6YhbiFdfYcjFC08hFzJx2iU4qnYmEn9AIaJJFfne6xPOpM+D6B5jOlEbw
LSmJzrmv12nn33wFrsz/ro791IuJnSz8BqKLnDVrFiW995o1W9WUlrUARVDa
whwNj+prov/GjMHpdcjoZDsr3f1t5aY/tXDdzMCItOn6nTlrwiAfbArQlHma
3zeAbrYy+dtOjyfkFzUKs7fL7kwemrQrvPApgZyqTsBg0FXyaVqhqNhG8erh
AEkJeNgdcH30POKdsQ5RVkRjhvPJxXYTb75Sxnc+DdJy1v4+RcjkbZsax18Y
U69sWCwESZUJQUZlSmMTrsH/OU7lAbDwd73QqfHKtru9NzvQ2R/m5RW8G654
6E9KM5Dv5O0Q8qLOgvXZlyfhtrfGmp53X/8W36dS5xZ5rYXGGJFmGmHNDMWE
fECLjt2gAAYqTDQzR7ZCtSNZjqH99O+/5iN8AiM2ysACM4uHjdekkVbxImD7
mjnF8xVPuCYo2f/ug8Cuq0Gn4womSolE5je2+qBecF8pJaSVgE7FDq/BJrpg
PXOKU6O4A4641lpqiHAOsbaGfeaiD4kFQQ86S3ljajEtNNponOzvzgpf4oMG
GG6yFLFwzi09gJB9uvuPsRzXQq9we9FeuPOCTNhKsEal+4tP138OdI6Z8xLF
CcTRIkXt/US2hKqBfkW/Dg9pCio275DUU/DEKSpw5w2HwfeXG0HfJglxB2TL
TgVu7Hv78w4xWo3jMbTitPWiie/pergQU7hpXwNSzqMJIMa+MIudK2s8iKKN
jq5yX6YrNsnaDh73ydX6dau6DSeZ7PuJnrpFeDzgr7dWLyMZEZ46c3/9vbW1
5OAOh4A17djeKoKNLwvYh6NI9lmIWDRjeroDJ+vI/X9X4+8s0Lv8ZhFw1acG
hVfycc3qFf8RcQICccNGKW4/TQxWgY3086SNkCiX/WFFoOzOZAAJoiEy2r+V
W1q24jouB/teRzNxxuf+18WZIRFfgS5O6UpPmf4wez5m/JXvqGv9jsJFspaJ
gOYmLrN/HsuoWCPDDu36VryC2T2eBgHvno6o6tqMcdBSaFm9cF3sTi0cL4J3
INEL3S4Z3IVGXdVLKXUxjyCS3QPv38Ejg/IKhKgDvoUjYKhhfRWkEI0zy6FL
6lr+1HBXsFcfZWpMP+lhHeZmFd/GQnMzj8pA+tRGBc42P9Z7b+DYorDkfIIb
R6GYchHIu6yEmbaDaEvxXbJu9fnkZXS2VvXVhvq3WJXxdkHmQS/YPneDcbsd
VzLEitymOhCvybI7aCAWM+tjsYzmBJlf44YvJ0Xag0CfG+iITXQXY34RxwX8
qhjBR67PjaJn8nmi6ei3ST46SuauKvuIKKC13v8eF5VK14g9hKvxYxNa63Un
kmVXvN/bnlS7l9UMIk8fDh4pp92XBnv7i3HG8nI9fpeuQ8dwEUMi/ZrzKLWU
g7KBHEj4lzBj6C3oh+ihAsLtDM/0wNoq2gO05OnoJfTxN9ENsRUGfXM4q3eN
HsLExHuhyE878bY3a22JanQRUajvs+xBQ89+XM0tWnY3MHuZDQSmrLFBwVII
S2ooJlgLm6Jw1kH7PshrvfK3OavaC/EduvWrF0Pfw5dBtDmMyyxriHvan3cG
ZaY0gkDvPEDKakGo/IWzMfmeAfivZDLp6/8Wy+bvvOP2zcytSn3gxPUc2xnC
5PPg0xSattjhyMFSvKbhi+6TI5voaaauMAvj/W+vKOVB8lSD2g4pFlwnmRLl
w/3ksVyAWKUSx7Jabpj8F2fdH/CZHIkE27lYoEhbbUa6ZJTZXHoo/whwqsiH
YiP+T0hCwu48oI0aea8CCWvzACke+x7Y9m/TljDsgXLk0S82Fbc9JI7tdqMd
s6rq6Ss3sqEci+ZEyI+QTsARaL/d5mS9iRktrZt+HHEL+PbzCy14glTYVSv2
wVDvhRCZFI2Dpusd6w3FY46w/qG8rbqGr/tBDam+3PIW1GRmGy8l3N+LCJF6
6OKPpBE7RdhcA7Xw4B2ipCq197Fg4XsEP702VBykyAGZxmJ7I75EpxWL2N8m
ek+yxUprRpEHn68cPufABG2of0WYh8oZVjPk2BCBRhb7x1Xr+zyAIYILkBEq
QvQk1ebu+fYBCAvSuQ6iiiVPZ4bXrIgCMuRw2byUWKQsVDWw7PWXfWR+XZvo
3+dgTnVUHi7U+LEB1EcNmeflqVYgc1DYFEwk9RMKljw2uVVJpHWhDzOxP18B
JTdWMW86RD2yIS66btWliS2ZdoHA0DaLyTaCt0NRtBanN3bjeMB83tyePOYN
sj9nVaeSBFtFHcTiKF4VoSlA+PuWQm7sSZA/YQi7Xe8CPdgWmqWyE/6OwmPN
YSuOoiajrkyW8yZdQ/R7xn5P4y0NjcKxZGWGZSYPDO3IPxsf4073qQJ8GMJQ
8bJDdkHeFQXBbnDJVi9O2KvoKiDr2QGRTzKSOWK2JpyDrpI3OnVGmqne2R2I
vJenpt9oc40zqIrjaDPCQ7KhGm98jdKKz0khOFNXr//ndT195Nz+XP/CHu5R
n5nQXSKoM3kSFjgjQBYrmNSPZnPtTjLKyelV191UV6AKEPD5g9Ac9FasMELB
F9HQUeYV1lxnhWgMam/invT0R9WwagS4rIlBpqWajq485L85RWSWVPidtNFD
cm84kvY2VFaBxZ/FAfe0Zr2jQaF9vOryKUBnBx2g3UZxv2KYBE2PcSeSqe2G
S3g1k6z8lwhZ1hY7p+Znl8BlRvAl4Ooy2TjZaudOSemF0elbhcgxN3nucNl5
esi47Nqe9qEdOMc9Lh3z8rZo2kzbxMSewEy2NWztVp7dRClcR7e9QoUrkMp6
CNccsmS7blk16lX92q6tSeiniRkTKJrnuWxOjz69mgNwYZt4PFA2zwI1OZCx
XNSxmXV+aBkrqVb09TbRoywPaHQqiprRyB3H/GRYdxMLS7OGKotFxDcZxwoB
0A7hQk1QoHQdBmvW2gXy5KfP7K4VyhcahFR5ZeJjYwEBr/HNXCTA5qjaPZ+o
L6S79dwqvg4vHmzJVQ/H5jdgTRunnko3/9wuij/zfMfejtl3Trn5ICV4bd0r
Xf9bIv6ITXskT6vcMLEbOiOsSdl4D27yF+fs0p6bM+t+CrnPT4pmW8CBmlaT
0QOQSkfF8iyCP+7i+hPV5ktiOmZFPU7EHPOUR7fOezOtooZQoI0dlFTInSo9
scysh+i3SGMI00F2IO9gXMU29YGKovdttATc6eqyE5NJgMhbupEwlJtMAjPx
zKtb3uMRDwHup9ORhC/LmG2wDGKioCMcU1pnr0HtUVR+NKauYsIXhKGkDdS/
cVv8VTH2+JQqO4z1zF8hpVYF0eeiDmLbRpanJpqiSXxxyz7WimEM3ajmIsW3
YEz0g7iRTgiraTnniqOJWkg41eANkWly6Xg6ciHlHdW/mhIpICVNl93CvhtD
oT8LDKh6MHGEmEEYHwCfBCT84pR3YCFjuPQzSdrmjT+I0oO1fgvUKmiJsTa7
GvR2I/Y5ku0dti9ggyrfK/y8f+C5h5FGirogM9cPDcDSkSJdfdsUQZzTkh1E
WPADOXGzo1Ih9qmorEKleW8F7CfSoL+xTWqhzGfYj+IJq99ciaW7q19YmTd0
KOGXcKBAIN3jYZCsOVOuhg3VqcCCF9NTfES3dLCMwTaWOEM3jZplt+5IDnIn
wy8948mocLwsld476ofC9qAvNgYRymippEXaW9NW5tgzh0ueuaKg7UCeKtXW
f/Szmt1ohl8w1RzcV6F0B0jR7153cILgrvnG1jURZxJUVdd+t8wF8ML9cCJX
gzcQ/+w+TdTN61VT64HJqbrkAT4KEQXexIKXCbR0wdaLjH5KedjjvZE2+9x6
MKT50ZMr7M1x3Gd/sLdfCH+in60wDcv78e+dQxhHN4nRhDtNUQBgp6CH8O4y
QMdEzKi5CYW8BuiZMWpZJQPHl271bliRXp8dLNLncjsQc0CqIo9dafIKedGu
NLtuF1zMFKc+4owR7YB3q8zo6Z7pdJzpvMD0eaSPwSD0VfPGIIRqk3NI8QGj
wyfb5mJhRixM2fyZWhh3EG+a/qlKNgOSkhqsZlrY73bYYQOvP1e2uxB8XBj6
Se/NNxheTUTLgT05aYFH5Xnw2ezwYPUoBJMAtg5vXkfDqqKDEUx4z6SJz3Ny
tZzMvCAyCb5hAPydnsiVMfU8RQJSVwcwJBf/Sl6uksP45gAcPGyk8/VH2ucu
tNfHmA+H2LX9yAg3vkB3FrTaCf4ba3oxyCLvPZCoxagxxyw3ZORYrdjM8sFL
mjftudQJdFJxfcCuHMJhjzKtfClJlwBdEEsLG9TT45YNyuE2CSIk0maAAlPh
YCm4tTtSLs4hk8HCS5SsOnOwDQFh0/ivd8dJ5gRkdeXuJ5od1A8Y7kVuxVK+
W6iakmr5+tpK1HXYiwPUxpvinNBjPQCkcfD8jz471/UbEEF8cqzcFNK/pl19
u0Q6UtFhld4aR/7dcCE0FpiDx5A54fz4wkSaUOoggmScRgvQMqdsFLwQpWdB
YX0VIql1EJm/Y0rHCJYNT/98gRY1zlOuK0Au6yEt/GXPNpmH46tHMvUGNiV+
WxQWiX7vxzXbF21Pja2yWXOg6zyHXVlpwUYsSBFEaCNrY9TwW+8OsKW1q3We
25ttTn0gStQP8luniwpoACYYdNw3m3HpnY553krxQCnq3NoIo3yA5TxPilgS
J9egeYFreqvbS9mlnqbH3rpCmQQfebK9Hl6KgcYC2Eb80uykNDBB1Hc2GBlX
VU0WdvDBN+sLzB+7A9KeqTMLRl2NETgiRACs5M/lQRY84CaBaLp2E4PTBpGB
JCO050HXgnr9YhW1LWr/HigZz8GDDl1gqTwzxhmiXg35ul/QShmgnm9aS2Cl
IrXyIKsnv45SqNsNFQCM20RXYfXuwVfUdqT9aYlVADazPO14nRxflS7M8jln
Vb1SmhqVee5CEpuf/4oPaFkt9+xM41InHxGR1rY/GiMUHe90BdsGo0PN/Nj1
4h5SfCh6QarZXpXZzwo4qVhIImKnwlv1IW6d/G6PmDBZkRDf/sjLr2uiiAwG
Hxe9Iwxy9yJl6/DnWJhhbMApLGBKqAFg1AfFER5mD7QbC0gNhm2LSCiRuVkT
dnFNIstVYdxvQHA3lYYjy3Qpis52tJ10MplHAQdIlegbQ63CoEuOpE681g/a
+VsZFUHT4Pw0DiCAvQIXu+/NPkcTSUdFFamtpi1IRzqBw3z393DrQSd7Y1mJ
X7A7f+gjinUkXxv2bC9eILLe1nMHHzQ+fs22AVjfIBBAeteNzViDOuFNS6j8
NEbtg9MCJQrzW7g8r/d8Ixeaid0I+wtSMeduRpXKGvOBtfzRy23+7PmCwO/n
orGvZpzNvJFWREnV3tpWbjO02lpd5VGKEznmoHoZ/qDQMB8x4EPJBknZZO4f
EzgT+OLv3yr8sE7qMJNEWfQAbX9ki2UB/3RUHoMJdxRSptKGSv0H2HErAQjC
foHbaXS4BQQig9IiaNsT1WdNsS8BXJJpecDoRhR8gnXZDbAXi49bH4Qz8vKz
//cG6rhqED8EyHFMv0qxvRYHJD3pdLMrCZliOhaUB3DalS5OBMsSh7pA5BcA
MFEFQgJr9+WbNq75feocLAbkFY8BjFKIpqgxHHgW/6mGprYmPQpfmTphQnNu
IQql+Ivwl9kndgYp8IO4E5pK1E6VRtb+4dq7LQ+kU/Y7mqTYIMG1xvWH89CR
IM++vCY949js/66WorFK4cPZlRTWqyHpL71+A4vizP9SYaTcooezOlB1RiUO
AQlnEVkM5ui4mNTHfe3sYBVc+eg/XA1qpAccjY8AefPLlAzSX38a2VVEzOP1
YPmrcmrl8oRyRS/Yv1LJmPJUKLvAiH31Ffvl9+XGIAKSKPUNrEyEI8nHed/4
sT5geY0XavQexofB707oFkzb5x8Vj36Tx+GEFovd3J9bUxOxOBiBaqU2X6UJ
Qo5i7ODGDNVhJcM4HljThLXUKV9wnxOzh8RQjhO/0CGBuWphN+D0NxzYN0MH
pX3HLTZUssXiaTCR+n1Y5VhvYwTKaRrcepdnk2RZ3QlMt0yVNTvzkwpXyHJ0
H7wRMgjvH6o2f64M2wLiSHWA83ey1VTXOMSYGx8PH2GMpFWk8ZTLPj79UkRa
BkoW5W+gIlB7QVOWr9yUKpTYh9cUl1v7TlZ7PXhMmReH5Tlt9XMGiqMOyD2y
UxS9I2EMPhXE2BdnwYi4k01l6SCcd5ZOhHa0yCLrkwr2F35jd2rZxPJPRnoD
I6IgkjyWuTIhtVKf380wg46gQKblmrlgdisfDjVokeFiaHkG/jt1OM3XvnhM
mUnF5KkPVn4s8VA3T4xlNqCUcAWX6LVToLVog9mj+orcmB+7LVfy/CaS5ENp
NTHVVYIrLCbrDgqFtVr84YkEQGL6WAaO/1oUdkd5qh4TFdAQGzo31BFgMHQA
6/gaVwzKyLEOmCVCDzIwO1K+PXK4a3YnBuNr/qn+MGfX20Zkhso+yB7XLj3K
lN/6t4L6An4Pikx9I7PvmaI2R/JE9prM2SzQQc8bI2lr6dQzawf0oyespl9y
EE/KwsSvboJHl+q1QuEhYoLDKZFlZad1qq2UGI4eyx/kTry/i2eYdnR9IR+I
vnn7HfEOL/ZdM82DSeuyL9o4dnJcktwyzdHI1jE9tutnymL9vLnFko4hh/dj
Ow7a+nEVuA0l/zsVWDYJ9KWaXLasaQsMcrsfOzgw+GB0VABE8egE0hl+PC1w
fFcntpwdiJJRdDqoOZUDXUeNwXxTswEFf7btmDf7wG88Ue/HK6UZDZUnlTNS
3ifFhyWWjZPgoZWCcRZu5WEhToCaIXJ9tQvF+YDDUWdBuc2TzMkvqt5NfLma
5pkfzrjiWoFlPL66IWLbTZFB6opfdNDkI1Se+N3BdlHGVtOhT8/tKdDbWqPD
KCOs7Obxtt9LYRRN3np/RgYzRPm8A2f8DCVUW3+u1A5OsApGjd7fsrudvkFx
rsFjAK9YmCwN0DceyuEPBoyCUhjxlmzSqE+7PMaRTiAEM7nJAFQSkpPRyzJJ
f4rQtXEYUAoHicS1IKMik56K98u9XNGJAnrNw4HowulCmW6m5lj3U5SPJArK
5dWAKqlRGkza39M2vSGh/MWxb+PedlxNkL2hNB5+jDfFZnb3KddQfXEZuhsB
0hvxPCikmAtgE2YKBTg1YK6vzafUw66ec+fNVMOHEQy9VdY6i/sitzrcBrQg
cXor4j1zbOefAea8zZW2s5M3Gs4Qb1/hu9ENbk/DCkPwln2FpGGKQX843OOl
sO4yCYpU2M9ftVgnBAV6lr8WRAG3ll6Dd05xZCnmSPDNjRrfRODbc08a0Dxa
NpJDvL0lNFEFHC+g4Iyy39TuyFQEGOzhjvNzNYRWrn+uIzIrxkFe4JSHeilF
KfZf6/3hpZFMVPrdzlArvnk8mie5tsVNKVPJpnNs+5vc2Kl3xLQxwCLCODMH
npx+fyB1YPe3NeFIgYilX9sAqamL8EAxtoMidkXyP4oPFeQungYh9ffSHy9f
2/y7OHvvhxEKVMR9rDAP2koJW0p+dUCw9TK7CGoc0GPIJXlsdwD2jqik3R8U
rZR5pXgw531R+N6F0fpgBKWsCUDvF3dvXDSvrY/8RgS/rH9StZ1DG498WFOP
tMUyBHSdqwZrSGL11W/aQrEjXwnta/dUME1a2vTkVc3bmYoohatab+Fi7Y7m
lI3PNVFu174nKDlHvzF2FIuqzdFz8fXzTmi4+M8XvQXIQNE6hFm3jY2BHoXV
At93tLT681SS4UC4DITOuW4GrwFijQFLoDcrWnawe+Smu9ofaCv+Rl8utxSk
akXlA7WTK6h1ATScyOSLAQ8QkanuvId4yKvR0M4+9Q8j0zkeoWeAVxDejFxk
kmRa4ukroGpjmtfPw/HcS9UPZR8cVd3vZW0dBEQjwf3YJfDhC2JkT8yRHQ7W
oCKVkExYUpBi3qIaV3pLTpKMHK/vT5Z8WWly/EqPVK1mg4jO4lLL7yDw/I7i
GHBxwLGTMYI7C3pY0QwbIidggh6tSa/K+xod7S5W56oVZfV0xthhdap/w4qQ
hn28vUkIIM6sGR7+LfZ06IqZDF2B+Skppj7XyFqiCkyD1bzx7RTqyjMPMMdY
UL1CZLBaxo1hFjYVnkHqxrTA9EGqUrXemXwvLx9PEKlGNIQb7athC+E65AfQ
29Z97s1qnOdUvz4I0e0Wi5oHq37W2H7d7pohNZpNBjTMStCmVIuj9CrDuQ2W
TDhNzFUGvPx6h3fWdkd3yMoGWko8wfYGtQqiKfM9+OyumuOPiNbQVHjkQUWL
6JyFARxd81kRUyCvz7PZ36U/2nnA8jdI5PIPtOn127BhBfqpEdGINxXDXUwS
fY0xvV1dENHypyhW/eaRCjFVg693jLb4wbOsbM08Xw0qs/sRERJovU+ebAm+
rSnozM45NcdcK3PUrRAJIVNmbaT1k7UFGBmN0Rpk/oKYBdexhO2NNbDcK8wR
fZCSJ5mJ3J8NDmgGCmMyDoM/NDRieggDATFyT4xsmeMrRq8m/+kOCr4N8eCV
rdjSrKrguKp5wPgPhDzyZ6UV2gDxC2uVQ7jcpflW30mJmtrFTEPwDhBp/Adk
n0DXhogipFc+is/fb+zCsl0UzpMsFu7nXzSltJOhJAY4bMDrjc/3mxc0ASd0
8Rn/rJLIDwe0G1QWSLDoStXI6D4fVztuThM8+Ym2cLgTKxFYa0eGD8OP8Exu
aaFhGscUAAXxtWJHGkRZchnTMIg/WUzFZB0BgpQ1JbuZX91ePb4zW3boWBrn
NYRdi9ntIpKrax+x4MNgzNpBEO/bTc2mJlFsDOsjK0cqViEh94Ova28jBfam
9TKgGnpdALFNZsRwAY82UCMX91hmSy4/BN/oXapFH91CcJUyxz277NvYmk/q
lD0TkWMQMFRgG+k1p8d2N3IgOeblTStXHju9/eMpxS14nRsurrsn+VA78jzx
TbG6jiN4LViDrSNR9x1HQVKZ3hFUJF+HdW93IkfL2alaU1XYDJzwjYSWBeHA
6CHxHQYUAllfCOIaZL1XBK8edKqOf3km7LIKi1XmUnnKxVPNzDDJwI1KUSkG
jW5CqPFlUsa5X9UnbwwEpx9zURh6guPz75T6txfaLzgqtPHCHUJA+ldU0tpt
D+BxqSz+0AmlcEkHSXzhNwluZakHD+P+lYgoNux/AOuiUdKTcrL1A3j6w23h
4e2k+sYWNWRv2dH0I1yXNNN7p+b7KNbNCli5vRglb/zsjtLrvSdZHFoOCZXm
wNMqBBHiDDB9g8zLisaSMRDSQR3G6f8FB+tcuswR5pfGyxlPFpky6XQLr8jW
LvTKUN4XvYsm1oF4XzU+X2QEIjFHezxlKc07pXKmrfb1q9qGcK21w2OIWEol
5pE13y/F5tJz0m5gTxwGnc3klLG5zxrD//L9Kx4lj+nz2Sg+3SfRTez1vUQT
WdbjaYmeykYqhaGkuTWXESaq4TcYFX00fRXcUs/xg3rS8A/wr2Dcxik0NlK5
t2l8oenYUeIAXqDgL0D3rkAshqtCbW8IOdewPuNmQw1PW5t2k/pAu+ST6Zn0
FMrMk0HdRKhQVrX7g54iXDZsjrE6vvyTmDkKrD2u+C+PmIa9eqcpBf6dxema
7aap1vOOZR6IggKBY5Mo+S90Rk6KwDUOT+m0bvLjBtWxVfF8LtJg3kuhTFW4
tIM84glPyqJWK9a8TVnfoudHmLckRlu+oyuUPjt+6+lDPCuyORoGu0+FggTS
1O1Gp+MSlpN8Ogpv9L5vqFP5aHOKJ0VpU4hmXEvrnJQhdCQQil/kjN9P+JeN
v+7MyQ/eWWa6Xxggxh91QxN6sO70iVCTGtccDepQ7wHlTJE0/zJm6VeSRX7x
SxWS14fw5olOmKZPfnHyC40esuUEyYeuUK3oD3cQvVqdw7m0gUXAZPi0dK9R
p2vzroe5FqPkPMze8CALBmR1rIjlJ0LOV+Q0vhaCwTeLSa3Fo01KrFNHDDxy
3uWEt6dPsVMA4eXsdhpfN7UB7kUYS1WuYcsoz3QzrqHWH16BH/IRikwcsFqm
B3UavQQ0EBpZG3sifm3lGBIdNtzeRTMGBb9KPF/JsuA2w8Auf9uFDkK3LsK0
kABm0YwSvI9OoVLbjZT7pMXS7h/XVEi7dcPmFdc2ZzIRZ5BiXoQ5MBU1Ryu4
Npl+Bwvwnx58oUtZ78mOLaCIjexCgpWvPntHf/xTrOnHCVnEOm/7WeauwpJY
3TNeuYWMsvreWgXjr+bKZ0cxON8oJtrZZcJGf83H7xBmzxe2ykT55II/hgp5
k6W3TNxBQUtqqjZDhSY/paSXrU7k98fS+jFiUYDOgSWup4mWFI1RzRW3OAKN
PkqAqULmk62hnbnp17rcwHxOzKR63wUgHY3BW1F4+0h9wHCuOg0g+W2FbcyS
s1PlsThQOQPMddr6uV2LFvILOH3Jo3bBSrKWExoQR0G3OaZcTD+hYU1MqNXI
PX2g4LqYZW/N2WEnGsEeziLmFK4GlIA7WflgeUyT3C1eHSnEPLHAKF1JFOia
xGH5Ndx98BsKhTX/5EM5bs5cMpE8hnzh3udY/uydN8MjvtlnbLnIeAEjQyG0
Ma0laYuNYRMLNsusTCUr8QWlIjrGdcr1Tex0cQwk2IYXOcLaL9iBDT9jlOOQ
r86w0fsGqG8yanCwFelM09CsUHOM1PJBYYKRgfWfw7X4FY/jGlHhj7MO4G0S
xwDCf9sj4TO5emMFxmPw+AlkcDMAq1hC3rl2huiIcGiBLS0+M+MRjgdPmb+k
jZnqmRGpL27JBTlxOm64g10ndB95DbUvMgki1Ll63j3Eg16kXi9AKI0Rh9Uw
hawQehS1AUyFuoCMXQ2QjluJzTF2Bwdg3B9XyGj66JCYsD31+7ZDJLF93JXr
Y+9F47MXABLw2KjimcNheKBf+/k4MegaTgVlnFJcAUyeUCWjKiBvAZIOLY8+
B7Z7YrRDSdrBPKPFoNwUIS8v92UhVndC4WexfR8f7C5zJuMKlnp5iBosTCda
dPx1sE/vsF9y7rVE96AKlEzpafRwPqKmjdnWa4wuZ3Uqz2nAdukb/aFt3xBG
t0xtJO3RauIIPeVV+XV2DAJqJOIaZ22OZaxecQKm1cLA9B0jGBW93yNY9RTN
+gD6pX6OQ889zNh+Jdppzd4XO5lnUcEXJFo6531XEXoKX77DRjoOayyf1rO9
KeSJ4iWRJab7Jt8QZDX9u1CkUI1Xb1ZWPfV8BfimNevR+cN7sYVBK3LCZF0c
5wPo8WJPzJ7pwRwovQBiGF4v1/HvdQo1I9HRXytBul47jt3dRuVlZVGseKa/
4oEYV9N79bYg+TJoyugw6UkG46qnvhqO1stzfkaDTUfLSvBo9//aUxuugRGA
jCSrnpw6+suIpwJ3hbcqGINQV0mQdIUR/pK+4ZjUzF5ASKP8K+AqTvJqSodG
RcgmrMQTo04knnsl7gFEvxaArIGPytFk4pS6dyRenS1++w0LB/AaYfD186ct
ZhvvfMEzU0dmnHWAo9BUz5t0gvjSICQtAHpenzLy+JKzG6RhHqBasXSofmZo
emkPiJWZLBwloWNZ5RZrZ/ksi3DkfPuRcOkjrcncMTu/5U2yPQlz06MaYIBj
450upY8UjB8FfneeCxfSfDW9QlIDCJzzuBZRkkijIE1s5E0GupYNQjNY4g/C
V0dTXNyH0fW3E6GazkK7J1FG3WBaeU2pEfq+b0u1VCveE2ueMbZsbV5FIktf
3u9L1CARAxsCND0ooCVY5pRviU7aV8+Usbbxv4ulZHVVwK+5UcSTMhwABJzs
9XXhe75YSKO0KjRTwMiXCEt64J33rNaznOlMFygjroQ01fZ9PWim1QxLu1VL
VnNvuyoW+BeTtjiBELd0opiSIuSIrY7XCt7mrjnCk9U0UelRURdwwDodNqtW
8OONv4v3T/m77y5cseWw/KsFODiw/gf5joYTCP2pVYfLC/kg/BOVT4WYTqH8
oOLJgQLgvzOjEOJX3JYTWyvMDo3zIxcD/ZMgSzyteyrvm4EwUJaIBa9A04HS
OU/1Vt3xOW2o1962lE+CTh64VNzUX7CJ8LtPP5pJ6vq/TpBtey80O1PQTC8E
1byohWBuh6QaU+J76ZLjITAfJLqtdHbffKTzHVogT4kDoz0LkVIKPYZ2smhF
QSyF2wlp4kF5Nt/vdKQyvKKxymG6xJ4qMQ9d1rFxlmCGiVWl9PAa/DB1lQ5P
2DA0R0+hYmoKYN5EA8y9OJYOBtbTq/VeD9n/GJJxWu/Qt7+el7hXRbC2YohC
mvQSE5cLxdJJc9cEpWZUnpgxihuEbBWF+EdBzYS6YNCCpaGaKJ1Q6So1pdzG
q92M477o0JhEIIcjX0xpiFEd5VLl3SfPH8TGF9VP4Oi0NRkyM1OfNCyey46b
L1eZ/K+0I2/pzz6Y6zn2vx28n5xcErqgjaqyQBy+dD1Bq2iom98Zkn3fkvNg
P5DNHfNGZ8tO/4A711uoA9Ei51nQn7h2tAFL+NBRrw/i/sLHolFclUqBTLpi
VoRe3LPtRofy88iIMK0MBGSr8fkOdexTXCGKw5ZmbYEuElthvtqF+3PMK7uj
ChtgCdF+2keCSyHbKsN8lTsGD3/3n8vbv/efLcxZ5B28KwK1z5355rhR8ndw
1gbbtfO5tptEhjErvMyJuGQmm2p6oPW1cX0fw0n5ossEG7/0bUUvpA2BKiw+
Q1uoMq0Tq9y0BLtvm6yEUDuXdgOzkQU4V4Go7uASTiMMgePfphlUdWkqOFU3
tyuZnnAYYLBpxbmKfBluoaunn1+vfLxKg/EHTmOB7ePihhOa1GowCF4oYxp0
NfhOnV0SXUsEqq6fj/pFSyNHvIMr8MNAn/4BlQWBZmX/8gpZcH3SQxQhf33v
G2/TFVcGDlzE4JdVhFWltbXVmuy7nRKo+PDg+dke8wmeedgBS2N+Owj4WBvJ
dfbDJbmaXqq/D4+5DMCIDN88LLWTlKH77x8QvzLYJ03NerAnWd6bSuf1IayW
FQCLA5LMJ2447epAJWzHTEIXbE1ODetGTXjp8K8wZirC0cZGIyjFwhOyB/E3
kerj/euztwMjMCBVPpO2vchlbs7frUiPy9HZRVh6lwn9Ny0ksWFMrWrWwaY0
TUfw0vtHIg7KdP1dXrVfoJnjqU5OvTiWDDnHTsoDH4GGnFm+qvGu0DJQOSQP
jHWimXhDweXJAI2bcEG754JN3ziJG7nf4H+zA+/nHyUKv8huGpyd1OzFOhVb
qoIvRiVInHIbGkSZLzW3AYxPK71Cv1aSbtLFcmsEUbJDI429ph07rCc99BAQ
5t2Izi3xKIv4E8Sl+K+ArFZ50j97yoJlR7kirj9VuPPSWTTDlm44F4Ijecx/
QS2T7mLBx9WxNJiQCqKcZrOutE9P3ez71wBeBIf92AIYsp2bubzVrGG2fzIT
CORuff0gzo2YFRHgXOAQ2zr/wV7RWN8o6ZhmLLdx8iz8ztdOV8wtpBiHAaUi
9XNVRsS86iY1DXMT7qIpNRZ8eBIRAjoCT17XjKEfuIaflL5Huv4Pml+YhNOs
qG6bWrHU7kGoRrTCenndx76FxZ36F0KNcW7fb6uxIhPFRXKhbc5TJRFZkAIq
Wge3xrLW3CVmnWX631VHlCk9LfVVF2D8+mC+VRAGr4e8H4WL4jLIiDQgpkVE
APwpXDj98cgW2LEd8QvCl8iBeCeAjHmkGZChzxJ3xbhh2K/uAkeZ7hJpaT2Q
PVHaKpww3WDRvk0zgTKhm/s9N9stDv2V5eTWy8WZZ6MSEtCFNC36u6bVhFEX
TEibM6dhMSxSUH7mapr9CwJnI5xaeQ+ENAM6EN+l/lwUv23b2OArFaK9fyoY
w5/xs5mBilT4jjqTFri9pxL74DNpOQf5TiEpk+/JeC/zBjZxNOezI5acTohu
rcwonUf1EVBVyagpv0++umEYMsKqPQtxFGSB4NiDPNfhFbSuABwWb43eGat3
xGiMrzVNzMRJ3+dQjnx7QkN9J4W9vVaOX6jj4wHVSmbqdHh+YWcaS592gwfi
LlrqX4P3/wqUjudKrsgv3mCq2wvwuWjNKutR0XiB4YMARzEms0S55BPSQh/+
w7DkaPWD++2PLeMUT1GPxRE8he+/aaRr5G6EYxUHhG6gbl8/NjUyy8XjSNCO
FAlAu5HzR0swB4Xno9PJZxzFIWASOKUi/AAIZ4Xy8Z3WZD844AWd3RYuJpDW
l1bl7HkI8F/deP8JLP0ZXE3jKyIiX8qyGyijhe+UDC65F7PhCBCgV4Albpmw
LUTpgmcGcvExPCmLukk8SAX60+GFFi9n6SLZpSoqJNKts8/rOYWdz+YL/F6P
fuxMIjhG53zlnD0K8GiRisb4/i5Ps2kmE4kH4p6Qofp6OgNaOoXEDaOB7z8e
9p8LfCLO8RsPgV1s0/q/72SvY0cv5C70YSq//pQGg2mWH9p4u4nRAFOsuwRm
L+7lsHkj6ROMfhk7XWmYFxplPc/embNc3FjW/Yiho9iVpHb52smgm5zVJQtp
Ke2qf9P3iCqGb2RwAM3Ok2Y0k442jWX0q8ASJkil26GV8ze86fGV0PKKNWmI
56olXF2Hbnb9LPof3aZtxgbTtF8Lu+kfWVmQrxmTU2lOCKxCgJrt3hC41N6r
l0HaUTOKUFyzdPQgdCIl0IjWzApMNDUW+R/hfFOIDBiiuwDZ6pJ43IkbfXnv
q9J9S8eLQ9tg7HHhB7hMqF2UwEgidOQXczWY1ON1yrFM2LN/dY/i1k/E9ei5
HdN4JX7YjVBuLYdqUs2vfdC8ctF5Ad2V0KOUI+DB13QESivEV8Cj4bmZ2wwy
s8Ll1KEAtLYzsd346lydiDc2t9eQLLojaowTnDHo0+NtppaVvf6PbnEj9GN9
OYHLpu2T8wb+HIJszbsCa3FiHc5Ayj4041Rfs58Sih63VhP36nJqstv60x4z
1OyAhj5PGk1GIbgmB3hB4ITITlBpid2qu0b3pLQ7Rt4Sjt11b2iQ8tMhn78L
5bUnlR3nF5RpoxDDWn9Ng0tNVPrcLw73iWkuYZPYfaSXe/HLlMye2k8osTB2
aqw0a+g9I481L0caMvSba+adsEZyBWH0QJs5V8dzWDBZOK8GiLIUkO5zcZIY
cBqcl2p91Vg+Sy0JWRUHf8XZTzKk5YG1BeQdrWYyJPb0+0gJJ0d1Ppy87/fh
oJFZ3uys3i/TNNu/RnvEu5Xr5PR3SWGxBw6MKdCgi1SSmrILTKIok2wYeB/3
Ibw0q9/gEM49lKJ2+mm9MyTRZ/MfGGT7JNgmTJYazMpNV+D8hpFlNKi64IdK
8OXuEu8roANDS8HOBYsoUrUTxxjglAFQeEKfTmaqTguBS2UVauKqG7+gRyYT
CCQMIin6L0W/KEInAOImccmApZLNFuuB/khR+9LdWIfIZil6alNfQk54pDiM
vHDcSBa5uCHgwlgrTD4SDRa6SBNaOfAmSBbuAhz/iwr9KdqT62oBPD5PtNhs
BRvab0E9tZkhhEYo87TDspLFOtMd4Y27RQcUGCoS+jiLmEHsBrrm/VnCxMMe
f3oVtKwfWP29C0QQy5Y/+1KBL5rlRIsJHzIdFt17qZxYao3/YV/Rmgb1BLc4
RRe3vLemx0aQix3Hpbm9ZE59IOad3Qsgsopr371wEZCJCBd7D7/gWYGHUib1
dfop2zReX5bAr7Smeorzp7juZiOVuAIO8hHk2okNc9Q+kU2w4LthMNUNQjtP
h09RdV12m5zTDytgimwvkhDSYmcVNI3+xv9IREbkI1jFf9uyr6wnDSG2atE1
tomsqkwgf4KJbgUwhSQRg22sCv++88bhf6dWEvk5csGjq604+bVZIZ6hiin6
PwvBI48WSbKHvIzao1LiH7KMpBP6hpUVb8R3hS0u8qCDBl/bJJ3d5HIv8kJV
feLX8VWeNrTltU2gDxfklh6Dy5XAIFNo4HF2YVFZraV008qldxXiH2cqFnFc
nSO/7BWCqMt0XJ/R0N1zvJZQn64A0uLsYtKjzEOJbX5Ho/OlMtINtssqFleb
xEhhIyhzfbT4xT1ZBwQ06fLLZi3FqjSwbTWNGPrqPKsDUfXpxwUf4a6lmB+F
uAET5I+ApZkdDrJIzmjmRoebF1Bcl3Hk/nOAIdFvAEOTGZ+hi46jdNL8uesz
G89fFnqD+23tsFd+3h0qIu3RXSRbSOmP9jNOtH/RZw4vkC1iGWwgWN0kU1xl
2vJbb7He/kCa4JYohTHgQyOLfmW0kVQIXB53naLa7Od/fyE20xMz5+i3yCGl
+KeI+8SIeUFsG7JUkqU34EPR0Hvlx7UC4oT7dAOt0vz3I8qVR2QGuwzyK0pP
i2/t6gHY0GZCJYYATAn5zcmIvKqfaC6EXUwj64x9FLGXp3RmTjztD70MHDZO
3wy54qk6UJJymGiddxC+GSaQ4KS/JD37K2hahps7KdGIAeiyMaofaVtgDyQM
0RCb1A2iOUV3pJpTFV86pJGUxWasau1kGmbTlcRXx6Z++TQaWrFMZ1sLKmlY
M5sjq5gm16jy3QzfEkwuDIAjj6mCULRW/l7LirWOqNlkplAiG+jBOLyUN4L8
cijRK7XtHQcTvGjKZyNveX4M+RKLcvX2TKHha6Hd9rSh8p/3Y/GiXZtdjy1H
/oRniNoHreOw3752BmqFRMgcttnuSJJ/W9VzmC5GhooDe1e4pIzLuCq6aWEC
QlZAE5KHlbPpEeuHsAB2CFbUBTsSYENsW+foTAaGHxCPAovMms99r3GsPIN2
vSwNwDk41SnsVgos0hHkFXIZx/HWdiYwPRoUQ8DeerE8PhPazqmmQuNZJLMH
4gM+QVjRWVjEhVAh9kjMnTE+jRMZlAuR3I7/jBI0OZqauMYbFOz2TJv9lkCv
VaBtsqBNGR6M6x8FgvHDaMwD4gmPkzF8FnTppP3QnB0FQcfiAGnoMPCAWJkx
l3bTdHHfTq0xtf4DLMYDco/4HMyP5NBk4FJdMESboWQyU3veZxOGLVfDTLWc
sqmuFylSiQCbEa71iAhukxigBL/4cnj0hamBZKGz3Pl24lGWB3AqY3j2UWYg
ca94pkLBetIpSObldLi8YEE/Yu0ugCqw90S9Pz054nJn/dKImxLsUZjDFIhm
hv5s3ys1cU2bXouAWWkxWS5YV6apVYk0/fkRUViAZbpcHUzCxLx6q64Mowgk
GpYWh33ZV9uyJ4EIqYYbiiIG0QMI0os9Xco0qIXevEBbqju6YaOEZz4DUPEA
9mtWvhkfctObW7kCLwStRdgm/n924/4Ho/ea4eTTaM7trsyVCCskpF1QImv+
9rK3svd2FAwVRhGjo8dArwctecvUMBAr99T5xur5NK0ZwuASwTSlEOgOvfd/
iELJtoIWA9uxfWVmuKcTOS1R6IFVMuoeBo390qgIqL25+D8m4usjEsHYYmXO
pRaUwGLBCJOxOjIR4OQbRrTYGllrQdNwViiPKtRDlIzk+6GG+T3FY293CZBP
U1dIMYlwPiOdOP+Hg5UqcijHhaEJ4Jm4tn9OL73PhEJljDJd4bAfSHAMC3gl
e224tDGD71H5hszppLpi+8EMiGHfJZoqStzQjtBxFj85NSYW99mK7eI4zANj
9SPYR9raSf7KXZrdVzOVs1kvHf0cJstOA27fmafb/YFCLw2TFWrKPnvB5OIS
/u7v0FyAZC9cdcJ4qm2arBmvIvXY2cYgO+87pdWkluWs8L4DP960vbC5MDST
hKsAqX4S7TfVoUxQ905dAyh6aE/4Q/yCnwU/k4fP0STzC1S8sIXnVjXP0ZlL
5bdPIxPExoPq5lesCMVpsF4XhghjdrI1QHpl2XdRloZhnnTSxhnqDRloKidf
2BoXmvvAIv8GDwgONgtER1CHOryv9B7vapWXzR0WG0S3AY39FJuDKVrOgigq
esZkPW2RoiNckqpuHP9+ObHeGWZqqPhUm7n6vBaTIzHqgZZOP/B35mUsMxK5
EoJ8ok2H9RsQXKE0XG4X4GpRs9oCaJfyPdDO0/TQlRkkjlJvXi679n5IgMoI
Iv8Q1GVFNyba6qUizeckZXSTtZQvGrCzHHgF2eh/E/MBkKooLZWM4tPcbnnC
xmu3WzHLL4H2v5paTRApfYR6fLdyiklXk+VxawATTHNuIBmdazfhlfeWa5l3
EnzDhH9grTPAdmZvngWREU22dZ9vYHkETXmF3VLeUe0QLJ4fgtZkxSqTvQsv
+MLo8dCfokkOe56rGAmz7QS53C7Mi+B+HsYWVjRzj0MRy4lT/Bb0/KNu81J6
aV97V75HJ1yb3x/BpzxrYK37QwRRBjNLAxlFPNk8i1UjOQ8B1tIt7qyIXc3j
J3zTgLG/iV65DSuv4wDYuOlZ1+L8WaH0T45t0lcd91NnH04M0LvZwVl8TTwt
81IG9rss5EUClRrhg6iks34mlGgBGqMNIb+1R54U4HiNJeO28q92TaBjdzcl
/frH1xxwcPUchOcjkT0hfET083wMcoA24LCyTyfwjpdp/0GBsFn9zYIyvqPO
Z/v/JgYhCn3QTFfyyZQJLfrvMZB4lB9FUnX3Hvg2ruUHntZDOMoaAoazI2O+
r0kZAfJhqgqJqy19pqJYOd+GjT8XURKPMNQTbJ7i+LHsp0peSkSjq6OmdcJ3
E28UB9VfKf3OWfeurC8pQPWuih9wRiKhFNKibmtg/pnt5iVgAFbQhiqWvwSA
RWYeZpEu8SxT6oIVuVnOIVPJjXl+GUTx+gNs2ocWUXcMPGZfbEv2I7PAHLrY
UtOfArHWn75XDkgHQ+aiXg4aLVOOuyeynCVjtMp8JWnEn4lBhOJGAR98vF4T
0v8TKz+z9lPxLeOXGUvJA05l4mDYeuaFQHBoeT28cB+k4PuHSplCDVdCWzDE
QRR/BHl6e8NnJNoeM9JfRvIkZnF1PihMYcxl5eYMjCL1NgY8Kqld5IQikHSX
9vgxcXGW3Fdkm454pD3E6GbkbkUYQRSBmsdzIFH6+r24m2Xo5JWYO96VVmc2
llISLAI0Rrtje1/+PIbfL4TuV51BTPb3XelV9/x01FcLjaRQwZ2/49FkfXOM
keVSAPODNscNufUV3MxyrWGo+Kgo10QKmLoHWX6cDc7DxoKDqKU+1szovOIw
7zTsS3y8K0cSprywF52qan6I5eOjTuCOWH8OLfTX3JYv6nz+CAxJ0WNs8Lq2
KJAP43kVmpu1o+CxdDX/Rqp8JbgPBThCVYOBgPnkzpSbGYlRdwPh+FPsbAZH
52TbO7VFpynNEPa3WMcj0p0ZpPZN71PXQpIuigNd6owv1CR4aiy1OEqYtV5E
JaVCquMriKjHvg3TTUkxL9SyxHtBzlHaIwapdiZNFw8zzjKXpM8Qsc5mB8QZ
gD/W+w640o/UN4sQDlMqyo8Rq3+U9y+JYrEo/ebgm9vsXl/WkfnG0VxUSMNx
IYqDlozEgMLz4EJ+vvRsICjK3dK1IV9jjEhNXV7ZIpV9niPq3iQ7py8CuKm4
Ii7SOU8xg4yX+ZtOhWdRG0S7o+4Xn2mehVa9/YJ4Ov+DLGqzns4ZBZJE8BMn
mQHaAEWuCzJjgBuQtyPSCR60AhQm0r0nMG8sZAm11i+Erz/cN9NxOISzsUut
o2YOjiriOZaffG0w+XfA3oBpXuKLWxVLule1LtmCc+QTWViraK5oJ31ZywT9
qkLGM5KE6wJWUpVflRMjCQuxMTThTwdP+/XO3EEi9PilZYQo1oklOSsdinzV
pf+HNI8WRn8u9MLmwi5Py7RTrPiIbPW6GSVPz9DoV/+icGY/92D8PML9ojr2
JKlF1QSjv1YHMpbe2/RZ32kPo6V+X6x+469R40Kmwe06ZXBBBaeMS0+I3Aoq
Jl6yrjNedIKEjvygo2S+pThEgvXsQlD9vcfHCMIvPjZf8WsXrEJXtZovR1lG
xqEY9o07u9vV/u9i7If124sXMxsCyueZTIvIosWzRJa+zlyz2ykZj/bHDhr8
bgRXl+EJhV0sJygT+mlzFL9ja1CLJa6Cq4lc8afInbxrcPMqdLc29Rayvs5l
vAa7ePPOE4RZTHbNUqJc4H2+5FXjPtWr2Xc+8rD62jzah2VUpZlpOJza3Bgl
65wtomSWhN2ztDAX2+iuKDs5IPcAmR7bht+xtaoFZeAbv70jIQ+ldjZBqcmh
spB/LCa5lBfKxq183ltcA0jNrZ+Y9fqpoLKfnQADrLs4LeO95eMmSm8/wiVF
/5MuEd2ChvKPbBgQGwy4jH7AZa3EnBfrY8DejNQSOR1MlGUit+n9KaJh1t4b
g3tZcNSbDXZufzSWTBdoJFOdbwCKh9YZPg+VureqQZNCL1A++cFEVBDA4etg
LU8T6gWHOX/POLn1t7KPyqY1q0Bdpx1mrDr6Dgh6kxiAgdAjglF5N2pE4XCe
OhxczVecopsd/Y7n1eT4fJ6XUu2f1IHYOkppW2Vi1bIjwOU4bh3zIZP63m0w
x+iuc4t3f3Rk9t+9D/bLJ8Pyix63T/rU4FGcFx8Y2OMbhCh/MsSVvVHhyK3K
uY5Y3+BB8ml09rMPllP0Z89hFtkKoqr5Ofq14w03o5C/Bespnzb+4PF9jxYX
PqvfzQ8D323UQ5DOLZdumqAdy31Mnx6K2Qosh72MXldOzz2RRFD2/C+uD/FH
kCpOeKghlpKHO++hqV0dHa0B2Q2597Ff1w0GHCRxFVHcEFlC9u/VGh+YMjPu
yqeU/q1pNqev4KiOoF+hFzrFts5puEvmOnltNKiw9k9ROG43OofOxbcJ8D3p
z8ST290lVF3iHrsF1kN6MFSZ7VJTvI+QgLzeI0gej+2ijYbTGZB22SQvq3Wi
TbPqfLAZO1zZx5TAF2Nr7i+Qi2GqzaM9v6d1Dj6e9awQpATN5dF9X89E6uf1
Dam25rYGlthm8uD5y3rDPm3y6xEWEoKu7/OeXWl6hY25hzC8KMeoFk8x6Jdu
VdHYw8OgVhbp3FglWmK6Ircsn5H44WUjEYVj6SAnnBJV5uiVLgO9PwsZ1cSG
JkDkgR2vLJCVTn7hWSe3cePhw/crpHw/Fl718RFMzoo1rGsyfGkkXzolUuNa
GhScF7v/fkJkJhsvNNswMnCiMbKPMmJ6zAGlCNsJxn3L4C4miWMwmgNC3lUs
V+boDNMRO/H+exXHWJmz3DQqh/6Ri33LOuI+jvPOFgUU96wFllBgNTIG+1w1
an4CfwSB+o2JsVG8dYFP4mt83blZnLRI1O7pMsyijbDVQVI1ITQGZGOj6gn+
LyJL5jPsHg50UI0LPDSHaOeVoGcH7XltjmSEU93Gu3Rjixzqyrgb08om+zzj
pnHmldpD4Ki7rGm8ERY0P684EjkpfT9X57oTe2fh/IvvCVuOKBpKWt7V+z7l
tQAm45Tp2hMWYbU+g37b5fEABm05H0NFx4vaDSX88QFSz741J5jnogc36qJt
bDb1WpCQdekwBngXtguwIkW1MsOfXMEWFIutaNWmv4zgLxglohQMyYPtHWmh
zaTFMVkWAAAvw0rD8Mg8059SmgKKV6q8dFRcuauiwWWLNgPS40opjF/pO0wB
uX6H5IIObWftHJl3L6/GICYohWRvM51v6cvC2l731YLWTo6lQNZC7WLI9g3Z
qkRY/vb2u8AwCXjwZQg3vCZ+HgOiRvyjM7QbH/77weLyCFM6oYd0ajtgTAOm
TPXe5DIYlhaVFSapm5G4gUdfLgnqgI16LIDGjBnvNXRznwSefa8Rqq3upIXb
4YPOx2NSzaTEhiOtisVsgjQj3Uq0gU8oZKsWeq66FqoiYSMFu302FH8EW894
QjrwZkpEkGp5ruRmVCn3Dj1Li/Nus8HgOmiVbS78coFJcfHNCOReic76WqfX
6pebl4rDrfDdYqPZ39r9lfIF4tzNYtAhQkqnl6tmAMjXzrcKg7tTxEC1lX/m
wVkBk1ACvRjdY8NIbjriHoMLMXelD58Jz3o4LmQn9cI2zZj+UYxDv5UwBAsP
KUst6DmSWzD7NXvbxyxrsofmHKpc9HumWMdZQqqmbEfBpmE4aoRF7gHxoogA
WEh22ktmjNuUCjgIJJCCe3fd/S9rH5JnzSeWvNDih8NPJy1cojDMPnDUdI7o
tI9Truj7gU3XPUjOWpyxBU2le9IJV4fOKqOHm04Y5UEGxWUPdMPVggqZUg/V
j69HR/SeF+UzDIUO8bK6e7TXoGQJqQE02xT9+mGrq6JSnNcOevo7SI/Ii/xG
r56X20jqSYlPl9lCbiwRtpBZpkDwAG7xiS+8jOGrAq34zEALu8JG9UZh/3gF
RWokZU4T28vmkpKkHtDdsGP0LZRI5Tfu/pwy7DiPIdCgOu/jZ+gkdK06zVtT
nBo0jHiXckjahbCmIuw33WETn90Hwqi7hV2aJQvQoMlyRUlE7BJnnvFp7nH1
f+WSQFP+pyFAULhLNt9zwrjVHmJERoCcYsN2WB8jhx7DyTH53ZR0odt2SRwz
HGl/fw53/TKRINcIZL6ZOqNis//Pibg3ydprH4NAPZJgvwjFNNMnMEKTpwqm
yC32oudzlz6ipRvmnOndu4kVcHawfBa7rI1dnSjfYwAnw5IiW66doOCdApYD
cIpTSK5LeiazLE2k2WGNpX+xhVLAaO/aPu0VoPSpPgHNzclblEn3Vt8pSYIs
uri80te49DTHkO7GoL1CQBhVSMDZgnfaWRbJ12KZfSfSHEoz591ss99aUex9
gO1rql/WX2OM3HK7LzpARUPX7E94PeE/16Ciugmmt+tE4b/byVlqwvdSLCYM
lgJuQ28hcQ+zJIn5yTkPDAV6y8h+jm+z8jJ4rOI2sY8wwMIob9QOSDdS6LjY
JmZTPJuVw2/2K1ImKkAQ/lxC4URqQNFyksfZNK26VQ/xC7RyiNHEBQqiBfTK
Kt3Y16wHWcLqZX7faWvPdjQ7ysY9wp8FWVeIG9oV92UFS0gRrad5wBqMUapI
e9HRa+dV9bmfr9fT7JuOcttL6a7oMcpQOuSTG2GzO5okqsbuJLra8asZU2I3
3JPOK2FZzy/sh6eGVoSxfIp5OdS2crM8U4Bp5nJmh1qRxheZJ4Q7MDxwy9yG
icbrMknfUqTSt2PNqJ9EiUN4H955W3qGJRS9mSbmkxep3K/PJ8VEg3XZFnfo
6vyVVJ4C3SpRKVjNwxwNmjs/tQUmQ1BK+Nev1Nm4WpVEwEHmd1ttwkxnDesR
X6DhpgiFbKV9+9yRtgQtZNDSPUBW9Iw15o3QQxt8cAf5sj4FmDfhIcxUNgsD
bCRqYNkgumGQTVqJubO+MmFfH9Bs1LMfK+IdXKgwDLwdSsGo3Ry80hZpEFHS
qRT6DCQX2VXlVovGf1DKumeUyv6edkbV9JWHAObQNJ290B9Wz2Tn1DLi/eaK
paKd3VDU6EbqGPnkK97l+H1gBeMLHAAZY/lOPR6B4kxWqZAW6huY+qhm/jlN
9xtM3xJydnDzVWoyB9Mqy8eQ9xSq4CNH0qRpasVRURbmGEJbL7c3WSF4OmAk
WTiu4wF1hZkjtUc3BRrn2ALccDaewBzGk+vGluPjTQNoJhJBNHsZprGGy18j
dp50Lsn3WZYuEVAdouZzPAPK/mXsHtEr5P3Rm01oP2WaDUywtcOzaewI2Azq
QLJTSjQKPZz0tFF2ZlrAJBMa6zgc5KLiA0D/prmXkq+cHsPAGgLrAo8Cfhwd
fH2Bs36PZDQaKxIuETaaaoelX7TNdHMAJVaIwylJfs5rfUB25yTY2uAj+KWB
x1AA8s6j/cXK6aNz4gdwJpO+kOK/jM5VBC/fW2FABeMAeZEwZJj2sXG3ABtu
5fEpQtqL4TykWqrIp8x7NGPmTpukZFmXIJjjEaV9n/Djim5P1cWIOKiZSqTi
wXCtfXd0yOW6v0FobosEORIaregOhP173+0n0pB1Suzss248N53kKT9bF7ub
KtgqxduyIsLxGTx9DHG9Y6dvZ5mS4yx2KV2YwVo0H4G3reHs1rqHUrP5+Z/C
6eUMZNBbqcCk8SircYK9SzBUhN52Vpdz5dGWRXKKfe6pIoe0WZCqgROrNjb1
RTUXpKID9KRFjbV/BP0WklxexcwB8ccf/qBSBLpcJUWqRIaYHUYTkCFCoAIl
O7CpZLawCl4fJQe/r+X8MgYTY8lbcWBOqsc9Qhys+XL9mcg4axoPugf5b3AG
us/2SV0aafac5iAWKuM1S/NKkhMq3s0ezg9utzg8S2/phB5KqahAc4b+zqMK
SUA/0PmG6tisUEiPQhuXZgIu2VExFrYxQm3yAI27ijkaU1qGnRcYSMISBWCI
Yvnx4hwsHVxH3uoMUt1v+KKBP6WHOvVa/jjot7aiB+Ul9WDyb1YQ7w1WfjPJ
kZXCi9gLNhERSkpbN6OL+21mAbmjdoxOddVR6QYen3y60eyKgkTCoSbQqKcD
mYFNn835q31tttEeFEVpLYFCQMe9q849Tm26DbwVrd/pGu7piaziZmsLzQZY
FGdpSMB5bScGGZbc3SyOTBJwDTIjsge4zfnw5Ly5LdHjX1reSme3GPlHEcYD
9nrlDtYUyay8MQR16QpLeXDqw0SzHFEkzVyHhkgBbgfDuWmQTqUqRyCaxLri
dQkO4bpMlFcw4XC7oeBel0w8jIFYrDCAjhIim10c9eReZ0DRxGHicN/7vPCK
zr3mSlLaHvoqMxihk5QIfSVrhJt94HlXxrPG6JbPC+YMM/XazAdIn1gxHdxW
hkcILCOEyQxtLH/12xICtbCV1HkrRpCZ0Ph/+0c+X92Kh2J4+fHVCZTg8++a
3LDN1ypZs3Uf2B6aOgdMdQGzdU3lnWVll5FKnptO3xpNn0v7fVTMiOqVD1Xn
2BEc3CJZlnp5/yxwP+6mjPrXBT9kzxSJhsQQrly3DfCaR/m4PSpFah1HnPPu
joDKNF85YrGq7wApcQFkq3oWZznr2RxtXuiUOp/Hgw7Xwjo86d6KhPVfLZp7
2h8i74ZNpWxBU7M27EaURMW66X4WNc1AGNV6QBLSNZyCI8onmIsrlMTifAKi
6Q+vGAq2fdL6FrI9CepWCk6nZpeKjBf/KlnLm8o7TkY6Jv01UIFOuHYHCEV9
60V9C+PRPNoXcfXyFjQVob2ceUZ0a6doUeD3Cp4mYf88+G5e0y75nNu5ekcY
xoD7/iFZV3QViLdQGWJb4mhjDozpbtXb7IUOVrKA47ipmHxlaQWbrxpNbOml
Vig2vUFGTBke1aqlcZfzTVI7G6MbSNmCHdHwvvcDSww9X41s1eJ1myA8GKIW
eXph+7qe3xplDptEmXVeQrM9btFTr+QkWPhaSQ1o/bsL/2a/tYCyh7mxG5xq
Pn5swOXzM/b/bJrJNR0Rk1fFCOgDo3BlpbXdNxrYvRzPloaA41RMmoehJhdC
tXAIMGZnmRB+ywV5PSUXcYKKpeciJXE0MTkoZo9HraUfJZhMGtBe0fEwG2qI
sSco25doYJbTgifo89xXxg59zfvsxT31SZWQwZ7OTe2RItMPM3KkA+0f9F03
ItQwkO2GkvJkhB9fG4MHUga5807GiyiopQIhTTDBJOJFQowqNU6+fE7XgC7c
5+W+sIPnXxnoUX1/C6U3V4ULR3ChcAhqY/bRkSXUW+U1QY6fAbhkxGjgFBY/
r5Y+1OdLlfdAMa7wjIMpCSzZEPwiRXD+6vdqlBL0YsZVyjkSd4dSfuEU9MCo
unBlensfpuKYka6NK8p2Jev2Qbt2yHjyoCgNXUBitLB/TxnZf9P6S6+d8Kcp
+yB+YSI8BiqXNPr+p1yA1CyWHFTfjNBMTCd96vrO+Na0IONMeCc2i6j0u/Kf
QidBxccdYXBcbSqyhT5ExZVIlKynKKvVUYIdoaeLdVEfso8V9NtDoOaaTS3n
IXIQYlyAe69wrxAJiIFP6P01Gf69FT6kQp8voNKtGWwuKBQ31b211sZkMtMm
vJf9ADf+2PjVfk1ReN7pl84m1w6yjrq9xCgN7qjeLCCjKUASSlEGOOS7sU5R
8pXRT0wsvcTEb1HhFWRxAj15pKxNA/o3PwfrYNo6V9TdEX/SLVO8zwVFlvZg
Mqdiq8qTJhfN0tu5j+ToFx8PdK5Fyd9VjOynSvrz/LH8ZkWo3dzxm7IFdo33
6/9nsorj0gF9I0+greOjQvEBUmW+fbWyzIba00GUyq9P30EqcN1/C3+LHmD6
/ucVMxD/JhChGnBNWkqpTTrcWVscn/5PW3gUNnn985FG50my5OxXbywem3gB
Ft7lkpqbhlR/DUtVLRGzsBbm4+kR7Grwl4PnKKfL2Vdw20bYre9G7P7+HWi4
Ln4WhaBrY8PgozRY7NwhR0QdYCoRuq9sBO9CZHhoMcEtiplDcr+leOtvEcFe
5Ye/8jUk6LtdDPHAMNp8MzoptMOLadryEPIocnF9Jf1oQnyQzepG5LJYUo4Y
0ai2b5KGFQ8ZQVqJHu2M8fib+lxgjJ2MHV8M2f5/4FYPsv6X9FoyK4JNeK2x
O2DvtPyQS+mjmbKInrwX0TnfqYsjxaWFPrqx4uTW1WLlU68bvt/kYGntZmj2
C6b9UqMtXadhso4nCAu2rOZjS7Z1nUWDDEDEjDH+qWo1j2L/hgmwBS+qd+gP
hLLD0BfDLw3EAQvavVKxASgW6YQuosiTCpxwUHlkgImFg6BPMxeHqFl4DXEe
7wqAHg7xmxSCttsxHtjTJWY4btAE83N2wPpfkP4nTA969GuhcRCqporytYMK
T+KbUbKV18Zg+CFVzG2FwM5HtxpxbZ4nwtVQOSWkQOT1GeicjpUsVFxacce+
JYApdRy1Afw7fPevTnZDcn3b24iIwWT1VNETwMmrfE3t26lRKnysBZw1vCok
yDEklbRr/nB5WrjDrSjdItEDVBgbgm8UEudsQsjIcVBf8vpxiWDXJ+tCZxIm
Erf0Kh+3OALZXxWehXzHVBX8IG8HY77NbGfOAbuW6R/7P76ioGVlZZGr6H9N
uiCKO/6qDpFmCTQMfR2ANYQWOI7RhPWkvQ4coNQ1WBIV042b/Rxjk//CLmbG
IkqWUeA14O14koPFE8K9dSZ+rxzpI5uLyqFpGahMvPH+IpfIjTjtitVJolRj
3mEDzd+rfodH8onx8R7rouM9PrPvB+UR4fBTcEfmivbcoNoj7XqEMo/eezLm
zn0bWJLzKJ3mM5pj8Oer3+be/X7ys7cU3yKvL7uGx2X4ErkON0em2o+jNz/v
fyaVaWk3bX80OevENIMuDu8sf+3QhilTAq3Yqa9MQqo8Em2c3gbGtPffvxgz
0Vcg2aI4WOMVEAD1NNHVxeUob3S19KmwCs0JCb605zB5C5kyU0ZCIlsUAV4H
jIsXvbqoYUtdvj4VMohtJhvSB03+Co0OlEKYRHF0VHRjKm/G3Tobtk/CYZGx
Jvf5iFZ9cfzEGTFNoV9nJSWHNowpsSOJgQdjemK40NeIkdvyFc86KO/Hu7ZY
rDg29RBXBciiQknYmsV0viyTvzaro0Fe9cT6SlwJ7DfOwALGpd/M54BHppnc
tp/YAPMzf2kcHV65G20n+/QiVOvTnuh3+vPiOg1V6wJeC1x54Ol4asGAFJUk
16iNhRP2qimn0L2GgwsWC7GrvaGfoF9pdIAl+rrRwJO+Dw1MQ7PCOuZH/M3m
pTJMRkA1rRUAgN4+PA7GjLEeFn8j5+loCZZF9nEnJkjFQlrFzTQnEe2xmRRv
nm/eRzNWeVfPENjCWlAWBhLyr7x/B7O51BI0ALv16k6jueqKYo3yEu1aqAaB
NhRh7XpgHleSRfTEG/oxX8Dowfpn2yNTduG1Ycv5NO6zwx1szEchZ0Bbt9uB
UAP0L00ZeW6Zqfuv5tvMhsWMN4wkH8x7hPVvyo1Yk7pUr8aDOk9zO8iG96VI
y1/u53ZsoCr+n+Hl/NPlucw0nm3WmJnQNIYl5f6W0ihs8Khh/rJkWDZBMxz5
g9zdiRPsvpt6cFFaNpfVpJ3tUHwHUDPLgsTPZ3GLWJW7rSNEKnkT5qLbgsLV
GahAljMW+PAN5FjNraor0Lz9TzcyXXpXyY+5Z/H7yXwf7mqmbPxHT+q2IWmD
xgqIsYtqEMDlgEdXqEL+Lua3FG5uiihgri4JfNvShV0D/TfUi8VhK1cuzTAG
29Cz96/e9/RDH94mv05KbexKUZ+Y/8rBNBmDR3CsesX3p33EDLNZTET8iuJ9
oYczjOJvVbS58DOVppyo4uESrpKw3hNj7JVJEis9fHZDaHmqEq2IgdYweUwX
rbkGdIEDex566DZlgJyVvem1FdPHQ2+X7mz7lpwrkBYyhsxFG0UfCxq4jRVG
xCQqn1/ltCwRrCkvz4gb7EYNhm8JoXK6AgwHpiuYwkVhCqQEy0yKKez6vdWo
9CsbANsURsgPOhJfTsMG/miWgEdACdIn3ZE8VwE7X/i8Qnb5eQ81QLZ1mpNE
HK9Y67pjGzB2Pf7lB+FBLoVhafzlL2Rng0fKIVtFI588Hp3/jH9rf6E1572h
v0CjmS6GH76cJ+RGbGZ8b5U/KIjlmcPDcvAOoH3DJ0RpfQzhLlVTPZJtQVwu
iBuxYE5N/opEyIsrhVtP9jeRVMDPL78eCgaGI9LPOY0oB9oX+IiJK+fLqj+y
R7BDDB4clxOycZ/C2G2zx+XGBoqXd+UT8S+sRHdOE1bmbNRuVMfuG8HPmgPd
PwYUZ4kDQYGlKL/qZ5atV8m/fLKAsYedfZPwECRCOevamaIsCUytCFCKDnOm
dqtNEBlG1EBobcDSFG42l0IzNtePfJpOXQuPwB0bB0drIBNLBhsXRtAQBWC/
tHcjvhSUzRjQlSshOdpgG6t2P5NvfVcWbRkNP2NkZ5caXxCLNTPPzcFG++jF
+E/j4iGmzwfZKnbnnhMhBKjh9oVGEgPXJlYFuFL6HcHmwj+r2kRKZBsq1YTg
FULFTKYnNMvWolPMbglRNGfkk14Dx3klu/wWCI+qIKUJIZxeXCBiJh7bPqek
ni8z1D/oEvAQAFvp0yV4Gx1DG8Zo0hh/PWaNcASBgZ8mk/pIByIHb12Bxsbb
thfEirqGpr0fEYgCAiMrw8h7J4DuMKD/S1h4hbvyFPxwwJos9OS+Oa0dCTh1
0hbd5+r35Z3SsZJq3IpfspKl6QZTa3qRjrnFyUjHhM1jB6DWH+nIu+rXNITq
ZwixKcxqiXS+uGKlaUbGQVmTzipBSo2l9wXy7Qz08ZsVhg6o/SVg05eZvg0S
j26M7t6S7se+M6m94vUcqjtc5O67GmhG51YB/7z7rvkOsDCsYjpcTDIYjOC9
UYO9vb9Mpr6iyWvEj/rEZCNmmYUGl1cPK3MtizYIa25kGtZjVUXH6oMBxE0b
d5WHCMht19RvkevTRAy/0dYOEMdSpPenKeaCYk0A2ONxpq5YQ5rj9aM0mwOP
6BDU+2qnrkQcf5wuctBSLvhC8fnAHIoSWG9Qaw81R07GrQN3Y42Uxzi/EtOD
S6RImufSAnd9p6ifr0zB1GnVU0D32pmxhEUwb6DbVbWgBipfw6KV8ADV7eDs
9Rd2IryZ3cUuyTzYXvUNskusbbHvcvNAgbnJLpfYYjwBJJ+QoZQjFB7mP071
gfooWo0vH9vgvgPPCmotcjXivXYeRc7NWV2wg207wSkrUl1rYFyKYJd1hVC5
ZA83fcx6M4StX4garTnku2gbJ7oXlg8VBQzlLofsicD/3jXzZzSBcj9Xn1Mi
m5+xBUDY0vxzkgy7JAuVUDDWpA+yDzMxFH6map6HS9NAP9S+2pziGg7QF7ik
2VF4qSESMuxg1nxk9e0RKosbnrUtQXAaqPz32ig191BjrvGSFz+XBugFcapH
g4ySQrqMfvJrG2b1YmsuNYcOn1o/fiW3/k/fdVVD9pSqNexCDqqgnyQypCWA
ogdaa5Xy94Q1MWooARSHTvvluGgLKqelx0bOcPmb4mLwDwUHiA1na2uTWefm
BW6Nzg2VcN5NmFmR0wmIW2VaLglNk0z05yaBtsYIc30CoRlwzFp+DPeSUR3h
edL8QjeU0ThaBY7CaJ9uBZmHzds21OGeWIqHlxGCunxWjdd9gb3Zx3DlcjlZ
Zr3F9nq0+Pl3MPV48KvMuTJXSCkB71deBjWkrWuRwHTUZig3soPZNBRg56bt
PNL2cT4NShcIbsNbFUi0Gvw+Ke8k7QPSflyqv1FA4x/3ArXWu5Pb+4QQKBgI
gmUaC+DKEHB1Ok20XWnGze4S+A3L8VaNGOcpetMn0bjLaTbuq4BzgYW8UmVV
YAeCEHSzIw19w0tZ98AWdjCHHkFPfjJUSuG+5yAnV6P9mOMkh4A/imkuPC+C
hQSMmsgJAxBAiBZaxUTMgKGIlTkVi0+QgWOa3GF4MKq4ac36BnpTRxQxozLk
uQiVXM5Z5htfkTNr8reWwoHodqMXOwiP6bNLYPZCW+N4lD2bZdSVOYxr/8QN
B4ua14fpMMQKJMy01xfMfClxBY9iOk6fYCPbYY5KY+MQ5cBQn+9JbEZt0K5e
9h27lAsqeXfwMFJiV8gppz9AwlhVW5aHr2TlpsK9GyLYchkyHXlWuguM6bEq
1J76uhbY41W7qsaUBEOhDA9LPv6yjLLsxz1SQM5CHpzrDIor/sboXQRWxncR
oB9TGpDudRDalwjjXIB5UdNZ9/TSViIevaA9c+JSdc3y/NzWINHa+NKzqtcp
kParwmu5ljiNG9PSWgi/XLS/r0Y8Txd4fn4nCO6kdsaVywVg/m2UCciZsMvA
Cya/SXGqPobHXHrY8njTtqgVbnikZI72bslw5x0HHTZuoYu8LAXKygz7pC3W
Df7Lvj97wqynSAT1fxxUTA1yCtkowp6gcQlHSGux8ikSOn7hkNHEWoP4gqbX
4gkCoIiaptMOQVAJcX2rJj2JHAuhHIw3h/z/YX9Vy2miRZBMHrrbFI17Vz3v
ST/CZdcDx0HpaxoJOJpviyuOG3SF70JxBOIdZ5sB8LUpqr0YyScWi/Bm7yGf
YSaCUvhGjzp0UlI/6ZbHR+7V0t8oToGs/FHZboLDV17Ook/FolWb2W4nsSiQ
MN25AWOXeMhhtjnJN1I0ttTB+5YeZklCddtm8zeXmVoZrQtPHizDTrc55rOA
vyn4ONpPc2c0vu2an6KAVgMd8T+OKL5OI/b7gmIAobcHmsU1CPqxCtAamphM
EbY80/Km1goI4YEPlG6ynzuxIbsbHIrp6cdZjDXqXH4SmcbVU/0j2jdU43+7
IH+r7jrurDGJ47zUYPJNdCYUe5qY7U7jEuKORBC9hd6sfrppqd+aTANsdktn
h83r5JxNcqyn2kpGMCYZSxAGi3nfYLkxCBTZfmpFXHwswq6MCp2KDbFDgR9r
ioRCPvFD4zSsxz2UgQ26DtXb9IyoYRFgxA5xsDqOSL+mB7TfslC4i7OXgkTt
05Sr2Mc8j3fTCjQTXxQ3H8MDHi3kGVzDtS87UbCVpyb8KrqFBJBOEiLfgpwz
lyjd4oevV1rQttUWYSdR0SUWMtanb4U6At3VSfxqdf25l8eiXrEgaA14FIAU
49vqMldwYSa+On4cSiD/jengXuR++z9cJQRF2xl+lKb88w2G4v6VxF9DN/vV
MzlRDIwQTKuA3FG5bet/V1LiQPF7RqC15iSTYhsn3QUXDFtR6UHhPMcsRv0D
hRXAkCt2kdAYtQe84yx2v4OFEK4A3i095ufmo+Qh/ZbyPwOBhVMilvEXCIum
xVSzOUFHwtADNFfx4ac8w87pqZo1iiOAB9OFwGGu3ffeOXOFLU723J9hjPGn
alzCWEH76d3ogrDpcBQLkZgVEaYM9Kg9qRmQuMYKNzCcUa0XmwuTXS0DDz3W
N9SL+CjCnpOgKi1DEBCmVVjI94/QWAnrr8m9IA/SU2089xHYn35xSF1JA7JG
+S2gLUiYn3nmJYXGxKXVxBaOcC/aDZ9rE/AAJsEwPyFpaEq36Py4j2OEhClu
VbpVrwX8/OIkJ143Wmu1TJV97tB8TwS7eHyBqM1Le3K3xv0QNd2MJubjvS7V
tJapBoDrkFRPw19XVaeEwDzGl/AYmMpVra0KjEdSjzhVUaTFRj5+DCwb04uO
pfYLNR+BWjkQPLoUdc+46nlmFiMvV34ftXZEIq4kJzZOSZTYHQ6OXn0q74FG
Xdktm7iJKMRV4wySNsVy1W3hHjxGJhXlyxCArfGN7SLDTf0AZC1XnPRlc7bw
DiEHPng98+Q1KEJNJqqsKTpOUoV2oWPOvBM6KivKxEfzPZ/t6UcXqC0AQZUu
ruIarfPwqiR1yN3+Uj88R8qvWZ7qntjx22Hglmv30RoMboPcKhNn0b7XBup9
7ym2oeXsIaNUrj4+JDIPDn42Im+HDfpbp1Dhl9c0GnA2zHuByLqtvDSbK8SC
Eyy4/5k7HJWJoOwoELgevSXSHwUlXCSphz4XLjqhjz2p0ozHNvAyMR+1WrGS
pZP5u3AT2v8+lUpATIAGfFLpboTacU3pJNM4Yx78SnshjgzJNck/9YmwXpkR
fVPZFhpD+E/WUenrYYKaxbgqNtc9mdcLUQa5834fwA7MvfBMzFDDXbdvpcBM
7AMB8X3SdBUKcBCB/9JMpMFp0mCr/9otumaxVzVQxmrZIhyDWWUwIM6h7mt3
mxn3c5WNaH1WK+uVUiedtXF+IxB9NbTVvrIvNSdv2BpuLANxrJBug6ldb3CW
02uQmOxYRRkj6Tpz53gL0zeRn+PJh0VJ1Nj1ykk1WS/tw8kL4XTPL+hPPHJ4
A6rWbS4WZWYjwypZZWXLZ4d1Z7bhdtg5hcAv/qSGQvR/myvpCjjbj9wK4AK8
OIpq9xX7zQ7gE0guvble5C4tjsPvhALCt9/sXC3UI173WafeSDMxSxHN7rLM
AqZPpkBmhqcMKHf/QhNwQVr7tNIS9g0QzZOCPBgCYrUzWqMbtjYdA9OzMYPY
rWCZ9LzYbkFjkTQjeGJ6aQ+iYyxs0y49RzdMmPWO3TvVov1idmWpKzykXepN
8iyTZfDMDWm3Ct5jUe2ai5PonsOEcck4o38yznNK5GQZDtjr6qSRUkw1bbiR
bOvxVM920N7ZJGy3KhWYesGB0APl5EbwprbNuhZPfy17KzZixlP/fM9xo3bs
eo2qlHQDaDAciKsJcvzqxngOHKHBLA0sagAjvMItiBVKnJsxTjUSUajTaydb
oX34++DoHgnNzpIwJKFzQct0XV83Uim1apNM+tRYYwe5dl7c+E07ai+hNQjI
Wn90rCqVBaABvRiuEHdG05vUgvixcKKWlJ4y0QzVw773YDhTx0wPo1Gcfnk/
GoRzuUsgNHgD+CZBZiqhKw+gT2dmNcTSzf6SHQ7s+eDsiqUdtUdCTlJAd89X
ESlxuZ0vtjXViM8n9/8bhrY8xEpvjhLx4mFhMqceOIY7cRJQiimKOTKIL6e3
sNvJKzjfT2X4XG8dicxEz5FqacxCItftbKB1DxOzp1hVieOO0rUrGznqox4o
JYKRSiiwcWBs5VyRAbdOBZR62OXOTFbF2HqQlIBRIe8/6WHk6IGq2XnsdrT0
QfOkDm8fkLVJG21dDJPbxbd0euIlJmcegtZeHVKN4dcKdMJgoUwCLtFOtnGh
Ko4NyHcvwLNHMeCnRfCSDba7nsHfVV4sQzdnw2rHtZT/K3ql5wVILVv8itNN
5Cqd5r6Ef6IU9rjoF0J32q6dIDFLhqxanRoAO9zVxzX6XD5kim6sRfmI0wrZ
NeCtkrY6UXLyGn1oLh9ig873rFMavjfK+Ukm6l0xxUXISOzVYV97tGFM0awX
uEmvuKZB/DGLqqRMdsM8eUk9UiqFIA4peSzaRQ4jBOC/iPGRu8hUGxdQM2bD
u+Ml6RbeRWOnhP4V+rvg0iLe29wQKZBqAMbG2gn4/SU1xLPpj8QSc/Fb6Spc
1Odg5obMTD/0a4afGgPPbpgd7cK4T2Av5eByAMp/Po1IyVQOTpcrJ2GOzFfT
gEOCl1hHc1Pwp2wnRRTRhHmKoKNsLPmmO7oM3eG2bXhuLZuu3XdODnMxgU9M
x1sN6KJMXK0371PjwiI5uK/ROBzCxsftFZx/iJIBcO2FUa8sQqq6px32qPKb
SEc0wpywTNdGCeZ7xQDMBsO4ig4XEqtPPqo6nBLHwwd2N7GdYKcznux2O5Xr
bQqGnCyWKJ5ZmJn8besjbaWDwVUv+nbB5SRI7SjMIxMBuzWKaV0AjtsreKB8
Jii18Jd4sQkeczx+nkQgChNKJOAdshMeLcE/9FiASj/psm115AQ2s+P/8cDd
auhqBEBIhiQpnqYoRIN6vST8jYYbrK3ye34v268O8h2IGdpAxEmvMGQ1crNB
zLY2qk2PLMN83V1lD5pHPIDajqabQByTTveW2EYGKX39qhb+3uN72OiSlQco
c2E+GLdw1PLdUUOHIxjEO1X9tGDh/olVcEsaiPh1FIVV3ikGUUTMNHS8ZgJ5
4QVfQAP68xMWQGQspoZkJraKO4IRlDBzjiYA6VTEAYYeMrG6KJodqAzvvNOH
N5rDrDA8MoH4mQeVlB7NqnmH5Y65PB5Z9gBtFL5VIbGCFwjLcixGMTm0euS0
pw0rmolfT3beZZXuvOThX3+qZqxwPy8luW51EG8ZwoOnNM2PU7P2cNgTg2Kp
iaagbanYrN1NMNZjIEU7pDkygxyzCM21Md7pkQPczO0JqbeMKCSTPmhgIw4I
UOozMTvf9f562E73xd64DehtMg1sfsWvrdbGZvZIis6N+g/VRImTzHHNxAYP
8Is0xiP/FX8iSff/rBtvoy9ljFCX3sXalGOCmVAy2rhRXHTqOl/I4Ie0ryy5
L4mG1Wa5/3C6nVAhF6cMDhYStBO67gYVlu7ujIqQZeWEWq6vom9YaMHkrui5
rsEHW/TRwl6oOgVSKS1bP0uOKgSLGtDA99jFZQjNi0EbCqtBf2JRKi11AuOS
IVmoQSCXh2+GD7fDN30jfnEXFHPug7y7+yzF+0rkHogUaTb6tJwS8JzwgRAr
8cNlMrde4AqvDk/8OLg6GtXyg0ZeJLn0rZpT0SBEwiptGEq0J0LNTLSq8P/P
+NZgtqmhr36rnjSEJuPthPptUgxdwZGMh2rJ9ECcgjX/xC3ypk4HI4LqtBX4
g2Kn3Qdf8m80pmMadhp0cx2u/SxWqYgCA6oH+JuLp4CFLyCB/QhIBn9QFKhH
x0lvyIzkhNXqA+kE2p6ZeI7fhszSFDGicao73uyKeTln8y8vJONJDMfiRnFN
mh3fd9a95Wj9h/sd7NA/j28tk0DESqG4MHt1lJsuh3DSl5YAed0IiB3EhzeD
vwvGCmyIz9OMapV2cJ1N68QsDRL8LKF7npXFaP0Aj+MxHOC5hiLyEAFKSwQY
J2Oe3wRliv3BH7W+n9AhukMLMLFYTpdjpcVT7lzFg8Jn0OBQBKd10dsMAhCk
+/BxwRpnugj8L7KOsZ8yeu8i0heZUuh/5A102jiHF9fVheH6jpx7gGo8jj3d
wo/IW7lDqEOuZCTaROoPUgVNnRElv+9setF4QMKImcknbbitvaGr4sGLM3Oz
54ywWvsXSYlof80Y7GXSNrJFMuPg5o7k/eRMFZcXuKWXhyT6y6Zo5pBuOqyk
65eBmrWs6i13ir8r0zRisMlse58BHXOj/cUUAD6ukBNg+VyFRuTORFmquT9g
m/eWlhpwFFX14v/RRKGnE8nBcdqZFuwjZswAvZrzKuDuFJpSQpjlQR2wIrRX
67iyijt5HYxo3zSzcITVfo4agcrLC4xpruau1yYbhc+ZoU7XUKF/DR2s4BCL
+UPcVUPp3tXQLjnFozjBLVKXqRdC7AeozBWuUBGWBtXhUBDo0L/LAwuMqvsg
tDvXqYBZFLdq3zofiyymH0s6Ayo6PTyjBxCC6eZqhg6UrKInIk2YBiTi2q7+
1zaQ1DVU+Me6/WLO3ZkQWblb4nDX3BXvxtsYZ3ssDyHNyTvCNS48PAVo5kbp
I0SCF4pNkYUNf0hoZvG5mlvZs5XWy2ZHsmCRkQCmq97G2FDCeMXb/p/nLaI/
c32f1x0a2GbhSLQ3vX4je1Z79vDtBUbgpTyMGnL0Hj/9XtAkpLs9a9ej489J
5BQNXOyd3JO1ARN7KdiHQeOV6cIYwc9J8W+tD10hVEFcyBaEBhAwoOJkWeM+
fZZyJFmq96MCW4yIAGtk3WFatkts8Y/JFxzTUWR1ziy2Q7Oiq5cbT74SqaeM
KrmAREfqGY8twnBleQDpWAYqyDO3zPdrarkHZeMbGdkR+SxAK1RLKMxwFZBU
JyQPhuChp4yK5IDns9meCIcsfiz7RjfvzMRKCYVhZRfpr/xBnXors5tF3Blk
357iFQ+N3zZGu+YhoYLPfbcFlfd4hlU2DwUzEGd+7MDdQS1shD9c6DyS2Yg5
TVFnt90TbhUNQoGC5OKLrTVEWjN5H6PjwiKsUi9Aeb+TsV6vuGGU4a0L2wQX
5k/tzECWgsqsiBNfShs+b2/v99TJJ34BbZwOAG0xa+qp5KJGvq9EDRQEcdfg
jBNHJ4t/VWeg3WCnwy1IHCCDqi0hsk8WF9b+3fvhrxY9hZG+kma9RX7V9AuK
Nwv8nQtoSK9CZb1MLSMJtjB1KLQIKSZeuglfjQmRpo4G/oE7NTH3PajKt/ss
JsLfCqgcPMkZYrlezeBBcCb/Tjt7GSHMhoP/9hJK+JN+89AwyFrSW/3hmu5t
OrfPOsIgE4aBDtD6cftBZzWDWiFD3/Fo8nqSJNmnCFF4EhxQpEnUAXvhvOnC
i8xMFCgf3s8lYEApAmolKb5RmrmW7/XS7Xpf/B53Df2JPzU12psd7WoOeYpA
sypU4JgDqV2rOKBkmBWEMxLFNYKj9LHNed9pY07+FEf9suxtdOA3dvuNXxmx
cWmz2uBgeQIO4QXt9UeFpT3pgeEudRYjGwHmDxBSa+eGfM3ZHxs3d0DqjXYy
9fFrtnlgSi8w9UUYfPYsp5XCXRezYXFK6u9zDVLmPHvIDBkkb/Z67Q+IQ+ob
2R22a2Wm5g9S2hUGuIU8o+Zqf5SHk4NW3MleuMY2VgOvCedqqaeFWaBFRtXW
NJwgBS9pFuA1QZfSPc66zmfMcg9+Ago1hTaSq5wTbpCqu6MR94sK/wHgyhpH
yOlmoIldu04IuLJAWyrgtdbrpVXJK+Y7/jaz5cdaW4k32YolsN7Ow5L6/a/6
BXaJaPbAMYjfDaLEhhD4O+rF3QW2A8eAc8tOSponkdyH8BkmmiOauRwDuDkT
QMDBC7moAwXuGS7x3NZAYkkQ2yyfPlYJ9VF9wtMjcEM1v7LMmY5wiEx4304B
MTXaZ5h1j5ENIhS5hs+M++RZtFtRNxevvZB4ccFatTTC6/d4FJp8L7gAD3hd
8nJKfCBz6s+ovKUPucBtvYFZChibfnjKR3Y6yRPYfJpGXYdEXw+pZSOSGqEV
24Z8uvv9xmbmkNaPbd9wxR47eqvjLE3G+bUUlUOxdJv+JNHwtHDtR0Bo9XBo
9tdtL5Ar5Qcn/lYolPHUgyS+yHLwuSyf5wWM4C3Po702nxjB/jmoGsnN/YEM
a/c1krV/4bO5n8KCJv5Sl0oPOEInCA9HVz8L4MGQpVCjrBo4hVJuuY4kPxxv
j8Lnagnh+q/hcjPfEoKkf+4V9fPZtl2zO74ZYpo+vTXBK+YKEKKbw19mmauZ
FZSiz3JI1G+mvFhvOgqI5OnXaZnApi0dMSuLLCUfwQLWsXP22XVpcVdrcwTC
aAShLKgTfFxLQFTKrtKxf4J4MHj8UOxlvUFZf/J/rHQWdKQB5SFIL2jjkDEd
F7VkL4xLV56Aq95Zr2iupM6YBTyIn/6JQPtvhFb+NtZc9uieqP4VLc/RhZ1v
Y/SE9daM8TNmF+lKPQ/40QtNev5201xvb9YzzoHNJCoaaIN/K0InzsYJRt7w
IGAZQOcq6mvTA9tIIyAdobvyA92zJQpMz6e8GTcesjg/Aeota2rmpUzXQrv0
JFou6kGibJTVMFizSl+6KrI+6JRshXmTJ7qMU+vIasC/zVupgKonupkjKGqg
rYhsmlibhWLEP91YqKNJVePvYqwaamAuUX7BcXGLQbpw7QooXc+igCjB9cTH
1Ed32HOdaLBEft0lKSRsJ+5sRK4bfWakmUY7nsyPrTfTcd2qez1ufsR1WUfv
+ilkHVCKub7VKmsIbkkQyC+Yf7qgXViepeCHxlIViiMR4VJZ+2zrW7JULOp7
AU/XEKW2v5/VVaYNaquB8CMU8F/1d1kyteZx47DFqYNTNipxrnX6fsUu6d6K
CgYv03mmTdKBGoHcdLb+v0fSo70bCIuraeDK8rUEqXFn2tyFt8sQu2f+J4LG
e0au2gNbgH9WkVJZn6TyI3NwAeR3LEVCoDzzqOQBmpCs+DVCAB5/izR7fSmw
kCglCO518R0Vb+7tidpJUfzo0SqH8piBl5u7goe5HDepzZkn4rjFocnRJN5C
twSqFowJBBO8rfuWx0G1qCEasT/HRg6H7BrrUEucbbGTlOuAT5VjSImw15kr
kwLjMwGgPEHdQbFSUPNElTH4DLBrBf2NuZW8Pz8PYmiisIk1axorAd5bNR+U
OIeNbz03ixs9cI1p3hnLp7hx2Dm0Uzsi3iNGbe8s6qmVCAgjJbihCSkK3zaQ
mQgEGSJKE3H6Buh54a45Jepf/Xy2aq3sVpYq0iSkEMF14KzsYzipO/8r6kot
l973oPlHPOn7GQjcBdMq2ozn3T4oft1EBP1nMd4zE9YHcFpi6co7V8ZQHkn0
vMc3+c9m5AUIIn1Sl0rum8/HNojt5RVk3LQ/C7kXQuJ70hq28JYJgp15nj70
jOikssCSI3EaNVG4uIjssgNv36xgDRNNdg7iPrAGfxnKZz7A3/yiVrL7iTRh
hHmFzklN268StWGYoOBdFC59FA79Z/VwcHII9K6wgQ4vAs0kMDMbTmgJd6ef
4shufSjX+y9uocWj0MYK5fA8fCUEPo34KWZQJ2+Axm848diL+QfEx8RfCOKv
Fia+Vg0er55/SB9n807XEv9SuNh+X3Yaejrw6CCaQrF9KivBcdtFYeL3JUiB
RnKDvOQlykRgSmrs+PLJb2NjJKCQZM8q13VDya7DpsDVImiJjsY9RpnJKG9R
qnGaxlGU5lW6rnQUikG5x1J5umezIYCICIESmsSDbcyL0nt0CFMpYEoLLC0i
wzNqVEC9LaMDtw7gkRmnAclIH+K/NWWyUIl4I6vIwUCgM424PAcozvdkXL33
E/EF7DTapk1txsauZGzk1h9XcBrfx7bJtWkqGgJuyQe5+53pdkkOA7QlCg9l
IH8abFk+CAErg63IZzG1eZ+YyFFOHoZt3m1HfV3XynDv6UGUZ9sI1HApNjOg
yedRhHnQFmh3R8mlIKrc31Tms7GSFV9bpxZTOf0UvGZngd/FOcKIqmbRg0OM
9fnV9u5IvBj61ymsWINL0hAV0Yn4DK/2x1xcWyzat744B02Uja34F9SsGS9o
P/NclA/SIMHhoWWztq2LFXIdyqtINonJadUb6GkrTnQ7THxP6BtTb95zjTag
LQqQ3iS1RsDzk8Bgn/SGjYinjAI58l20c27kVlULl92BCi48A3gfIMI4eT+f
E9Ag0BmLz5GXzCtn5Wj/nv6FzZRbYPBLudQEsPHoWUq0DA1saqnd+DS4Peoe
G+UVWUsIHTOdIKMm2S4GNS1cjLCNQGguiYXO632ckXcB4q8Gl+lR0S6RP4BD
2H/NWltzFJmvR/OL8VP7xzGiKv9JtnvXtHbUAnqLc5kTN9R78rntIQVfSq0s
9UXl9na1B+B1ScMLhCINCC6sohLqhL9ktGkrooqmc72/ibWOKvq1SJwIRTuF
6cHBmbpx92H2opQPt7BFMvdzaz1WghgN724KohO/aS0H1oPd+vliBj4JgJDN
tNyQaXntcZnUIcb1AdOLCaqrDeSVDhSz/iM9h8FBzwWCP71rUuYf1hcEiTWR
NeZxWY5RQxhdHEaaTK5uok5d19NvaEBepGYdtvwexOkw3oKMgkjAYKFr95cB
Y/WTv00yDsQZvqo687L727z7NQ7somYHU/N/ePNm+cl7ael2Qj8Px4qhS+bp
RE8Z2EK5ddiemoN02R3ErMEQvEmsTlpMaNn5hnGZo5+RudUxmWcsdsEdqiyq
hLG35DJhUOOfmranUsxwL8YiWGsF6QyY4FiOqhYJ6jIr2TK7juWlt6dBMIRs
taXwWR6thtq569CohrSGV1EujhMzCAfvXONS5rkxF/FGAzyGFz0f93I9Ap2P
d+po18ylCDYfqJ6x8p7NkcDBAFdwXcsQp+yW3kFD+dMFNAoAG77XJEOb0nit
ovBguMwLvnwy1z+spmUF7/VO4YqCQwe8U2hzuKGOLcJC1h1DhCmeOb+lYnU0
AtpOh5Kb8Tlu/C6eNCmJ2DHfsESPrT4PS/WAqGo6q6VAQ3b/WUj+8kvneMch
6349MzS1Zo9PT9sAXJSXYOGTtkZe8ga2taAZ+rzpebmKQ6RhY5c4pQUU2hSK
Kxe7PWHCIyXMuCaC4sMbprXNEPZXuKF3b9/4KEoPAhyqpZfaKWHPlfYVW9x7
I9a4FPOZe1W/7DQ4KzaCEpfZcxMNpF1Si1KeSINA29ImkTlPM65jG3RMPKeA
MYiosESC5StgHLMEGi0zosDTqRW5LBOahZIBYwi0Gjyg47WNdkX1Uhx5Dzjl
GKsM2Vp2vUrBGzL4jwHauWC1yTGt23JymtgdcpbZDQMIDpFaUdIzU1u+pqds
BUmWpcb5O4Z28Ps2NIjHTBG7aQ3NGpHbJW81GM9X1zAWdaoq9S9Y2zbuRI70
7WTAJYuoL4acCO7Y1CQiZ68W+rOtARsCOsH3jJ+69uX6wfqbIpWB498eL2DN
08Yl8CV5Jk9ca0yYFGcosVba2syFbd0tHU1CfVPqDJRrYJH6GOfxtZ4QTXAS
jVfoz5fMgI/wkWBLYeMOaQWfFc6/p/3kRCNh73+/J7PhAnFTu6hDULHa/8Tw
YfY9WzHbaREFIIwtghg4GHDEtd8O43NKp2zpvfmQA+DJP69XWmvuu0G8cXsb
oghDLD8cLtFLN/D+IrgXYZ4ZLxCl+prRRtNghiPK6PTzLzVwtDQPCL+H9EhU
/FQbrIuQcGRPqtjtUFtMsI+EDNvgFy/kbK1bysztBt/FZAle/EoIrMIRxx53
U9Yt4GjSrQnhP6sq19HmVPtnpexTaUJqqgWY9FkajyOhf6/G8eivWb/C0rMz
V3PZ7u7C4KTFURzsPqFv+algvTbCz6RJbfKnXEX4XIF3ueiJznPoURiigvrD
knV4/c5EeA3sRsrLO7ORrXnVf1YDwCKUBKlKClOEITR7hFIJM00fCC+5YKdw
n/x2Iz+0dbYkDls4vz4t/TDhP0n8ReFnQv5LrTlsHaGDGAjMH4Ozeldp241w
kaaTRYcDA54dJD/jDZP0OyS3/SFGanp5xH7yoOlKhRCXA+8iEl1o2+WyM0EI
eu35tBYJJMd3zwJDfTVyU8pW3EX9mUR6laLQe8jSABWbFqZml7SecUinBOWn
5QOWdiuc9WFYeCJzN3SU8AQdrVWKOpxa8ITFqBXxyTaZk0prgf0efTyXnkPB
iW+47Z2FN4iLlQt9YAGavtGbrQhGvqrX6ImMjIR+sGN84RZcw0BCrRCY5N/c
q+yTga+8RBInoxBqzbMnQpOkTC7kgA8sy2/fjYXzm08FuXhylrekbf/V4r2J
rMYIwVpmJ86oPzP5lqCE9pjswgAbF9OOmqRVeajtGnOp+kbqXfTmdHIWDeEM
Q7NkgcfaQjJawbtVKYGySuvDXDb8aKwYcaX7YOTB6nRptqdfVh4H+sB7dqF6
dsMcwvMyr5BHxgwdgvpuLASqLvCWn/R1JQbhSxXgdZO2mV6Ss2BEn0yPpTKa
dRfnaRVveSkdFqZyZMERQhosLvK9Sh2zCmPDKjgVS74NvydkXQ3epkBjLyiY
pxg8dvOV6OYdQuI7C8k06q0fkTAWWb9LfmlPXwpb5QxmilEkmBcX4zFmBPo2
tn4p3ozbesJs9IBWx4avAPyVLkzWfRAIV+LmdpCXFolVUsCKagPOUHL/BnfD
13vE7fiI+36yg9HATtHIHGFpTeZzPvG/DjnYbadFxsyQZYiBjN90o2wlpOgl
/MVcNAMVkbZDjtH4OE1Op1aCDddufPy2hHgTs6cB8L3TVVtZb8JJ6/MfdNnX
PjH4W1WISNFmLj2gv2/vcXT32oaPuTv4ofpwsYUTp5jZZzTrCqRoiEJJnVC0
OtNKKmBwPaGZ5pHn1dpbTThEZ0NuijljdrnvUALz5WDVjws6f+Mo+F0pVEHV
Zuifp1Myx09c6JJV/hAFUvTXCuIHnzPPESISs2zlEuMga5R1bqtzh+C9RZgr
2OjMCvk36mtdycYs0QBEYsUDXTcjDnHhv9nim3Diy6CWQDMq2LtMnL5+wNWZ
qiE6SFuKTeHcy5gxFBiZMuc7lt4PIbJQEK4sVUG+gAJhaF2Cpx0/YtAes4W1
Qk4nTETj6+u3xuROJe+ery5vBAaiyVCC26Qg8qIcBo8R44GNEc7NxR1Y8HY2
TzeNuT3CzhJsqMSeF3TrgRIWROL3CtG0kdT7OyDaBUQDaAStsdV7gqCl3MN1
Ubbs9AqOSzUiPvfZekAAryYttBQnF6y03OoDkorOg1DUuxXIOiotGWRlqzY8
Ymny7EZWWxG1CCdMnW2ER7nUqYo28hDGKlI1SD1vEIadzH6fhA4mt3FMAgRv
KiIHzg90jEzd10EPYUuMH+btGdWTmEiwbN9haXwZvmrkJ9xRYuJctshL0/9d
FKMhLSaFVJylkgXrOROeLnJ+++xBymcNXpLm9FgB4kFkJJj0kjEBo9m9G0DD
DlPUoiwOIhsSkx7LmSdYIyms15p95M4rWaitUARsmKdQ9dzzEIm9azehfySR
dzLT3+2MhMATvJkZDqRWrLwagePm/+IUqhznCqaeF14WfUDKAd9DNM7Is7Ip
xDIAKrIcXijEn7q1SMmXM2+iGf5eeHMGmJ6N2OL5C4QbeeM+Y1KjnhwO7J6x
FwBlPdnVAnzYzs6PTJVPpNxFaL55P9a+uI6B8A6Py6JLJz5+2Am2ddDUV5eN
5E7UzhxyS/TC0ClE2+13HOk5EH1rAXUzCM99H85dvoRvY2NgoQZSWrxkZFti
eWrBPhfss7UMFcgiYyy/fTPMszZXhdwsYQgDH4OvOt0vtx65KUHdbvPgZ1JF
UzPrl2pbj/hHnsuqsvULoYHOwGKRP9W+yahB/B7O6IrsfP5ukDs+I6Nq4u18
QgZ8zNBAljQKOc6rpnmAZcoEsHWdpvMPYkkuaPIc0Bz9HB1pueLPmen9OArI
Zi3CRIRuqSqG3kGJUElu9XdqyWMv1qXL6b436pW+RAldTHYoDd77BFvUxSj2
Z1Drg11sDSSdIpvXKgzECJxc6DIVt/N/AowAhv9Qm4k2+EU92gDR9AbtBrzj
JHVgewgr9hfgDjUN3NHK9SKSZqQclW/XEUhQ+NEHmG+11Y1BsYFEQjvWtl2e
Bk7smfwJPGZyOHoRb5GSZfeVgRRDcOfekydmi0H9l82CahwcoYjGLzBkiAzd
PUndfw4fbzRpaPliyyldFnfCwV+UG6K/6qRVKq+0m+4obJ+DOfeRkRdqjIOi
Libclsfbft/Zr0hewdaskw4R1ZjWvqdzSJj/6hDn9KtWDQBxCfCh5eacbyj/
bj8IAxDisbdaHN23Dvutxd2KWsq/DhzORl7YLtGcCNY/maOppQQGuukv9PAo
qOmYIRRvZR2pijgRr9cjT3mVn9rxF311+lgDqzVLT9ncDBn0hP9gVVd1oEE8
Qc9ekY5b58FXczLF6S+tdj/x9CMee1MdaK7mjrmKoUXQG92Fw9rtjUOM0edt
kewVLJqQEK+yiMIcTFNXKlztAFS26mcdl6QwQb6IVCnXiuSIZCAhM4dkTl6m
XGT6rfwwMJPxijEA5Az+ugV4Xz6Bp/eoqGZyelWKV6jayQVa6IGFYhqnUs6N
9MIHeWCP8U7vypioXJVYqZxVfytlz0wNLekfLRcIXvEawloW+TQoxBI+ZLff
hQCt+tK0z5pNnWmFyg3ul1aJm0o19x9H2bbJlrhBrh+i/fVSxTRPFu3a3Zbj
L2SPNjwDmxoq1i28bc8Bw3HNt4oLhfjYe3kTH/A7xdYV0RfhdigFs7DvzLMi
Oe0lBHc9+9Kc8UlghgvH8D1vQLqVhD8tEfVkgiRtb5s9CEdPBtTUHT3VfITK
p62WrioBXj019+jlf3irgx8FCEvK1AqULZ2S047ggxtpeA9fXgebYo8SPa/v
+v2LfNLlL+X1+KpxIMU7OEwIbo6lwNBbrtcD9QZutyFeWYPZdN3EUri2Ksf2
jxad/W03KguuBJUyhqTMf4fe3Rpu+hbvrZZ9u1GztkyY8tPjVcpWutYn070t
xd3cH+rArf+Dx1+w4vnXrmaLWYfC5YMbXZ8V1esKNtT6AYxcP+/6JhrpGBmB
/rfoBbIEOnqJGoCprbTlq3sgJF5MddnJg/JFV3PGCzfHHybmTYZfiB6DxWvd
X9vAkmCWwsD6gGjv9loftO+Hz8K32X35qJ24D6kMAQlr8LY0PP+2Dr/hE3uo
w948KLkeqAsaAhMRJSFPTnX0acJcyeeV86+uvaI6MQr53s/KgMGZ9qoId07J
c7gdxPfSCJGae6tT8lEOPqcX8qyIRSLIWAoioWoNoBORRzfdiuI+DYVZxITn
6tWp9Kts4y6Tlxb81iFuOcK2ei9jFRTOuzJ7ce4xMArWeRl0GxQXGx+N5fr9
DLcjfj01vp9BvpBofM1w27Su5Mwrqij5hWJCUIcFL+0k2cyPGCQ0CL2JOUa1
ygtTCEOY8t8PbAKOC2iWJaLm9LhVSLHrZXT2hvG95KURtpVuPqeJbBRAYGrH
IVVvQVapRrJvg5Vzj4krRJ1aBVepqiReNIFT7vBp+L/MraQBQMHAMu6PBErP
ZCtVP+JUCebbi01784r2uY4bXV0e7b1u+JNjXfRRaO/WJEiYaF8942PTbdKQ
tOVEwRCzQLKkglWoYM15O2iYw4b+15slfsJrwM62DD1jCiHSurBiW6aFHMiP
55YcWQ438zriTQTiRnTu0AkuS8F+D4MGmSCC+ZOMvEzcE1uQydKMrISZCq4j
cj6S/U5A1w4xdXH4+c8kh5D3bnRSlt/vF1qt4Vp/2nnF6xjwsr6fgx+m6/3u
g3jevwiUZ7xCEhhVewGF4FWv5nPkyG2xEgmn3byzAJK3w7bGU5HCoOdcy1uX
1S3mW/BgUcmi3KV7M9WhOnRdMAKw6qoByCiHbB9cJpvQvZh3SXv0P6+Vt999
pQTw0h1FU5HJeD4qzW+df7yj+1A5sqd31xZ/6h5RonXrgV6htuqu5cmeRfkf
FcPayYOWoTFUvX0++IxU5LKgpv3RGgFycE7fIpJcBPoElkXTfB6mcyLLtKo3
bFEiYRtGSBsjiBNjnHgXMYmBtgtVzjIUY6LGVWOO0jSxf6exOftInKefLpg7
Afj1bMO03dAnT8FxKSTaQsGwFguvvmOd9Kj8cOec6JdoVRkM+C7+v0UghxSO
VreIISLRhSm6EfWQDCIG4NTfsM2Dqf1Eg8++1frO4nl5k+Xc1nJgJU3+b+QZ
CKL9cXi0eyb/MnUuwbzC1sDzSXS+0unj/JM6QpK/Mrs1WjDs1gz9FdeQemlV
/KZFkFMq9DqNx44UhAX2orf15tBRCdVFbVTSyJ2b6a4QoN5jE6ro3G5uiNu9
SlRxaamBgzJomiGhrYrpYFcQ3J9WuIDRYXvrgaHKkByCAstlIX1LQoTildak
sW265VdgytDXq/vIWKmv3LmVH5TG1k9hhgFjR4XLmvcWC/rOBTPat/qNqWkf
Bcv6vHJ6siHvakP2uiqxSffnYKlcoY7VuNC449zwTCAX2re144tuxJXxc3mw
Os/lvQ0uBr4ROv92JBAkGkPIeNSlPeI6LDZr1CRdHwMcbbkWaiwp5cVa60ke
5cm3k2OQAvtrULzTCkhBOFoJC83sPbMjJ8D/Y7YfhM75xJERN3rNSDQ/xA/Y
iat8ruTu5gvpK0dz34qD98Iff5b8XMfgtXwSEyHpB1uel4Pjw8DKKWOWQUt2
MJCfZD/YNOgnTNJ4RmR2B1blohlJtV11mCdv7EzYRJZzcUCCWu+po7TDmtDX
ojbaS15KLJm3sbxtC8F5L0f3ZMtgLPAWbvwXPjGX8M7j0HrzurOOM6/NDWXU
DsC9WL3P66Cb0wlcQYkSjhC2lCz4NkvpKerrt4g51e565fNGoxYFb1TOJq7l
CekUxrb1RcFGp9M6e2hFLz/nMeLH1bDiP0WIEX3yaJC1mZhnwFssQSOJ/xx2
louksMd6ev/GJjYyjNiWSHUSPyf3hQvNRTJuKC4Ov/kHdLKJxFPZORJN1iiC
d6VONqKR60M64V8qknG3nejAEZdXOHGSrF1UL1zrRPJUspSxdN7+g/blXtNK
cF3bQG3mAVguX2gx9cw07qu0ZxEKMXSSaQI61W6kfg/CX7OmK40BFmH6ubUz
zLKTUVBS5XkvaipceqA7vc2ZMP9WQxBu18fASvpHWPID5N0w98vEWt/CWWk6
+23TjXofd6K4zbxtl8RubUnW3Yszw+b5hcvaEqomHlGABzf647hzFD+uFbZT
4jNMlnKkd7JsE3PZtIFQhkeBu53HUcJj9M4yg8iZvGEpyCRr3Wk8AxeqdVbg
430f8xKjFcYm23xQIgPq9AzK+nZYYx8eaSP+Cl0VECMfuHXRRVxT10nDdp/Z
W/KrXkT9ghWtr6SUEjuS2Ln4kkYOg+Hk1HBRGgW4rpOP7yU7SzEqsOKx7b8a
8gSyJaHlOoHiRV+p3kXR47aibEE+Kqw0y3Ze1h2z3kmOv9cW2RRwgph7JnR6
40KD+zq8+P7BcH754UEHFjEkelUvoGK117Tu6iFQL22ZdMZWrg+oZ9E/Qoob
1eoZfsaqYUQF3An+Hj7wbEVphbHxXeujBZ/HS+uDHSCyQogEmdhXgWQ4y05M
t8cESY94tOs8aA2bs5k0PZthyNey1U3bkeyHmTHd74IUDXtcLzGC8MG5W+wd
OUALvSaD0F5RjiHvBlHAKAdL5kfZqElDG/hzD3/atRw395vuUhCORynduA1L
z9mrB0geJ/0NHRK31sFI4zffli9iLJrNHXr5LyRZvm9/6c1p3Qwjnw5DjEwm
7dcWf2mX0K1VPfCQZP/K1ndajaiI3osMqdtyxzP8GPC3N3RGtWJcCNkhpH7a
iL1gS+JWMbc86nMBdU8HSfPKRPXvT0oWLxdC0VF2EDTgiCVNFsDokEJ1o5P/
xgTqyddDvI5Tk9/hMYX+rjFXKc0O+5f/nGj0pFxEwo+IXJacRSWWy6rt4R58
gHsyDIN34SPdGF/BktEAi5TzcSxP1QrIY8yGo6+UZKZdC+S1qiqaNzTx0CIy
urTLeyA0YPjFaQvEiyaVMtRjiwnV3JaXhQcb6SXwBxeFlb0hfvjTpvGzo5ni
zA1BgkEWI2DkT+msyD67k2jMBtDDz2hRRUXEDvxigD05aMaBTq6Wmf3uCMxf
Wjy1otbB5l/vrtjMShT3hg/aKRvR5ORM57FgGegiF5vNQm16gbUHEzx/Kiik
w/mihlCy2AACDLhn/jYWJMKBr7YzG6D/eoweQjO+9kA/22BUOPARJ9eDRzIq
5MONDfbww+rGea0si25Snda5VB19ghttEaprtzxgvUl/bTLYA1y4D0GeSRQK
EKyEhF2ON7V3zM2pNFQTO9VYTW6GRCR5k3J9aPrRGBnEFYTFU76c/6jQPU80
px0r4fIka/BZONwaCyh4ZdHm21/xTzfbiSmSzQtJU/ld1XLZd8puDpMcgBlH
LqA8pec6iuJxOkdZ+xGoW9FS0bcRyRqdbjLiZUWhRzSXylcsbdaSajyEIT7S
sU2nqrDEDVZsBf8mshZ9mSApKrDSPb1YhXfT1apMPkg+LTokOAVOW0GJGM/W
d0cLXHsxB1ETitJXIc2n+1plyXkryYiMuiKuwcy5RLRkrQFA+0Mv5zf4tCY9
aYjKP8P/FwSAoJjroIcJ4kT4QdUQFtttp5a44DVbzW7P/JC96qF3LXSGriL3
k2ctb94kJ8AgGaDQz70w/uamrtfCFu4cMKzSk3R+gRDgXXLXV46psc63UHxP
ywgSoBqw+6wHvG+KwrncK/pusqZS878czmYPsKjkRQTMpKqZRDsMsHpdGrPl
z6jhuFD4RCT+rpfMR5qQhRE6Er23wb1Mh/7Hk4lDCvYkMa3P1oHnDEe9cmAf
vwG59qR37FqlyTcRcn9+pa4sqaoIl05YLNVZR9qn/jmN+LIYeiPfYA8GY68g
AeNVuRoTCoLLCXocdvnAakpNM1Ek+teQ4yH3jnSPZUZct4B6IozSdzZ6TWPh
WKP6C4MLHxb45YYF3PwOuZYR4sqPtx6VsrAUUpoZx305Zs3N80bxePzHlHfU
NNpQ/yxrnnhkdbrPV2Q7ztZ2Jg2nqP9ZFuBCchvi2xPwi1MHLYFPk91wNNnt
TE9PBoKqEmJsfKn/MBdqrbAbJrOMCvZchglVsYB3EF3wI6wuNzvSevRBDZTY
4NboQHZrsr9JZFckzT2hCr+TToWC7wX1CPPOp/W+sqzGmX6WUiK4DodzF5qR
OXNDavxE0KhQhnpsZTGYEkoJOYUwUFqmnZ9qK8byaQdW9NsiJp7df2EJ3T8y
mLAn/6B8yZg2AOPWajYf6cXjuZBwH+rkWr+W7ePJvEEqT37O9H6sd/mumE8z
zmGA914qbtb9LNfAUiwjZEhvhOCa2jEaGBAjb7xU7SK+t3F+kgY7UMlhev+L
WSxh94S6SRBeFLgPtxfLdRR0FBnnBa6Xh6Y+hWaoSGSyhsCRt2j7EmBjsX9Q
xJcCktknm69NHyXfzU3oEChDU5aOrAoNJYmO5eorchRzWW26QPLS1I9Esqep
9G0ZTfErP+yOM/hXacbU9zA89U827Ll33FBi8Fd6H6bfBt9+UnWZD6HjvNNY
TvCGqcMaa9geBGXj3BOSPJYR6dlqhi5n1cgTreOKYZqZFmqmPQT5W+8aAg6q
xE6H2w5lLeKMD1pjNJlT0dxjjk9ZBKYVFuDowC6BCNwNdkGIH/SxdkYfoIPk
8hhW/v2UEr3xQgEIK662Vlw/i5AGGOfmsLA/x4OnQb+KxRgmnPjMd5IPtqWR
QN8NwK71wp3Fb+ib+80eGJvM7RloJlJWkJOOCqqNFQPmGFIQiIGC1L82oYbO
7PvVmVHKUOJfHvkRMA0drIC9NKruKGE6raQz1Db/EuvNNBfMwpw1yLMv9MIt
X8+jng5KW3jjBpRKmSIzuOyhwFOzExz8tcWXipVGZ0odTGli3U6CBMzB/TCF
az/plGTOg5qcFy1odC5dHWPa9ORThw4kibtE+MfmC/VXYtjP7+GE5vpKK82l
BvZhbkKIzqDrD7FUo8+hW3K9vdgMPlJ7+NjOvN1ODhCCVtDyk3eWrWjqNMq5
9NIYF63yX4N+ZD05LON+xhwoTq6thcJmjCxj/QhI5+QFRrUozm//z2r/gJ4C
BFcTkgl7PMPkRj7fo+VK4kbTmhupaHAxIHux5y1biLw2CaKLX9HxuAKNC+A2
43X0wc55YDOqccm/C0/yWIhV/FnzrZuodwbgSUZtDssbNFNCc1iH1+2jU/yZ
1O+4bo5H55uXosyyketpQGq8cOT9ePswmHukXBmKqKkC9cOXZHakh3RdcQeM
PRkNONyWPiEIXlXQBbw7aepSe2nAt3i6arPfAjhW6dwcZR01TwO85Omm1TuJ
ulOPoTqKEiyRJzzgsXJbzKwuFG79fNmo5pK/x0U+8m3mtlQYQYXTnFxv4gL4
VeAmcqLC4bweYvpw4w0K422Eip59oEr7FdglBw6fT/2wPkGkRZ87nsJ5w/64
aqabfTz0Ac2oMJ+87EZajBz39gVst12AIWD9XGaDUNDs5qdcxeLHcMYYz5Vb
S6N6rNUn69m/myiaIfgDBzeaOkqKpG/JVDdFsCCWbZ+RX/HxKpBULbImw7zx
WZl4aRm1thZnvvo9bNcKfLl3FvdAqnEGkC3JBg3F/x0nsPQ9IhcDciLTNZRi
MaLqdHUIuAtRmX5ymH32vVajPuxl3rtBktqsry7H3AL6TgPByibNI+vp6bBL
BGbKxIDA/Er/uUqrFWMmh+VoP4z29kDYWAEj213pwxmPINVSZxjUjjelAGdJ
ItBjd50AZvXePvnPZ3Mz9y4L5UXtQYN/xmUGousi4msRBYRIlFyj7cgkov8A
sjduvEaHH6r2UXv0y+56LnPUgwM4o/Qw6eLk8pOx9VgHx4zAImY8aFKr/K+p
JqRg6jfz/zPq6rd7K9y9Vq9W13A+dg+XN+3hNnx7ADUAYNgDITSK0+j/PF6G
A1S2Jp+KeCHKWB4wCszOwJZKZa4GnMEQZ6/EAPpJTM5AAzDRFpfZLinFpC10
c6DOePCUud7a2BgylyIVqYV3zwBry766rBJZyRQAX8kwxvsF83uftpIgWTAW
xJvfX6CkmupnUVfbSnqUi0AtV4QxN9P7m1Whj0eflkgjWYbaSaUbVQXYE30P
3U+4dvJ6gKoOGmxwefDD4zSBTB9P/apLV816o5xYzbLKL22vFl+S1lJuwaiD
ixbAbACQ91hPG1f4sxkTm8pWaOA910QrTRgrOK7aehYiwaWA5UJI+8gIH3HJ
OYz2G7wxXNn+5/Rh1kzzT1VFbtj16F+Q/Nsr/jIbwTdx6HVEgzINI4Hn2B+t
CKwoA+xI/NgC6ixsvHzt8tXAKdBEZyNcnF8gKn8/7Fcorod+ZAQ570LK4MPK
A2ym/feJwlJRkDGuPajdHqf58ehUWeu0kKKg14CBuChcisMIX178lbqG986l
zOfV0z49LU/9bzPuzInRGt6HycuKs+qemH//DHj/fxtp+9omMq7pd1ODtdtN
vbg63Io11ZmQvR5MAAIqj4XiNyPf3a2ZHa+r3ys/CqrSE56Be+rI8wdB/lJ8
yoogIM11x3JwO71wPG0ihkG5x021eMKCxug53KezW/QOAx4PR2wTCp6afYLm
uPYLy0BYIO384ljgdBVy0c682tbZFJXqYEFkRmH88yEKKDHV+jhx90u8XduD
52MvxmOhFknipgyuUfLrqA1r/QEHo537sLc8Ar1QoDuTGRZ1IY4TE4YbsU1t
nt7uRfygn6MaqjhOagCAqut0flmvoCcf51+uXApB1dQvbN57TsUGkoeZh2lJ
IMLMovUkqrlyc4HiMXz74OFieQ8mcP9KTMB5bJ3LOWeAXXVwaFUT4LBx+FN3
IIeRyAFVNxA0po/VU1v6TEUU+Zy/Jlc2tl+vp3vYOGyG/ckhGlNCYOiAlyl6
AHOGf8M1leDFCIv63BgIyX2B5j3vVGFs3odP3v/QYUsByrNbFpHauFdBR/Yb
lYourNWE2NeLbth/d/YuDqQsux3PxUgw8NfwRKxT4+khYbNBhVYXggfUz/FK
rlxDfR1M+s1NGD6WckOHzH/MUsnzFf8HhtkyLvlasi2XpV8PXk130awUvyyz
pkyKMVwTgJaLKAwJkOe2+4xAGLuR8CXpTm+D2vojZgDN1foXTFdmyJqr6SWv
ShEqm6xU6fHi/qpS8fUeoJ8TLf4Hm8A3VfL6t3EgCqX0aS3GZWkiQybVs+BJ
41q8BjnAqExULm2xpTNhymMCg3KgmsksvQRaVby2L4nLBaiT6q8O00Nq4rUs
b/5oQByI8WLAtCEFtOYZzSE5KP/VmSLJGgsJyNlsVb683n8UdXptrTbJzp79
0tTG+MTf6JYcfD3DDJw3g0Ol5GGQv05/rjXEvcD1dGz8zxZa6aBZymC5xbJY
7Xuf2WGgENoOBwGnOiha/gy3f0WSo7iEUNx8Q0l0EufZxMAQXcd4OSICKXYg
7WQEtrR9nucW4DBPYS1ZUWrtiWG3B/8zTcTmmsUFnnanmdfli9Ol0GocXXDg
WQKToMY1K+WDEvMyiydX5bHnXqQxhse/r56nMGjhGVb20i1v20rInWlHSGtX
n5dtwdo/9qJIkzmygxkg2yd7+J1R+A3105BpoV6fCFZjkCdWas08fpNGfaqr
dUetBFPdZ/R+/mVgPXCl/uwSjJt2Vkf9Dd9oOWG7+oSJ0HQCTSsAceNjpMKc
38NrXycbh9fJ4mfTX5A0E61eTUqoUyXb8uVFex75TPhso+N5SzHDYkPeWZNt
cSKlN77WsoNWJlK2C2E7W8Sk0fHfxM0gA6Die3J7MEOldzpHLLAxaIncGqMa
gSlPRjMYaArGEIum8kQ4zV6pEo2kZannaKGpyEnNJU6wAzE5KNVD4alYLyVb
6sam2DeZ8iidgJRR60JJmS6/Ry5VKXOyHjvgHDqRoTZ6Jm1pPvu2Kffd2pkF
0NKzSaN1IXwfreAYXaauljjZDceA4Kxw1/5mbl3pfscotV94xaYV9Tx789bR
5OKzViRwX46ZyzUUTKsFaSeASQ21GjLxCUu/LH9ypE5GeiE5ydXuqd0Le8K/
LKVWt217GbDpQnv+lZ3aBDMXfyvpB/WlyP/lnYmanPX+PBm+bwNH/8E9695E
2DuJ6KHU5BFmnqWcRFBrO2NJeFaO6RxNlLsj5PAu6/xrEdRL7077vKHj13ci
mwwWNjQC+Ig/ui82jdlHrb6zyXRAAQGTwZKxb8s6BZ/P6mWzjx34ibIwVs0p
+on77fQpwQ22ecJ7EXXaWjgn61PTyg+0/gk10Q/dmxGtZkgOOKHtghLVWiVP
09W1PMmfGl4TVXNjqgKJyfrEuPUPjzNlkZDUD8gi27iG7fzTPa17O6MuF1yY
ORof1/DM0cQUQR4WgIPZJ7VZj78aTiYFZJt5M50S/N4+ZbjwHCcJ8aNHXfAe
KqLJD+juJDhgQ9ikgdFCbMNXntzuJY0+FGfypNYm5SCFhbeh7lPzu9RyOuVB
gksdqwzdMBWZHKM2lisnBZYoxm8LUA+QlsEKJTT4nrzYvH9Nheqzh25o3gSP
PSOCpTT3DP5dydNkvAJffdO41JFwxO6/5tjPxE2I/igb9ZdtooaQcr5z6yI+
vZ7VmUHIzuXQnLcLPQnTSAx1e3CfD2lyT1JZyerRmgaD2aIB38pfhyL5S8Hy
P0k7QFx6kI5YZNzPYgN4hZKreyeyr8+SJi7ifoj9ssbcrwhKvT/CURW4LN0h
6EEdV9AxzEUwH8IHZqTsFeeFPv6/li4QjBTUSvKburHMmB5lHrixInoSPpsr
PErTeRidb3hjXUZfwMl5xZ9dFfWc8vXQHmMM3XNhkg2xiDQprWVY5alZQvNj
aqr/zV9jS0r2OFjlVd/9MInmtkkcWReMaFsRRtcH0f4+cAUdynQn4Wc8zVJg
QqvDh928PE4MOAUZj+pMew5bOkDrsFVFSFcIQ6gM8MASrh/say328I8isFtF
ZlEAQOUR8gP3FcLD/PIGQK0iQ7VuuJq/7dyi+PUhd2cAG+iEacA6wvhAeHUt
yEvX/XHNbVAbk+CZMaOUp1i/Q89vh86KHZ3YWawjSIiGFyttQgfXQkhFBWbr
iLdkR2hfCq2fTb+QY1LliazgXYE+yA7ov1YKytZ9amnj+RcaMmZ/Wthxi4av
GmwqP21fiXaaU5yWSzPTzV+9dSKDHAOnmkfGqRtBi4F4SwopXCrtrCKc/1c+
MWwVE3PvSkWB9+biSSlDoHQp4/r8wCupsuPhiu2fAqZzLyz9FyJwb57XlxqQ
8Sy5lR2g7bvfXP55LgLH/H5pCWLH8sMAgeXfqobFOh0wzBKIOHJgaDHvMToZ
PA3xhmGJPIaoZg19U2wGuUx4B5K6rkkoE/Ejs7eVRPpan+INT3NclcfAPZ56
myfrvpIz2iEvItGsR1jWnNOJLbCXDz3JbS1DjJpEXBPXf30751Ws9XBbCDyA
KCtERD0T4H/IuJo2NzxvximNKDLXjWwyIYQuYTymPEC72mFlI7+nC/sBjgfv
JbEBKuFxDf96kL72UUEpZOnH4ZdgLTuBgxoQIUKJ1NESgHclOfMSgYW6VL0Y
CCpYHcqUDUWOEErpLkqj4WsAZGs0vwo8Q20ptzNsfNKN/lDSAvigxLyoodeg
Vh7eDiUEyadc3Ma9r7dRYLQojKgJc/Z8Nw0Gg/OZ7lP3T/HtjZPwpXGo71Wg
vMbeBcqYNNSPEePgto9e6kipXimLBxtSnjCyOa8dbFGaPK0gqLK/GRrCNyHA
ELBRoVllEM65elR+w867VkdW6M+JXfOMUaJhFibHTtgdYbf1fG8U6jok8/uS
PlozYFedXQgrHPmuz5G7SYUsKtSJ08JwrWWr4HR1GPGKnC+FS0sFqgY/Gidm
XWHJ4csUB6kYFkWa3dgVkzte9unQ4IqY56PLQiqmqJK5/bbanA0p7fpbqwEz
tLKcHGFkFPLK+D+B7X6IIvhenrezQVPeVz5qnhfVlbGcA/SPys1pGn5Sj5ED
18zUKOYOCv6hLZJckI/xr6dXt3+HiaTJt9/sTa3ZWLhFXqHwESBkNMkKWEwT
8SsTVYwxbP0ODGnfSQmDQaZRYe/GlsAc1Ys3JpXIDXDB355TUfVJXLgSL123
u+K9uCpilsipcm+tpTd8vo2Uv1bLw+0R99FChB4J8PYijj1XzUO5TQXgvCd4
Z9I9U3e4ch1yvFjli1Ua+RM7ky9XBkpHY9JwvDLgDA3L957K4GuN3uo3XrK+
7JGdb1UmGgeWcG9hU4RkSJkQTqETdFlxFdQmNLCPp2C4tmAd+s1WQGOnWzun
kOiGy7JP5RgWsdRYjQ0FahHo30Fvx2ttAV56SnwcahtklORFQ1ltK19t2miR
ImKWPiCCEB6Uq2K1LSSlYtYmif60FLlYbAe5IkjDU04AoLb+IlZlWNIxvdKv
oEiPxQjmSn64fU0kSKDbWoJqfJMNHc1TcJzNrXyDhz5gfwn/DEaQ10DkE2ib
ZMlwnJ5YHmCZc7VutXRm4wG4rzwG44C9QbrQfMa8QB7rOaaWzT8L8ejfMQGo
PHWChyV5dUph2IMd0YGZ0pMivI2svUleS7gT/j/AC9PPjqAZ4EjU0nTHeArr
QZ6fUez+fNMP8LbvP9jX6WpNuIpzpA3agd7MGSV7FBR/boEclW+lWuaTlVWY
OvNcXbxTZgAJI0QYmfISJiYrCxOjjdlTyBSwMaDV6K7Fg9yh5ZwTZjyGmn2s
oCx2llE1HLJqjrAiK83S3zLUEOiUuePUVTXScG7JgWpw+HEwdqIez5ez/Tgh
xuGZjmLixpDs4ciDjZPPEjjC2lkPlrpt2ShYSvVrKnYWhBX0MBlBTx05zfgk
dVj3hJbaL3EhYKnPricTsqnKqxERaPv+rU000WYAmx6Todt4aeljqkYio6yQ
K3Arse5T55jTqQRel0YaI3bfOtJetMjHLTw+F3PKWRIxY09N5HSSGwhJ6kqC
/fn2PvWwmat98hVZusGdJlnFDlGqyj3ySCah/DLKSgynDXtoD/cB/vVfJS5q
8Is9FpZU2XlYAm68Bts6HtLDyjks8OHQs5t6dTW6Z/fYP+Z2U247Of8kETjq
4B+wb4xb2u7UM1MA1AJE9w3/bT8X9qvhOKIpkWNpyMbMAQ8nS3CZzk1SY/0A
T27c5W1Og1tg40VCVJKR0Sagz3ZuyvmDnfJrQiSeCtrx2HfYlN8i0Op5WqZI
0pDJb0jJojaQH2Uss3eBMJHNt8V7gcXDN2BKVSGBAxkkxq3Gva9DnnAIO3jd
fjcrv0v9KtAsgf6JXcIkUv+06pzpsmKpuXwHANBax29w2nfWrPYcZ+kNVN43
FKCxTKuEnVugmA5NRvXZWpptWFpgA9vchCmQvFlZnDiUgMP0OfvliiCnxoyj
v9lQfjOworrHVOrPUw5v0eWsGSVJRMQQnuGYDf9dr/LFTM9J6QRydmxlLctt
R8MJ7pDjqAw4sXyp0jwLyPYt5BJw5UOhTBFux+pM09FkdLxG6W0h07TmUcbW
8qlvtJPSgUq7uLxIhBy4Z/L/xTZV20VElJuJFjV0ee1dI+qP6I1qbsXf/5jB
pTB4KDxoQaXiCd5N/hY3pSBeFNkDmhGC38n4PakvuN5LY3OaWWm74p2OxM5C
8oyqyewwoeKPPRjUT55q0sLBXT82xEeOL5lYiNb7tCpvhHokn94XKQdoZCNu
Xnb/07rQCmDKCbdmk42zOldTEoFHUHOwdt+cco9vPPMbuZXxN870sDtz31RF
EdzXZ/KMcU89VX3cIo8JQrYERE/5NgsvD96G6spaFIiODQjnLALNzEMfFA2F
fs0odrGPfrkBFopA+SKz2sfaN3/n55wzkRWKlxD93qsSWRzKMKZhTPbGFCoo
YINJ8amEv98x0wKRYgcRETwi5DODYBITjt86yy00JQXbjVBTt8YW9X3k7GFk
yhd6HNNw9cQuqSNenbs4F/o4xUtEsGPMvO0Y/4bB+fo6iKozMesZNsI8PM2w
3Pf6t0qjzhZPZDa9zmzh9XNjjTnCceIaIdWFjXdUrsSYTdZvkBALhjGOJQ2I
bvcokil27S/59b1iPUu3P+cJkkNkwzKXu38R786b0IiL10zDDY8K1niOZwu/
i+mz67Mvmt8ya7XfJ+OJDIwP3qozgjSBQqyc0JoFzXHoCzuH8usoZlkluLTS
VqSVgVa5XiA6m6mKdnucizYoarmKeYUxOJTh3u92K2GPg9K3LwMpfNaLxLZX
86CxU+fH2M9e1Qnuh9+deXl3kAGKIOWx2pehgB2XTxPuDMAgvKo3W8o4FD9X
jnBDOEENyq+apue/UmMfJ8nXmgah5T9oM2hevhMIxDPdA4MuArz8qT74EnDI
MkT3kWTgrEETQYe8X/msaCDqVjByi+lG+4OmT4Si4/SCNo53lkKibk93Kawp
oLfRkJB3iIsULv4N0/ZKipvlUiEZJJv6iz9dKWqAB8+0tfgpgV72JlbCswD5
YM8M5YfDkGSs/Z+vdI4y3GwwM937b65BcFK5I3jf8oJZcjONe+4rzJSzNUZD
V3+wkqJnHtHn2xt4j1/eiKhwMgytiStvY6SJ6zyRp/lFALT6s5LMR8FqPclv
lWsKjtkfCpgBJ9EG1nbVHvnGPYlsY52FhHbnrcTglpvDNGdW7y1v1dedIqt0
mM40+sn0yrzQltH6x6w3DAMADkfHiz4lmm/VMfiFqfAHL7oyT+QibBCkbhH0
jiseQtmQ4/pOr6AEDVF8KmTx/1Fbc2C3HQ1gKxEYsxxsUBY+b0dssCDHK1ND
1ESxIHzdQA5JRyuuAww+6EwniBSdrViDaWkTFnMp52a4BMz4pSmTMPI0SQeD
Yi9a+UPXpoVzViJmHU/6dt3qdG/nkYwS3c9QZYxCXrEKSe9/WCZcXEbZsRIL
j9kG1vzoOubscTzePvufSAWpPydtlgdS3VtqLxdy2w6tgGym4HHSKJcnIxBG
Pru7Aqi9i250T6180KTI7rZk1KwrF7fQGI1pzDk5w6dPZD0Loh1Clc++XBgi
FwN7HvqbrnVcZHKiV3GgXidClmiyPP8xVQYNCEzaKGh8mTxienHG4lN5jC+g
8RMUhxMtfgdEpa/jc6j9mQmEQFILCc9fqpdapKkLG796OWuYYA0OhB9tbxOm
FgsN150oZvOxSxIlWPvsl3c6qOjy9wBQdRXaC/tiBeitoC63dBnC6mrOe+Xl
T+yuhNMxRr1B/FRhwDTm9C6BTFERsCuF1mEk0h6exSaCz5gc1YUNcRc22VD3
rJgZ+uFXw7VOM2ch1FstwAQHSMPKpvGuLMH21dcQUzyivEm2eIRpoK9KP7tp
Vj+mWCWyuRiPwgNM14eiOeF0jJrfiKUBB2meE3jnQ9JlsksEUQSd5vByzUXg
uCRwRo2+HUk+wG38USHYOQvOwigzwnzTy44S8E3DRx3QgcVqfsS0C6u4sW4m
jGsq4HM51ZOfixVFxWddqQufWzpyH/Tp5kXD2yGW8qIHb+Vc9oosGAYg3f1e
1a8BFl5R2EImcd8QoVR4/dnW/DXfIhcFEnqTynWg1rXAJBHUHu332j8mzsP/
I2MLE7uelPKHNt/zjwK0g5pxf1XlXfr4oekIxnNnIytV2xiFd2fH3h/BVFmL
XujBRFzfCYZwmJnfPUFY8JTFsXsJSwp+zVd3GiDl52MY/LiekG6Ts3uMKgSW
vWqZtUOh5vf9CWw+axkU88HslJFL6Cu/C6gybctafJ8Pv5EobKeCfn9s/aOH
Kt2HKcx+dGvhfEDsJCYCAQ8aCNemiz2IUbfO67ydiwkGDAFbYmSQu6COwklS
Hjqz3h+k5aeureiZlMQJtYPlvkXOzKMOZyZ0Y2SXr7hZF9ASI50UxB29NvnS
vTSwLL1weDHUosAD9LPHK80PtAw9WaBvyvu4/TQCXSCltakY3J+PvS4Y5q2C
iQbjhCxjK5rw4Z+F7eIHbIQx0XTGJF8X7/yfCCttjlRnNzKj5YsZshysIJgc
i88z7LfGTyavM2z4LjMJT8b17Met68P3YnNUDQpNjdNYdGFkRSr7BGxCYLdR
bQE4fJA3YU8C7NQ/JdOBswrv3eUZHgPFlUNUAR64vkYmJk6U1Wbg5I2AmjNb
LIpS9Zvp1m8iF+C+wo2fefPznaZA4NXDYjxazB/iI20FlJhV+O80sOxsasHG
fIAEZaB0HtxhCWuqRdZ0VhWJBQ74r03DrOSAz3Fnoj6k2E6ranALf6V0D8tK
31d/dKXhv4papz0jMODVl/SX4mvGEH5kFvXr0VuxVmkdrrtR9VYrectbUdes
N4LovKCwYDAJutD+/FsBTGXBv/i/HvHhtt1tHbeYdJXNKbb2i8Zi8ngAsMaQ
0n4621wxrd8c4z+OaMJiPQDLTx6IjkkazhHzn2DDdCQAHs8uM7Bqcn8Y70u2
XESEwEkNwoj5FZREy6YeyS52N2MqTAIgK95qYhJ2YJh2RM9AMreMPKL5H7uV
NnRI+lI6MnQhi8D2H8SaOG7qozfRiENxBrJo9f4CUIrRLxf0JMdqXEfNCgkF
zksEr2RaR9xeTMYkcCfLHvVViTaKIEVUqtiEACh9LEXh1HnZvhE8WJlv9kUa
TteqhmqvzJTBjWIyCl5ThjzOAIxPws7OaCKdgDQuyg/QzRkAPq2hebsQZIRz
9Pi3HQ2uztDFr+nErMSZItfpLswUsuATRLMD+eC6k3/u9ImyHHRuR1v05WVC
iVxHBQTi/6em1/fU+qj4VzWVf+mkzZyV7xFIX3k+rZOdcR/XehqD3ilBvtqK
P0O6VLPWYii7+ewkW2c37aRPtY2ZO2C6mI4i17MiNJBzhQiCHkxxin824y0f
lPP4AP1QiJX5Lw9AJlHJGITbc7VfEL2hrI5wxZOztEeI0N1LkbccSL4M8dKz
wTPCKwVX4OxeUfGpj7r4Ye3t7ThQK+F1F9u6xY2uUhK8EEGopFmxYeCEGKJq
5OnHoWtYxhxMJWKgVDuxnIhA1hwuMnBqeF1/uhed6mj2YpEubSNAge467qK4
bm6FVy2PbRj7AR8q1Xtm0p7iHstNgfOSCmWVy1qdIbtlcZTPMnX88Hbc+x6S
1jJz8j1L2hu6jYXUyGBtFPHgQPmRIUZznERpBeWRubqLrrPQftOQBH35eQtc
kVN4JcWllV+O+GzrM5fr24BIoVRah7KU5xydQ2o6JH7rSb1CONOFleOQh4Vc
ODa6bsrq3WAMRdVX7VoPCscozDb7MmJ96jWj1kawJI7+RcJhi+juSCldQp8m
LVQvO1uawiYqYk1ty2ROw4iSc+24jOrhSYsj3rRzEHd1QlU43i/fh53nCOa5
gthoiKvB6zrqEf7JC9f4UwTj5DU/sRMVEAF0gDjm7kMV8njg5IdajqHRcwun
HYCXD5g7gpW0rJay3OYmpoT//Uppm0pFECYV9gFKgQDOtPP6N3EsvWOh+Egw
e2gxnBllmIyUNjU8Z0kLPBqsoaaNT3oTlmxtJOcX0KiWp6aiDJB/iUCjlFI5
cyssjjyrTyUH02UhePTn6xWq05zdIiToSm+a+b0Rnpayp52UWyHn3JQVN3W7
Lc/+yQhAgAUSWB6QV6svGXout5lEwUwDiJh4XSFSDi/kfzhBOMYmo/CwGqpx
bGTHAt+SjO0YdU4+uOvCMfc9kFXi1xljiaJIg/CD2xg0o5lA1SWlOO5CLU+e
NNHfZcNdj2Qbbmt90OBW9BEKkht0KLn/vXjCApLGcqlRJDFeAtYBeROTiPiK
7nECtQAMRuHBUqPi4r9kadkONtguZEk2H6D7haPFISPv/2sQZAalgaYhqhx/
88+KOUXqVzem2yqHSXlzaZ9TT2gi96rjHM/CCmKnl7DPkU+jyYAPlAMU98eA
/8IDELMWPuRaEiswC+Jzid/PRip22KoajoBprrcXBByRhrwwt0gg67ybi1mR
0R6G4sqhysaID6J9BITFqYVBDIQu0TF0LBKDN5DSkzuzrWEuzF7DCZw7Ij5N
Kbjg0nllE5whp7c3DCcF03mtpMEunLJTuH252qvg1JcByu+lrpK0ytdqbvsd
Eoz29VFbJ6B/RN+/WnWRxxItjDI+cbDl8puEjc977FqwL78s6ODCQBhk/Gjh
0z90DjGF1oyGTWIaGbXKbKgoLPR1ha8sgdNR88/0qCJFbJUQSimF1LkstWzo
1QeCDytrL8jOeOfUUCFmW8R2bufZ22nR2pS92M5MDlcWjqqeq+3bq3fzU5xQ
HaLnd2R80ehBRvAMCB/9eYxvaC3dG6ELxFfAalGIuqJlMeBsWf7V9Z33EvwX
sqlJ3oGS64SEv/8VW7FDV11OGi+64b76xr8v2cHhzJIfo8PMOjOQoHe8t48h
k2VWbLPM7Yhx/Fk2D/mHK4i5Jgpk8SL/V58KfcblvdSeeYGd9eJ+wNjZLBzW
X8XFuGP4rIYaN4UyJOE5W8KRTiUTNszdBdYNQoQJb4V6JrVHXpQoyLyYIGhr
tN9mKtAiOLiVmxy0D7HX0KsTaHsSNXbtRZjKMgflBz2p5GqS5dIW9e3BuQDu
L8D/vUVYI/KEdAXu+S6GouWdQca7QxzWsmNJpqZECqFby5wFAIG6l3K5l5vi
h1h4HB/c0L9haeiUDAK6eoE4vMdheBmGShUU9FHOp19Wb0x58k/ADqUPlItG
QmM1b42jJ45UoWLfnAi4FO5WkA+Xlsz1rp/K73iDOwpZOUsHPy4jlAugtzz9
i6N1mbATsyZuXThGe6S+ivRZCGhtdD3bD8LJOvLNPe49kJlZSMQlhVSiqgjF
qc4kLBdI0ARYQNp6vPQdD5GSc2mBEXVmW+Fn4qZ0gp1tHi0VaDb1XOHTOktL
l251G7gl2O7EmKspSs6c9LCBMDnT2GxLJe9qO/qeIFlUW8EvfWqk4juHRyyu
IHa8VRXGpiO1Xg0bUdJA5MWhmt+he5Dj2j1iFLAyM0QSkjvGBkfmDeAxiYgV
QI+Rl3B/u3JUgs4SEzvmPLRvt0/K83X47riSiCzXo2+V4RdNo7FaYfq4pZUl
HBcrDNltRtRnK2F/FUV7gOMgC/QHhd2A5ppgxCutzR1qO+CsNFgR69QiN+61
4Pg4iZE+2es+/j9ws24nbWo5+TEFrKMVWmUfY+8dTsMrUihGdz3lkhn98vlF
tOsspQHuKv+R9D7FCMIhiJlnh2whsYfAKY6SwtGG4Kg6/9Dy8qBHsjhTcSIe
89mlg2rkH35Yl5tJx3YWsnzCzHH8VzLTfep0W6AE1wCSPaykAEnvsZFp3E5t
yQqGNptaZAz4XHtkrQPyH1GuJn2hI/S2FsxrBdtNUD2v3VhsqN08MZKrDEmg
JKopCfXr0phqqfF41DUOX9YfRZ2OF2142/s1pcXesfmr+94JLHAR5DUsedEn
U7IDBVgdrD6PIhPNeDrLphAeFrVri3UUm2/KulnNVlUfAxuwsVxVgzkfhieb
nxEMbyFDQL3V3zluNqtBTEJybtSCsdKCJheDB4qrCwAcNuX4NmTnvmq88LzC
TgiVcLuhDztwbytuulG6eWnJGQrYRJWglrT2mVhxLT1vM5OHS5hJynq2Nbr2
oP9TrRTj/37DI4ZndeM5RMRH6oYuvxsy2vQMnYvbAmQ48PSae27oPAVzEwUI
xmwaaGv5afE5qjWERTiXWRIQEE/W3Yjs7uD3V/KWUhsxCsr5ZKSbUQkGs1GB
V5qptjfaGi/xYM+EWre8kPlrjPjvrdGvyWIfsKNZ+jaRBz5kxkrj8iAynBR2
L74O8RnDj2Nmq9unwbraD+bP6/1LU7GltT1wulM0jnyMzX0UDa3cEfQII0Y1
tEI6PyY5YeSoRRq32LnloWnKrhL7JalaPKOYsyjrs9zQbycM21/OWJ6lbDji
mtsd+3X9TIj7nLAhluNnluwovL/xTafAXUlm2v1DMjt6O4jvTtk2XqfhKqmp
H2vbcp/KmfjkYhio6I1fbelLLpJFgOyb/V06lc+m+QLXtpEqb3yJxSGcCqJO
7MI7yVpBXgEvKutNe33gZXjXfsoxiEYemmaJvh5N+ww9SIBlsTt31vZjO33+
fDc0nt4eBkZzRCpR1V/IeE+Vu8L0KG1EA4oigq7UXB1/IWycgPL7fXecxMsO
re653hnqggXbkpYaqosJcuDzU6LAkFwfgxlWv0b2PjxzAOnsDA6EXUacvZA+
XBOsrFh/oO8o1vJPjM0yRV9JC9Y/rPhWO6x8Se7H0q2Oovj6Jfv0DkqC0tzR
mb5fYO5TFi9redf4VI0rPCtfjQSnUk6AITefx+t6YGzuT3h/eMOOpmIpWiEQ
0NiJ0EOWYH066IVmWNL4chzPjNxbhN4+5Jm6wdZXC89BFg/vQstSH1orcTUJ
eaw+JSV9YQsvtvXbX18GArTinD9pgqLIosGGt2asq+FAa7k2W3EWcpXN4AUR
RxnY4rI4Bw3oqOpDrvMzcmsNYM0QVGjT5Rj4VfZxZB4ExV0GQVio0EVFI65/
rFROUVuU+ywiaqiqDQ9dFNsqvufIYSoA720AGUGfB+vrGifWXPqucHUvlYeN
ajZ7pkkjn9US9dwd8ooM9A0vtnPeNwZk6uFJ7KXEGhL12XPOpsMeuDAw19Wq
OB3BphlJzrYuccYehMcMLHWkD8kdz0p+D+cV3qrZR47CvMA2WWQR/runUdZC
xN36ado/Z+ZFlkZp+KbiCRJMAqmbVjl1Yx5ZQrO2x5Kvqc0hKSCiXamYNHDi
oTqRe6OSUs4DxT6vPNWn3uGyljdpYwOzfJ5UzF5rvqS3n/xCLkAzZH4Dw9Td
TUA3Eb7+9Lihy9VrN3YFIN+Ou+NdmiEgOlYFCVPR63+18TfxA+9akAAUtBa3
RsV3F4Y5Xt2fMt3f2E8KSWhF+G75MMQXtHObVjwqPNXRoyOvRYgWaqLSrvCo
ZR+f2ulxMKGGg28kbPCineN9JRGa94OQZtsJvKg2KfFZDFSZW8WmMuCNw7Gr
KibUWz0IhPwlN1W7LgzNVDpVS5GGNR1tah2mobNI2lW1bgn8AovJ2gn8vOX5
s6ydQ21lRwJARjXtdf43eyTdWqrZLANGjhMpq3sxek/UykSDJZOgdVyJEbID
WqQTWCRcWo5m97uulGjg2iEHXQXYJp+f8rcucFHVeEKi9QTOHnbpX+cL9Tsk
p3pMEfsy7RxNrxbgo+APcsFndgcOBCJgNLOeOsnG3qq49Csplb9dd6CDsm2l
Rctm/oKcLuYF09MFBaSdprUJjiAxQpfp9KzvgMcuZDl3w9YpSlET9jRYSoIU
h+EhpOIyvaDXI6rmU+iUFG6SGoJz1b9+nuSLdE0iOpmR7JZ/UM136x0CFfoF
CZ7+CiNayvZBTB8hYu5Lk+L+qcruAeKbQxdKboxitln99qcDcJwEfMC0lSwz
JKPKrIzO7bSgBljqQ0HpO3YJ4lJfLGjGFAVR+P6Tugge7JdjVP+mDO/NSefc
tXBP3yWGomrRa2F1rFZpLmYxhXd3XSziH9Mly953uGzAmTVejPyZFoZYOXXn
GAKC3Ns+huFyTG5Zk+F8JEJltIJurvZepF/HS4WDD+nbp/a0XLw1ID4bVg+I
64F582lbPwpdCPP2zWNwzR+wQjmV4Lc0Z2ZD1NAMl/DfRCYxOpfoUcZTW0wi
sAWo/ihXWx3QIvt6V9bWgzf1T0GHFpMOm9umYPZbrIxXGyCKIRxo80MD1SbZ
e9ATDoh2qdQ1x+O8S+FBgJ/yZeuslyZM56DVU5YnT8zoFdqnuGk7kzYhmhHV
N+meyKkRsH+tBvQZFNenJ6XOW2f1KKN4wOcjJsUuzaGdslczbmi8RzoMfTcS
1px1C4CLUM1Q8MK1w9i8UyelG9KIref2zC3Qx8XsgIeWsvx+i7REhkH9tP/K
+q5DAurNw/TYNy+27PMW8Dlh2g8+97g2gRpxt2LwL+lZDxWi6XPbKlsIlHTB
mxOt0Qi4QuZmj+HK1qMhXyb808ZV27119mt0L+MS1NiZzvRukcdE6B1EcBg+
nSxSXXKEo0Zf+Wzlj3Tc2N0kXdKaNkqXW0CaDbyyttn9NSZXA3qUoaxTgvuJ
dRXck3j2088pu4fImP2TTIdMYkVsxIdNYWA48Yd586ZlL1YCWcGBQI4r/Qfm
n9Ue/+Oxjhj/1ZpALoliJRuxqptLHYtsAcVHR8xXylpkJrMyCh2AHpIxlA4E
r1z/vNDRCXR/d0tjcXYcQvB/LNwn1FfKyFEkyxU+dvseglNtLySrb2D84NsR
k1Ho3BT+0Dou8b1Uinxtyj0cuWC1+ArbBVenkueRDA/XOUzVZLVj6gie7FFz
il3Sqzxb0KKfyfBwVi8T2zIxIkv6kwq4/XXg+jE9upSSTpy/6eyWYFVrpyxb
gu3raVXmaDrkuoITLkPHTNhICCwXhZgF0gtFectSIE0VANiAlDt7UkcP16oL
P6XbWOt8I150IejP0rhVLM3kXsrNgCcge5mWT4My5TfMaHOhuaPHz0r7UTeX
aMDW+H5uQT1PtI1d8nvpwqJLTE0TxQGYAcbHp4K1kSBIcyaowwhIsNBEFYw9
1ue6+pCgr8esJzLtvMffciKSEMbVzCjPUrJWMDdiWkG5REMNJzxPcyVl1e1z
rhsCyNYPbwcSsfQzvyNaRnXJL61Nyp7z3hG7yzdSo6m1q4apo4A2qao8B5Di
7zniTl9p/5b3lbPd8SvGwoe1UtSOHno7KIEPUI+O5axDRKDkmnzirRu4ZUSZ
VrTJH8YXRyNmTN3AqZbzU0PPoijrozRm7gEnB6QPXISgfKS4BHKAq0jIDdPF
5Ev313IEioz+vvobb0xx8ZUl/ewhlm+kd8kjf38kMRG3sLOIbRli41Brum/e
r05rQV46e4dsS9PrJJ5j+aWDWWGo3R13rZeDOmaM4BUXjrhwDeVmuA11n/yf
pnZ/HdeTI6klQTEXPyrm6wq9Y9fNuOkHkF4tu/Mxobsm3qvceSlqebXbbZ4I
X/tMldRQT3KttfJ0pRgGU7a7OQter9ptKpIMORgREhaMfeVOxGXYjZXIik3R
3CfVc127hIebb4cAnxMCj/cBM75zWyS3OdESU7FAPZyJV/EwGoNRUeRsyBBL
8S/yi44untq8DOSaVQO44x3EXykTo4vxv1mVyeUOlNPwdzihnlpEEoo6kXa3
8JTem3Y90J8YSyjxKUHkpeetJh0DO6AqfPmN5cL20tXgPb184zLLnQoFcqaU
79X+ZeDHqzdVi8v0C8ISHdYiRvzwmlledcEAMcADOnqdCBejR7rK5UKVJ3Y9
Cp66//954wc4kxcmHHmthsOUePePyDPSKMNV3bfFccUSJvLYUPX/BnAtXGPz
MAkQrbEwQBTb+YFSdA6ahxRUh3Jzj26PfQAN189yXzSLR9eHhhDubYk+XZe1
2ruBtS5kqFOvmZrM/db9Ep7QHQIw4u/BczghFVLbfYGLFChZB9MtpEaib3xD
9PyuCedqNejzoY9SF6K2KO3LXHFJ5MicxDsd/uLBxnKRXvdV8TpBwxHQv9l/
cohUlnavKbITKDzOewQzlvCNQjwiJD8Jiyi+QG9tLK58ew+LWqw3V7bIX3Uz
GX9CpHBtyAgV4wDS7g5sYjQ1rLTv4NOL3FNFa8RTUDFsvz5IUfT1JGFbX+ZZ
bstJOC/OkEOM+2ycNuYQaU+8by1LNP4MYy0PIAJunytqPSAv4DBjRgN/emEi
4Q653LgSRJgKQvLMpatG8FtTHFssYlUcv2RCvwoPRW0fGnVHukBOI+hGRjO6
pVqybz3W9WQ++6NJGIPUfwVeAz7ESq4M6g12m2QS6Tep8m4MFbmfbV1QxirH
mtuWyWKjCIy7aJUOHCT9u/ZC86pcNUWdhNNrMZSUYTaGYyisVCkYJqigNbko
N+ipr2Uij2b8lPH7TrcuMJsOHKp8IMJR72sEh2/W5wrx2PH9veDB4PcazkHK
boek9l18kUdCyQAMg8CLBwHzZvXLQEwMKsuuatwZ2UhRRUuNrtIGVIF3+M6t
hk2XXSvdJf4lbObYQLEDHjMKjqy6mDHIp+uWd1HTQeTsVr7N99kzAwFSoS+g
fkCMYnf/H9ZT684NXZrT0Jo5MANql2SAbZ5ngxQrhZqbwE0FS3fWGa478105
gmOlh2iDcuPQb3b489wBJ98RyPm45CiCiivWfnuSwcPuutVo0a388Hmm48yx
/5BUJMa7Ub4xUWQePAP/wJXvYKu0jiF8FStWEXX1k6HtKKKjChiVZTk8JnlQ
zh1mOPLmvgeMZAJM0jveGluMDpjrK+NN/HH5AN/VC4GgbmF9BTOsfnomT02s
fdDT8XqpMk3XVRxM9/h8B6e9wdh5Juq/3+XItyLzUlgeAorJetHEazrHYOxQ
S3jDFoYMfJbstD3JwidkyxgjJkhdGvpGDdwQLDLfLiOSqvIYcCecD+IxoMsw
bYM/DqAeE53iTsyXJ0kAuqsU1i2cqmt0v8xp40Fonb5xSt2EEVD1b8nKnjV5
zFjtCOmpZqxmZm6jAf/7onSWZrE92vxfCwBJWnD3Wzs+5X03ixKNGUx5Ez5H
muMWz2urzDNz4fsidelNDqCmimixIGT4NVoBdGmmWHdYpkACh+QGplsJJ8Fo
5OvXrMet7UD+ZcE+ZSVpdU6vDeyGrTBMf1RkbM2ZPdMTeUbbydECF4Kg4Rbd
ReipIpg1BwNqFq89ihE24lmHTh8d/h+TJbEENglK+t1JjwJlhgEgdD84rouD
pmCEjRTp5c1IAflQNyLzJfKmkOFdPmIs6OmW5UzabNw3wbCZhwOO1Cm6iicl
jEnE7L4aLf5OvEstu30U+rPNlzWFYpiBczrI+W3oyM2Ixfrb7p06TXsN7u/1
3TObLKsVC1qJn2GD3af+tT7yZ8xQr9uPp/imfE1S0lyX4EKFiXdTTCv+8nJ7
1cnbE81IWRGnyesOE3L0c0aZ8BqZmRumlnQeR5lzePTBVXyPotckNylafG3X
93slP+UBOsSvarrRQkwJglKqY0OLI0svDZqZwafn76nAbiXPaKWGammjW1qO
KceducJh++lPXbUgRLVnkUC5WYLuyZduQSKJVvTnZtwqQJGGC/BqVoAV01xh
X3Wg95fTAe3uNd/oz6i+jTg6IWlmE9AamHMpb/Vw6KZXMsujKRp5jvY+POYy
Ujuz6uy5JVHF2n3D0MwT/cSc8Mo3vgOv4EQ4fMZBGT16KoHSmH0DAFuvX+NH
jMZUoTYv8J5DeBUZCV0fQl8tgy0EOQGigqorHD5w3SR9nO9z3RArrjvYiD9J
NXHzfh5WHQVdgS5bRWoxSK7vulRFnmPQL7GSq8kQf1Sw43SrfYZgnRuLiTaL
ZEghLVP24mLCzukYwBRhDZNWFAx2gALZ+WdvhmOTdljtWGJmSQ67kc+jLixD
8txNnrIPEimpSkHcBrjnZfSP9RD5eiZgnWh2QB3ha/a+A/Om6HO5EvKk6C3J
qQHAoApYZZqfXtv0bnv+0ZiY4HLEM/dhwgFOMqnudshnvJPb+sEj+ZrELzBH
h8qhv3FpnxBe8IxBPpXmu5XH4d4+XXR7EDPgpP9ctmmOIL3q4sq54Eu0Ohs5
GQ79JmWREpVTSObufzFTJgTMSG2RvCVgcW7L8xAoUJYVYEWq7vqXOKPUQOed
gIc/lcI/zhgy1/TUQgsMLybXDGbrdnwITpTu+oYeRIq3OwyGWadwGpC1j9yY
o4O+MLByGTkopFVqdV+yn+9p33kEjF5HxtJ6v1vN4lvGw0ZhU7V7P9v8qER/
ES18gRz5O49/QbXP9SIu3jfi8APNDoy2Aev6u4ygO5FX+uadEZSudc7qjpcn
5MwNQaO1oPXNa6+6I9X++e/zrVOWtwGdwnFlkfqpAgIWS5ByQSO8xXE5cNPC
fRHpbKq69tKZ/ELRCerfsRJLE1XE9LrlYAB4q6zqV4kzsjCZYWGZaJiVVhJh
zA2Yi6OBtVUTnisw9iDk5Ji85GpHfuswrZdU2cdkZRXxfESHkp/FQw1I59Qh
2dG7pxsWrNT3zU9FdQDwY8OvAnpwBX2c05xkfoARCZ+gneE1enti6dU58qaO
5kItSgpRXzplaR6F34q3RK3octmx2KOW4ID+wRczTtRwD1ZzK38HNMQTmGvM
uHUA0tGf441o7WJlVJojoyhM5mVVtEN2se90mZRxoKlFWChgAldFW8cUshHN
YLKFBev9QULO/TpLpfVrj2EO6susGIwlEaPOJpHLaolkj5Xl/TahKW/vocFQ
dU60vOPUKAoOKc5/g+N/yXeiFfh7192vJ2/1wZAERwumghhDdIyPzEn99FwH
bwqSZSCnq2NPasxHV0PYDIVqNJJIgaiGUam4E1fEgkE6RyP9Hbm9e9u1pEuw
AhHmK6a8kuYRUvMMYjfl7SxhsFqU0IZyJ0OUnEvQvUvanDmHCKNi6YqG9Nhn
7lx+HmjWA5tX+ua0N13gA6bY6/Q47ybwt0BEIyKtKvrPjFqHij0OXmvhLoO2
XV87xhU4DAi1PheAvK0ccpsFjIWeMJcXOEcw0V2YCWfGVLzucQLngFrZAv44
dZokK6AxHvGBji+AbBnwlHQuFx12oYWQ8oDj5TjKSIQqYMhK5q0H88rptku9
+6YGPBlHeXvoBJI8OZzA2XH5Bh40rnm+vfJcFuCkQ3LlcFAkorfymjw75GP4
o/9pRXdp+53IFj0zENFey+IqfairdiPKSHjs1CCYD84z9epIRDHmwmwNMmx5
pvwN1p3KRwHMk0MAxVkT/JId1OgIA70vDSby7XF6EqHbX8nmhL7E7bCmZVzf
2eO8WI42b5nCwcwqrpWCI/U3ctk0U3XTveLBT2BBvNvNkdOcRkNm6NV2C2jH
rpF3qq9F9iPKACLlPhUL54xVOIuj/CbvbEraBU25p1oeV25ySVXuN/OWbFD3
MsVtlBQkmZVjRrqzuu0vwUzYJGgQK6+laX3I4D3256vzhd28IC1B0P0NQpc5
9coJMv0BmdfxvFFRtSH4xXs6gaRAAu2kYpKl1/2atEJLKUCYpT00L81NzxvM
QwMmFnmg4QevAX8+SiL1UV2PJOETKi77fuvTU0hirSHY6RWFgUtK7S30qPD0
3ddESbj3DPeavof10R2snhNgU1uDd9GZYaEqu2e31MzH4xxvuUCD7APq3m2L
GBepCSc3myP0AuZA7Bol5JHFYddm64weJGUW0+AXrUyQSOAS8Wo5US8Qsd54
Zbwz5XN8KJajZStxdXloKw4YisT8Si25+u1JReZX3VaCJ92AvKb7+XQ5jKRR
o3fklJZXEhs6Q1A1IXnmGlqHwfbz7SvWkGsKs6tif2We22Ot4kqmUSqqFPbS
N7L73NGVmO9WC2PX57nGrBzai7/fwNEBC2YXVEjlmEjwDLP+HPNf52wkkQgH
2JXqyM9mvqotvlphCjug7lYqGNQn2o2PlQzXDfR43g+9inAtujNkXmShqr/6
/GVHda3grH0VdyAmQTLyN7ZBbi+stXncp+1vanYjn8WXFbkPi8iDXv4hw3uL
GgnV9R7KYg2ZNvQ3qMiIObtI0ifLMWLaVRB+7stbhxlzcmrAwHcBGZ9iX+pW
HUs8nqp0lxRJtxCr3xRPIR4sO+OtN3nw4cdJHBJm5GbVQTqT2Uvg50r5vv9q
gPb2Zpz3iB2phRr3TPMk+/5o/sx9oYEWJE1OZ70e9ArzVU8jamEBkdvqUwc3
dtm+oUYkoMOyye6pGkc4vWByyKd+miz33Oxcwc3QgzFtrsvE/adT4F8velxA
jVItic+mxMcmek7ZKpBQYfrQFxMOGc8pHRlRqwaQvvJEH0KDBykHLtwc4fNB
IqdWOvRzk6FxHuXGxQG17Wu7Vz70phwSWXlHj4sinFBWQMAf/7Oo8s5RdU+v
sUjsh628+0WdmGmV+MGqEQLwj0jbMhKftI51Bmi3JVxRS4uolDLYlwezvACH
/RC7INJCxghx86J9f2g2WtS6d/2qZNCB2HzU/pw6/inYXDI2BQaT4No669U+
6ZIRwVcRM0IhkJXuEj6K678DU4KUwBui13aeKBEWMcPiUOhrQKzRtPFD8tov
ackOkDmF9CHWEoYKsdJP0b7rzdJfI9+7wQvVGkZrzD9uKbn5C0PemuP4yW2p
PzbmiJGiJFVHEmQURFQI6dBF+vdbhlP/DXZ1mZbVqJvxlVSND3NA3nblKGtu
qshN19sQGuIiEuPbK9RQnIFhgfusIOouGbJn842PrHHLXGyuwSMMIY6PsOMQ
QCVSVrLcXare9DxRYyotcIvBr+7CM+pc681QxQApWcnMj1fHDLVltZcSdrhh
IS6A+9U5wKhSr9fvbhh55Ty/RB7uGyEGgDneIKrSMtxTAgtrl/F8iLaiFTMr
5ufkk9vom783kEzK+mrJVoyv8JLPZ3gvTh0SMuw7rsnbaopDKOmtfAgBjbmM
p49r6GWqtdOuJNldW5SFUsTOqhaBgeHU0hnp6CsgQs4P0GTsS/8MnfzVrSFN
8GmQjACCY/ShsYxo0QTvcK9pIwH/kUCGKCa35B+qDZZIZOaJViqfR3Ghuv5l
CX5glw3Wo3lLH6VhdNRVbixc7ZnVrzIlafP+VpxM9Y3wYIR3PyC7/iZoiTah
aHH1Pvn6SfZ1Po7jrfpkubljqX2347L2VvHgZ5y68NmjBxcnrXY5kw5ox4Fr
QwUIn8+0dDodwCHJV4hWE9gYdjge7sUd2KK7LOD7S+886CMyTv6u3nITtsPL
ZBYGFLgQndOrfVi58FtFHMni65a6onPd4CLmYs4uYJuwwN6saC2R2vEfGV21
RWKCgnYYhFV2i53XxZELp41JbS/wsdn+FZeZWjmzh5Ik3QfA9+7yd9HeTAZB
1XrDLgcWKhYYpNdTjokFsFzmxhJxJkoe8PxPwelnOysUm+sSf8UAvxAhURhh
1qXfNSsiZY5DkCqs5pIpIznMMw8od90695tXU4gJ+7wBHQuvscwC1uvBDhC2
4y728XTVYRHOVrJQ+FnDrQ/jNpTonqrbXsBqxDN4gIBn5yeeN+kOeAcfDofA
H0WJkAk4W4wWITKWOeoFc0vSlhwuJz0ekiI1VLjhLKuqQsBo0G8Yg9k39BYt
aAv66kSRWgfKBcW5Um9do7nPR5TWCVCtHtzGaANP9bEx+LSXWWtr2GbXDBoH
LQCZI/hST08BWGDhBXifxtHFA+jO2KxuzPLJ4uBuw/Hr4upBtmwhrfRs8Gaj
7rup6px7cB1zU68UBtmakNc6OujOFzR8aBZvEUuqcqpE7AGQI7t6KS5ysrFn
qVBtvXhHpBH5im7VKMRQOb8w8dzl5Pz1lKSrXxYmTfAjbP6oXG4EbPdfUQKQ
jeeBnvWme5RxHMn4SnX85O9NCKwbwukHJfy80X/eK286n6iq01nA+kPAKUeR
6y1B53Et9bKzgW5V0s6ZqcpVm2ZImOPLBgRUI99TwwU6JAIBxQaS4Xw5pWhb
oWuD2PXfbYUthRbIt0joF3Zj3Cb1bYnsUSEQ68V6G9LuGPoI6GxfWBMZEFdQ
Y5LUDWDfRTdiO+OokJDLaGboi0C70uqKZQhqHsClGI7BP4HRmqo1vsYdw0qc
FsURbQN/EqM3rRake6YH8N1oyNryKJmTnmF/4v1VORJRGImRX5/LyORatoW1
5IlI6VL2wZTCtsV1oYlh5Xi3X46+74F8Z1JLAhjdwrvx0vNSg/TdmJ0GqG2K
uaLj/Wgl+lAdftnwghouU+CdQzjXSaWcQY/tNTRfEbpfP+ZiPNrymb9VQ205
anxcj4GjwpzFnD+s2Kx3JA40eUEQOxM2SB2mYMPEYSVGh+vqJ2V7mZwUpXmN
rtsazv3Ol14egl8y9tJXfcu2soJQrOAENTaE3wP6W+nTR+G4ECjXaWADnVTh
3dxjxhO0lN6Sz0ltkuvw4q73EUvXq5xffzS1DQGGP0dhbkQqDUop3FcgpHht
q7RlCsCrLnxX4PquEuxBdqW9RVWhWBy9+EUdmngWhJvTsTQ6nMM6VmutQMG4
AQ5alz6IwkQc6zuhsrDKmLjC17G/v9Na/cyfex/INfKR8gPqkL7zVjyGPcZf
lpAQvSsWSjxrUJ2w4Ux9JAVdG2BjsV9BV+NOYzYZQwV+q8737KBx2eLkqaT/
FtgynOhvrUEqIos7O7mRYn7XYpBCiYrXa7N8aqPD94+5d4RgXXgTui/4uXZe
8EqKP8q+2irmKRRUmPPbhfiKJiYdJITU6yHJoq+p/gvRyX9Bpug9EbNulvd8
+7iI+m2Yf6D4bQ4S62fX31qBP6cKwfwiA4n7/SNISXDMQFnpqSUg8+uKXnGo
x0LqlQJrq4mYzIvo3TKujumouMY0AYyr8nugUED9xsFpYy5xi5wjWmoh+T3f
/VZiPnmMGdiEImoE3XsgEm+ruGosRCfefz7DVlgw8hcFej7HXhH/E7RBEQas
WCqPHCLUlZP4lSrAEdp6MULyQot+MNQo+VKMofPXoKCnv5mjLQvmLxJmS9DO
E0GwGJg+YjQGoG66KQq3lCILRwlW/5ljd8HZnEUkHUbVuOIQ4WUutBgmLxDz
60zxCyAi4zFU5HiwutSNz3DgG3zktAjOH27nqS/AEimgKadyN2XyEj+02LeP
+vCrS5k5NqRJxZQeiEmDM9kfZ15gTKexj3e8squ4TT2XYJMFPmu9y3MUvPnR
vS/OSd0xj/822+lhV/wVAIAHHl/q0qsbPtTnc2eA3055slsatsgHXIIQ5xfG
Z0vYRDFm8soneV3P24e64MEcMAZQkVqPOuD7xtEkqLc9amx0Kz8h5SpiXR8j
r/tA7I7kHKkdQ0NpZEs5G34F6BIzpRIZ4JIrpuifLQ+t1TM4Xa0GLDLCOwMz
2MUqr4Jxs75K/ggyr1OmspnxMT5E8+QyunBeigZsGne1BPCjHiG8hN5sWspM
Cc5N0LT8BNivbWTnKvewwVu94BjtVmdb2wCbYEDU7laZ32TrJIxSzjLTxR+B
U2egTf7B9F6VjuF2xSzoRqc3U+PbPXUlhip4FLWdZPAdGt0jZYCMOeyCztD7
S1wFYSoUuDHeT8mqFCYtYAWUaU3kpB2i9Ly8CrwXGcFKtT3CFsvSdeHuzv8T
UB6RB+P1vf5sHnbXnMCxC/opnzgZUH4cVKqxISTICNqmHLOmjAhYnvKLGMyl
9xPY9wWm4IVzykow2lVnZLOO2bYkz8Xndj1KLf/lLaDDivi+5myM/haiyUS2
EpVEZOYgnAgrOYurVgl4ZdMM1wmrmj7hCgm4VvGqdVYyEdQuM29WFDzGWdNm
tmM8p2EFif1V0ZBasbwwSnBKCv7njy5OIAE0/8/6zYGFbP+Vh3EiKysw/Hhp
T32RFIqEA0Z1E/wDmp6sEhS9e1ylTuUw7pBKH3l6VOUPAviQhojxRl2/1auv
VluKG9v0BaNtVOVcatdszXMr5SbWBLzHsO21wMI+unCcj9SvAo9cGK6ntXrX
dnOw06jQ9BN75BlTG87hpdOABEBRMK1juOeWugD1P150I+IWaExjMfOPZ1MV
LPE1DWWltajSn/bbRMC/dLb7WyXTc4CaEBnHnQi0uW7c7nKFw8LSXJGpEYFv
1v8vtXk3Jp3ufKk06hG2t56UjD4418uOK9oSDlIAO/tJGlNTMCiYuja7tHXK
WWwqDtyRvEQYaK66gbkuXdQAb82pLJmjmCJnKt+oz7kGS9FOkYea6WHfi1vr
Ke+lDxd5lBJEmLaW5nteSmQN0C3p8UsHp8WznRlL9mU2y7ifpwxbrjdBtmhC
wLRxOjUoHHkR0bkLWO4C2W70BbG+YIdcwVH/nuiM7P1p1XZA9/CW5HENla+R
iwZzCBfj4l5rgDd5BXrgrgG6a6c53AeMVrHL+Hdfz91TrhJuo0ziV+DQbM/8
4JBYGaWBlXenfQcV4uahWaJixuKP/yex3gadYurr6elqvyWonEUnwF7KH+NG
H0yDIBKdGleVkribnj5Qq+2B+DZUyLG+XxwmyTxwIRN5WMsaHPsThtv+PPzM
PBOIrdB9TIqpBJxsVY4+etVWFAEshc+HshDgKUF8gS5feIRzcj8AcxNVXnjq
aIPJRyG4BPl0NOQnTVf9Q6kU9jiWH42viE90RIO1c1NzNWA61tYAvlRgm0k0
IGwfBWFMOiQgTe59awPivMTIZJE5uenR9CMs3YJOlkIffrf9XEN20P+Nq1DH
HRYFsRCDVINnwU5jCJM26c30SOh1smLFKZal7pmRr8PD74ZZEgSzApoDNZ9c
IFrlG2/UOd7a6nqb/DPb1nehpry1PH/CjvdMVfP3/JJnb+Q10ueGiUuJtemz
wYL6FIUqs8eMyMmQk4EoSZj1a7LKE1mTP599VjuxTJ8WMhlN525er7kwAcwa
OGVfrV26+/bmGmFuEJEErFtcDOAXlFibkOiyNW4tVrFvryCOs8sdGsXGdmXR
gisvahQ6HMzhyt06pdNDnpsBBVDi2MIQqtc+w4fg4yj81jws1AsuzLgOxYQy
/t3mTPWZ10oolcs46DEJWIYfI961Zo/KhRnEzYzrIRCgg738AU21FKUs5dQr
+FiPzlgWz7lcd+4my3o4nP9iVLHCOeGngMHOMm4WxnY9huR5WW2fVn3Zwmtb
tVHxiZij6wwdTcDJNCqslXZHJJVReKTTOJOR91fTq7P8io6kA1vjzmmUXLi6
qAZHswgQgk1mIE03IR7K+lox3imlGJBIGShrxRozJEpPJHzRSFDfyD9H3SeX
TldzHq8NGy+XaDn4NMJCVesKZ9hCpcxxcblCeew7AW1UxU8doiSAfu3fP0WZ
mOM93p6QMQA9bKpupWeEZYX6IWByZHKwx0aOn8g7AieOOsXyZlg5kzX83YdX
tgjfGEi6Z+ihkXy5I1aDafQlvx1FzjFVoy2npBvNOKWNLXtjl0f3Uuy/p+J/
6Q2ooBhgVLE6bXzuB6yC3NIlcy2Lz3Fa3MApgWvfwX657JY0EuESw8GrfFdd
Bbi3OE0QN7gp8YcldoLKLKFhpyA5VpPaK3p6lKFM5xbJyq2vG8Ie9jZpgVhr
vCXvy+1f+Zw6h6pQszWOLBpHkcVfWgZ9k3dHeMRozaaBHWTInTw1aVwBQmqA
Yki9lyCNAgKZ/FBKsHYb9j/ZP8wPm07JCulhpgsKle5Q3Q70K9p8Etrp0DQv
g5Hhf7jplzG1MkMrstKOLirZk6jY9tQNvfxsckoXtliIKMh2F0AuwpoysJaz
QlIOAgpKStU5P2+FcR/irBLF6fPu2+YaZsASQKjwcccXTSj+/QxwbkBI5pHN
PL6orLijamSI1IQxqo1YlEXX3IXssoWJd+u5/NPDeS5eGX0OgzDMKjBQFRhJ
78cDx6875Ywzkh9ylJoMsxTHHPaV4LVJ/LDDgSzlraec05Hb4T2mdM5gLC7c
ETFYuFX4V/FV9UfYRe8r4PplZbzOb2jFBihpOhhH5zaTHSiK75ncLIY0Ag9R
iqyBFtjBooX7wChn453gCCcEC9d3wyBgQtQZrpwfEyIrTlFn1ONwSfEpFyS6
Sz/9g8muFr7LkFaUrOxsPNd3Sq85gtCTq3ej2hJ/+HAYFJ5FRLTH5cUepFsU
q3ulgOVFktO0BZBvqJ9BSTuBf/91SMMMIdKQHhYPtLTaGyEC4zFsdN9CLFnq
GGLg1DdK66StaIjgEfftKm6veo2AXdpBvImjAx+PLmJVGHKoZztT+MKX/lGz
mToY8MSsxu1z216yuYIi2hnxz6WHmS3dtPPZFnObRFmGqCEeCABsJUFgrsrL
mAVu4WoWW2Nm5Wjj/yEu4DiypeKYvS+ejAUWKiHxGpsdxgiYskvXBqs3don1
Rs8BSpHzrVF8rDef0CRyoGUPp3pRRMsswtfzHLLFxoWPGximGn7wvZlCdHAk
fp6jxFF46JAie1GlXg4iTGSE8SJpyYbUR0FQtaestFPL59W6zDn0N2hiPsr9
lbvN2Tr9KAhw3UrzhmPo9fRZnZefJmenAAgeeC+/z8kHeKv/JwvFwszOcmOj
OjBrbPyl5GvBUEPozGPlj+tV78msrgirt4y7S8UxoIXrHqyaPFYD10QGB0uX
+OAgk7lfbj7UcZrVgJQqg6jYedEI1A8Vt7oQSvKdLkmdKlFzT/OizA9VoNWx
a2sLyPO2jXLlL+Ngft459bz2e3+HUI0JQ6XN7qiXw1pG659c28s3vl5/T36h
6nUyxUrdn3Hhc6EVBqYy+UbAYHg+VpUEmh/uC/spNdRPyWdtwJlhToEiUEQG
J3uXbiKPufvN+K169KkzbQEDpYThr6tWBlnQ3jC3G4GVTKk49C0R3Tw6D+iX
ARYD53avFH6WTItA+oR3lfeXXiBL1K82ofhD4leBUiRwjY42CwH0gBgj6ntM
7PExrA4m4MEnqIdek3HqyIx40MdsuGwNnU1MWhPSuSzoO5wz8Y22adYgjhdS
5E1w4q0RuxCDoY9SXdab8KxhX0TNRUBhX2mm5TXnR4bjxRGpfHnsvCJ9NSH4
9gYEXW93mFXu+KpU+52nSu+4Q2U5chdV4OuK41KAEjOeBsiSrn182nAKxZbo
1aC1wNwTqvGMQkqiD+SHBTkXxag9qR8PnNdxa77rkSxlzUp18d7Yj4+A1AkJ
ACqsjOOCkNn4o1jgzjgLhy5jYHkbj185MFbbWmv0FCccsw7Jicl+lx8Ne29c
wL3sW9Q3CTdZLnQxlJNjYU/tPaIbGlwKtw70Sfj9SRAYEOhOi4NLlcOf3ccq
NGXX5PZdabLVVKJv/P7NOBNq/Pis9jB+lQWZUy0b2k34dnSYdnIy1YyhYHeO
5xz8Abhq96SL62/581mLBZ2HwDD3ygF1tTSrgfaSZQF7iVpVIX4i/C7tbVjT
5zGnW2Z2IMWB69TxaY6UrGd31qeELtgu0SGCCvnCdvsxT/CKYTv5yxYM2nbL
gWtkbwaJv2qBRXW9uogCmuJmHCtklLyvxVQGqKJWYKMKEfdW1XQC6YAeudvF
X2pJyOr5yy9lCSgu1X6HZoZudbIoV7iri/W2ez1dv5igR2leIcd/tcbUjtTB
02diZzbrwdMGUa3OU+AAoPYPjNN+Zl8clE41omrIsLTDDMLb3QshWBNF+Uqk
naVVMq6SPxikVoLBxx0LcxNHWLHSomeEab7qC3O302H2rNcUr1o56F7J8xh3
tQuv73or1LvmMh0t1WwtrpWOXvU/V0hrrKCdfsiiO8xRa7oU3WbprCPY8bsN
lrzv2Q6uH/QZO9d7uPzwbnVljQONaiy/eNw7TYdkZjeavQsxj1tGwdK2ltkO
68PM2JkFJSoP4zmqx8Dv0mpq22rXOTXs6EjMsCs4Xl7XNrexOgMWxEX9TI5t
pjlTHe8cN5uMlBGj7lY8MmpF72oe/ovO30vu/LYsUH7ipMe8GRnd007Eqpti
2uvDAJTctJIxQoFtxudfoX72cyK0gDpP0rU42W6DdO9NapAWQHqS/w5LvY94
MgptEbfPNvcwLZB6AbIKWefPYKT9oJ2wYyza1q6thcio4fgCra3NsRJ5pj8C
JZNXN0O0NoenstaQ1DHaxNJwM9luriU0bXFA1AMVrr/Ng4Enxou/FU4AsyLX
gnXXJnrAtQl45viAE3eXZ8QouY8VacATdDw6+MykpNIrBlqUkxvZ3Yr6v6A2
inoySRFl73quCrbyFcti4zk+vyyLxZPHMY7M33AP/HD/eXubB7k+TyPUCF5R
5TBn0pqV4mZKI/7Dlr/uyoOOPX8I3gT6qBP1ETo4rMBTeGRTFn6Ovb/x/jFF
bQMUg6lcnI1BF6CCpKGk83RHi4Mnfic5zFVYDtaRhBXVJhSrDSC0x8GgPs85
+lGJ0+W2TILW5bOshnE7ySmr0Cv0QCDLpIzdI98RH5M4HXKbP88+oVH7jJbE
vkPYHcO2SVSt56/sRJhdNOONIoCyo2b9rGNYzkzZpJsGkMUYPIY5sOvI/4bR
H2KgHhxTSPnTVcJFSbELO9DsMp+Af5AB+UwRmIAzbLjTfD+UTvzXixt74Ssj
c25XiSYqU4+qQnThKwIStZBCauJndC8UkMvaN+e8mDesNlX97WQfV2PsiXoa
SdB6O9CbBMC302m3p/q+MnEQSG+pSvQeaycS3+GY3Oa87KE29/RxJLueAk3S
wsLAlVGpBiJytDX3VdC1uuNWN8W1aSHN9FlIonSy5GZuC+yPre1h7HzJaoyI
/qESjMd33Lmyuxi4kg8rxiCQXHXxswZfI0IdIuIBwEQ1oMmgtbMHUFaHH/DY
RH4SjX2X48SP3ltY7+N+3zqxG4EsckBOEdSX5hzUoaqXSCP2PYVsIfKSUWC7
+3+2NqOfnQV/PR+gtxp961eg7Nl21okOKYMySsMpkL83citaKHSv4KJJAiNF
bFeyatvpdKEcnSkFASj2a92nFQrbq3h8hNqRZt28O2fi0d8B42E0S7loQsL+
CPNijkM2c6GAJiLGT3tIHybi4aVHkQ27wFlYrWYzgqagNAc8bYuQbSLVh3D2
+zOVoHK/JpVRqpT1NX40Jmr21kqCvlPzauPUjHyr2rXxABKtw7VyIge0BHzV
MzKitUpvI+KjcoCaYD56U+RA2/KoLoy5tSMweaVuRNfU+Doi/Q6sWQpSNtLJ
EGIANK13/eI5ya1wTSDj7ctFRcVK4cJFmyRPKHeaT6ojouXoBU6TIER9yoRp
g+zMxsAE3WwQ+75NVMKQxMJceDOoTNtmWYSa3Z2ImyqP0Z0YiP0gckKA6+sd
/fZ11Q5TfT1a1VeW8o6IkaX9rtiXnW3KjGas9U0m/ZSt60kD938BImWd7uVq
CwCGaKUqZ3zcKv9Jkc/jzcRUa1ZYz63ZAS2C5q+CWj5VeK2p6A7jQKyef+qd
apYMVIBervHfMYRLWgq9/zC26Lekg+6rK36SV8qpKyWaQX9GbOxh7jCg3JVd
4TZY5/KWP7CS7c2ICM4//2s1yKRNB6Z2d90bedpxS5h1bfDp2RRfNjjyvkXx
QmQIQgl1CfL97NbwCIsp+4xHZTOkxtLOHXeBNYYCT0XbnMWimHq2xVBZ3TTv
KG0WkfP2bYsoJDF7EApYqYrwI+le4+LwTr5ga5sdTVpcRNMBXELNN3bCVeC1
IhLWP6p4iz9A3pJ50G1HJsXwzX8BTWVeIJ1bp4YHyR4vJxoAljlu+buU/tux
Yc0HyXBn64KFKuUriUOTKoqvs2MRcvCAwDPDKSUCc4x0S0SadDslkzAFX5yl
AqInqX7HIo2lIIWnnzaEjsYYxRWC9D/l8kIH8pN/hweEBfZCXpQFmHnMeVN4
qwnHk1uV6yGH3GsoogmD0ZOArzdygmUZRaj1dUpMjkp0nkZVb/FKgRJrm26V
7psDWX5mrharKMt3dFWYEaDCo2SbLtErSGvLyfjsdSb9TaNAlwaoP41IMlHG
kroSFTgQXTx2tDdj4RsgCToFmYEpMo56MPJ0PiVatZfRfmlPDqSNnpSOrjH/
uNXJLVjGicJiAz+oSm5pbPJMnMgMA2xNRhA211+i0+WeTbuo/AtOFSZjyJvq
f02PI+zU+0nk4FN1K4FZzCm3eDdOoGcTInB2ayXJqp9g71dXi32+clzLpib7
/3/piTPKzHxoZyZjW0pRUlK/2kE20ADnAvKB3VAk4mqw0WW8I45DkbNtRdlv
GJxyi0iVo4u8HkWh0gLsTYxCbXykSmkaJXVKCTmafDffo6jJMv+xQcaOQGWT
wrqdlat+aA6VECIIQJeTNl1NB/Ub7X1RNjh2t6zO9JZy8AFTrKs/Q6aeNPPA
QKzYlTPsirzV0WRaCxPuwYLT7JZ2/wWaf8E0PoIAj9uE+dWzvOj3KnP8umg4
8u9uChkEPk+9KU1uSNwVyDran1G68kyiEmi45eobIreYeUNU5YjGtVgdw8W7
j2wdoOWMR6NzEUo72DZQ59ntCKN9xZYAmGUwZRrwVUKr0YnYuJl4tzVzmUwd
tWLek+Z15dnvKuwRK1w/tEIfHmRGc7EBW5hIcrricVBy1zpeP5n0dB6LdZy2
VFQEUUTnu+xYQEnWVGuo82j5H4x2pkJpUFsIvNEu01iYxgG/UZsMOS/D/6it
gFQxaocZoMtEcPfmYjA6XthCeMZoc1PePqlrudi4J+UA/PGRx+xsvY2aN/D3
KcXxyUqle7G6T8qg6nTBhu1ZrFMEKkZssbdyLDHuxpZasuFZmNWiQoIR3WIV
IEJD8DtWVotBcBhDiU5dIDau/exV+21kNQr9NVt2y9R8qDLpqwHxlbuaM64I
cfWQa4r97tFXnfOx0i/YEuNxgQbAkAlapN4d1qD4b7A4coIFINtPxO/qrNwM
QxIJh1mA6T5Uou9AVN83SDy0YauCcTu22LAoATCg21nyRk5wGahT7PoSXuYB
Fr6QfEYmHZbVsE93ShEzjYrH7N0MjT21V99QiImYUPhX125S0owdEaGahp1S
KY2AzdfOMEMa6KArxq+kZTazSY0LKNK2rxZPW7+vQlfwjW3CHZh3LngN4i7u
6C5MSlKZxE5r7+k8HtnZV97BuCOsStmLlWbCpDDJCm22sy7yuZe4kbBsr+fH
t2ET8Fl5vZmMN/wZc42A5Xra0II7ZK5tVofCi1ZFVxEroRK/yk6uv4oIfKq2
IabShKKNG/hU724R8HIgQA/wyELvsPUntf5mmVGmwMPgbqrG5HYskJKsjsXw
Nbo0ly6fT/dafGAFwguD9MKiM7ayckCm6cuBzGDMI2QCvAI4bm3f71cSUekm
sBmy6sdHQq8oMuKRHuxQOGmky4GGF7sJnRbroxeBc+OBH+QOleZomS8YR/Us
hESrVCA3idqe2AXYwQ443lKC3QGFnrRSKDdLLUcjai/sIRRRyjQqmBj/siBS
OAvgbdQXHPHo/WBe4rFzgkGornX1ymbgdCuL60+lK5ua5Ex5V7LRParGQu1e
Jn6Mao/iUaa1pNxwB1l5hGyBLHAzjCnzc2iAmGBVzg5qHtqx1oxfLHTvEMiD
Kz+zMNQk0VHhNMJ0UhF+PPb8KGcG9Q02e7L6LfMWjsBpAjoqQTRxenzklOPN
XB7/EtdKIRp2ZO6mLr8Yx8VfPYmKhnFpoNy9oB6bZWkGpBpuDZKC9UoxmGFi
097KwGo3ybOkCgmItzYwaO46prUhEnMZxyL5koDLBPM6gy0e0ciPkxtNiK2F
xzBnDEEykJI1s0oIgwyegCBPg14au9vABrIHynB5XUXC0sCiRJmfNBw5mdb2
QtdASCKsdOYOeW2QMjHbvStLkD5NkwRc6y4A5F7uQ3hbFdddzQjxGFl4cT2b
6+sfre7rm180xtpjw5CgoV9u9xActoIk+aPLwNgBxxJqp3FAi4ikJaGZTDYT
NfpVhZS6t2yO6u75FW3+Baox+7TzwS1+jt6ZT2tXLvrHkbFBBu9f59xLmazb
Bzgj/XneuBLz8HvG4W4dKrMHcqzOFmPV1ZLsPKvzppyN4mppLx2g1y3AGE7H
vH5RbsUIwlQ/zAWNdK1k/irUEHXTcZ0FuYTiTMymcc/FRkDgeNzW8uECKrW7
tS/zIueJAqAzpHNWCKWcSAD8kKnfbzYnJbQe87WwV3KhwCs3zzmGKlQfoqKz
3+YbvTLJJzaSrrfGsnrzSRTsf7ZGZutk5vYFCo+toFbKy6A6FiBjOP0oEPgp
99tFrY3QPRdb1txDus5HDu0vYkt0cEFm4TxDnvCbrm+fXKiOdNrn/knlx0yH
ab5GZpVJBbWhXkoyhjeluFilbAt+QykyqitmYWe5LwdlrsZQxeX8TgmHg3Nq
3FohnvFr8Rd9gj+fpRFqYsElM8uPVo/doYSuNobhi1A/EkXuoa0NsA2xIKIE
4cQ1DPXhrXbCDyhuyViCHr3j27d+PdvtLmixi65L67/wS60shmEqOO2ueaiF
4xoW0nuadr2VCmp/Xqp8e8jFJQlg4AD+Txkjl+FWJGOMVos8Rxyc9cS7db/Y
Qs+OKIbK4aWJfT+VIk1ZMMKb8BwLZwaZHgqcHAdzDiqF09o6C1XUfZmkzR38
tJQLsWXwg+yHpkSVf2P4PpzA1kOChFNEYaWiesdi2ovy3ZBuINYNku4hPX2L
mRQGTYNpRwruHh/fW6Gpitz4GZm/yxx7H33Lu5hL1Qk92qn/6DD2n6jzd3md
lPzU1dk6wJ5FxclDpuHoh9rEe96vPgEag1x3y8GGMbX9Hpf0GlCRzPVuAFLw
PXx8D39EBDmXueAskBdLTKuqLs/OPMbVPrlXJJIm3Lg7+wxkZL0zazCHnqk3
+X0jv1KT0eIVBNLX2EBbmJ0UAv8w3DSt2tH+mf1CAfelTNaJux1w8+eXrQeD
xEcS/oeNxcdJKDwJgVwLhNvEhZ9r6QMlje5p+6RgDjMCiRB9zZSRnUjskQ5i
xWF2DtPEhWcxwR9Nc0+WFLPCBB7Luz6mEcwNJ98WTSGtBfln7TGImkGe/3r9
hx44KQctOxFopT9lV4VwR3AIP6ugVXxXZDnFufYPsOQOhr1ohI0sh1OnApLD
puRsnXKr6IZdr2QXJoF3qtyvYQNujaD+nLyVjPvvAH7fYn5Hu119wuJKUnYI
pxTxeSqO0j5kUm/cHhuPVh5dMEQU8Xh91UHIHsuQWygJ3DcHmGsKyveBEusy
NLhqbajG+MWbViZI1uSX+hn4Z09HLE12y2WoMcPASYtP+uokYT3FkgJNxEfI
iLcuHZGwAXnsO2VqgbDHli8eitWVkXDdOmURzuPLOI6qPgahNNLLbGTvLyEO
qlA4dO32BOajUhYIGfK5t00PgS3dzXGerhOczbmGBZrglVw1ypJBDdk1duCr
xzFQ/1eSqGBz6eEPY6h6YRrUKl/fF6NlWsatkzudmq1CaW8AZAWz+2Sm+TXs
nERK94QbpIKJv2XhT1gKLQflU0Y2hij+WVo7x3sVR8jp1F85ctnScroVXTCx
7xOGwEJiJadRgFYbD2iZLNO3V+1CDkEYFdo44dNP8Itlpsnn+l/NBe06D0jE
tyTzZ+bGvqNmyWNbPpx6NcphkIaYf4fx8ZrCYgIvc0iZ3mlSFHKs4sk/HhkP
dhZ8H7LjQ/OJYk7dC9Yov3zvF3k+zrP5KmIh8Kw+f5lQuvPdLJvjgi4syLlM
+ZIwKn1NylCjz7x1qWWIgBoFRy50dD1UymoYGP+ujjeOejHBXKAcTNVnMIOw
7iKEwmKK43DNIDMt606EeIsg8Rmq/2uudnuCS9TcTj/L4tbWe2fFDQmlhnp7
tuSEXAWXgkFwwY8BCVWIZJBv5OYp5rd7EuNtEvkhUao0M4JHBPTO3JTqFTEP
+9UP5uaO53MMBt4pnG60hELAKi0cWn7kSwt223bg1JreQfWjYqGogp6Lzjuu
jjZv4g7IewYgwvlGcIGCX4kuxhhHQjzWxwDiuTBQn2bg9IS3RBM4Y9VYiCwm
tLUZ17YfHBcqh3OS7hOXQD75R6nhU0/+8e+Xcw8fXjRkbhMyJqfJ/GQZg4Gf
ih9abngGmtDME4xPpsYR98ba1uep6QiMxJxWLJaVVIiKUxMELwrUOOx+Xn8S
bKzuWGJHhJU19jxRTGBRqLNDfDnF2IIVyVCvyWKxxU0V0nMXHYv6LwwoM9d7
Yv24HXtTJFNweVPtnd6cByW43xmvNJVhYe4ZB0IMHlKQ0EFyeVVU/kpfdowr
+hUV39TyuW8XV5NgGuXsIpHXmhJivc939igJiGVOMKGc8QURiPKijGuWiDKG
79rVQXEbu976PqCa23ig2B22W2/He1w/HHEqqSM1btQpc4uJGRT+p7qvL0zW
h6f2T1p1+yZruNxl/z6b0B3fnQLkVP3CdF8V6yBQ36q4IMKDdbqAK2J1g2+H
g6aIXY6gltis0akO6x5bKXi3MNrZlkM8sKNBgq+3R5XhLz7DZMd8uvt6Q8pk
8xComsWNjNWq6A9nC6F8D7GMbmcm0cq5a7r0W9UGT8e0RNXIMS/61Bx4glsr
dTVnob8xKgvnN3OdjdAg3tFSoP8/Q0ucrbZu/U+XIlYfwbq7El1EdrmHFqSO
7zamNuXi8mS5sZN6PG01qH9y/D3p8PBi65/qeKl9++WnRBvXQbFSH+wspblG
gALhKSMgyclV7ULsMPEwspBbkHfnnztgCUkgNlv61nv3pha2+hf8FY0YaJx5
mhBtQsXbFqMMuxlWDzytHsxYpLDeiE3r4UtvdA0S4Wt68HXvNvDbVuugTY0M
I8CQeozriyvDnTHdABXYiWO39xYmGqzc4aKcsoHM7EdU0WPdkU941psOD+ke
n6zKPSu6btAAQv08Hi1ugKNAhnqB1GGIW4/K1CgZQ6ee7pq6VFuuN1wBODaZ
OjUk7CLWC+bbii7nam22uTDRC/4mKhReY/r9o+I4PMr6GSnjH1VYXLbfxgrP
OLYLFdMa4AVyNjKZa/QGZkv+GaIkMXkdz4o1GxhI2VKUputA5slPBT2txT3L
6o2/DVyVDGTnBK9jAZkI1Bf5brRVTcxxLztKyY6QIOqUVuGnD0EA5X9CwlWq
Gi+0uTIjw/rvvkKyCdYC5S0VQmrt5/61B5B812AlrZ8iFffhH+M+HsloPLu+
oHMFw+zG3YNziTDdnpJyDZnSD6fX3Yk9nq4DD5CQBA+0EkUtYHOAdjktfXcC
RFY48472k3LcoPRT8K6AKj82xIqq/tAVR23qwGFgLtu+38OVXlpbTI8Tl6CO
U75nOm6vsRjEAxDsKMx/MeH/2mpPEvM2vOrgKAIJ8QqKs57J7DHihkVioIiS
IRp65bV/b5fkFNKYdlckrvM5XCgg9+Xx+I53bJ94oo65YesElpt8OOaDccij
SYUsYCSEvh01C4UbgCkX61nEFylwi75PjJiElaSMdtsz0d6rZu0nBsshciVo
EBH6pRAHVQfDpL6eK0xRB9ul1bHnuEqhZp/WqDD/uwsgW3WPrlUUSCjT0yjK
hD0pYgMN8GTne40X8xBV56KWiOsoVEfFpNBsj5TI11HM0cxFVA43zmRcypVi
RhFWFgCKx+n+kr1mp8E0Bk+7rixMlRl+0BMY7mUPO6429XTepnWaMXg4kfHu
dFFbNKQCycEL4TQMtUhcwdYOTWhRv2BC6h60EDtzaEj/EgeMEJLMiQXUatZe
b9/xSCsCmSiecEncGujlhxT9Qlpi+SO4d90RrR5bm7xcx8oY4WEa6uyfFtxo
Sr9FvM2roRoWuHdu1kYziRY+vPmVJ7tFrNYmwYBzDqNs8evsT9b1wchTWQZS
60Q9KrEkGbQRyiM+jJtLuo3EhB5MtfhrJm3O/5PrT7xAJD+cM7sVKmzjhET4
/lFei3Nxs3wMkOiMT26f+UeS7zGgRAzrhLeyYJw8qRNsK6VMpcY0s8d3heYM
MrrvkQYmAge7EWAmutgTg2K0gPbjc+ft0xogmz0yWzS9rnlIU032sbWyX1tE
qQ0SmrI48q28VF/ijoaXpU6fCZF05PBpBmOQgjqVZbS3lABgwLa40YKq4Ss5
mtNmrDG7c7tWbZNomkRPnTd49Io44CrbUFCOPhZiZOtIAGrBKYrDYeKbrNgi
+2VJHmvAswfn/fJbcbWllJrfrs7y1Qn+jQZP2JRsIcBrx85ib/uqkW96jBlA
TNe5qMZHQc8Mxq751UaEAXiYtkoGmz+mENaS14JPsZIYuo4y5bWrj4uZCUsv
8JuJ66+4Sl+RERhEJcfeFCsuXHjrkDkEm0xMiaG71TDU3thkD4u3OxXQCeAN
ZK0w7GkECipPm7lqnQU7YnTU2ai/tsl6y7U11/0jbKcXzxJ5Ha/Vpq/XPG/w
nsSxBM23WZSJTaM0Z6t1BXYDI9vsIPms1Z0BCsCg30wcyRkHIwrCn2FMjY6z
uEpcbddhuHwpK1GTAIB7aRYpkQGFC2tYgWMTq0zbviy8N2uTbvIoMfRzO7cn
7Z+IVqCUFPH9/7+Y3SiIhkCqDm5r9eo04J/uh/Yx0SkhT3ropsyPyXz9SMcR
oSo6YUonqCWGQtrY0zz8eMJkcEjW03l8HWzOAU3c7sUG/635x7UWnBsmxBx9
ME3w7xG0ZgLTuE6h+8fQiCqz3WrdWU3LSPA4RM1TkYYraFhonIVFsP2jSX68
3Oyltaoft8MNwHKd5/OjfTFS64SnkRWBRk74TFAXGksQB+QMMSYynXAwXLk8
8vMqjbj1SIVKHtXgCx20A2Bm08u7EBBRGAXlG14n+0ULlZkeKsqHjBK2JN7j
vajRdNl/44EKdt40GG25EOeXXQ+rmwayzUoC+/KLYHs38SEig5GancnqcMi0
W8dcBUupPzH5bZ8JhCrxxL2aWPAIgdUq+8LjbEWqYyqziUYHu2bsbLEkXTEI
nVnV9RMMo4GxJ+9IW10Rn55acPWgARPlS8Lpac3N7zB97f+uC1s64O4L700G
6HBslu+azTZLxewBHWz0ZBb6n9DiZoO7IIPUpZ0QcRmedUgdcunJEOY+mQCK
mjBUIhCg6t5WAX/tdObmT2/qzlHNcWGPJh0P58zbmIlDzMC4j5ggZ2q9kqiA
uL2BSr/hciRy5Nyzhe0AmsmLg/80wm3B4Y+dbdmW1S97wGf2/juyod2wFv4r
D5hybTGvIVMjcNWWde4fdJBCdrVHN9K9cbAXlc+b+pMqqyicJwiURZoVgVnm
aiDEKCFxDuHhAtqWccyUFbs8r2HjnZVeatI8XWZztuhcXYJwnJghvW6zWkO9
u3ixQFXnn3+FLNQLopvZ5rKLxMbmfKI/rWXMdH3EmzrwiVdzedS3PcjwrRK7
b/fZxC6jrVDQL64ItpSkwzxEFWgAHgcvWYpAOtUQPsHw6zOBdB4L68Z6mbnK
q+OuETYJ3LdLlF30ikXh/XhlRWtAJiW02xenPWgUb4fcnuCgs19FnGdfIU3w
YbLFbNHNDB3Vv7B7unk3F1QWRbXSlOhT3hqeHtjKkWotw5iZMkZ8cdEPraWF
40JoZQe7gud9xqKK8dBSyadMMJuUBqlZSHLLdcCSUoaOzyc0WREI9Z2rJS0r
If/7+vTndABD3mHpnIDxmMRhDEFaFHsIPP9LfpYaB9CO+CgErfrFOXO9u9CQ
HsCNVZ5hoqpKnED7UmoPaclOO19KuZXLkDl3lfkLyLhnghmnCLNOD+VK2P5F
2S3wVVVeijzjYrtO+XjhDr5sjqd/iWxkvoiAIAMnbAS/QRd2aCaDFZD38aH+
e9RakMKh7OLGmEdCwb7F1GLPg7/QMfk7sdTanAWxyuPlN2g3JUZJ26Ca/d6e
RWqsXkkKJf5D1/pVmM5QUGA/2fWMH8wEO1EcI/MZEEsY7KgvgTneISWHzsDv
YTCD+4bR4fHR3k9Tt7afye303kSvDRjmgps4Of50BTYnd7caI9l6Jv/KHVFm
Fc3Go7Gruh0WcLvGkgNFWuvQqd4/KveU5BHkhmJheIYneb0u+hGVhNervYZM
0gEzCo+P2dnUfqk2Q9UE8RuBY6Q//jOviW5up7GoxckmET6FKYgrgw2MjY3e
pz3svFZfe14fmI1+vdPURMYaiAvoGj5N0G7sd45IgPjSaf4qizgcLpJ/Ie3o
J4F4C/hgqeBaFV/0VyG/uMkRW8TWAKQ2w7my707W6Oq90+pjIj1V5V24IdtK
omGGXFAUwVYZ/cFMJBJkt8Yr5G0qIwNEHqscYupvc0229iC6Pory9/RV1/Sp
RyMAO9BtE6pBKsxFWdpadXj53IoTUjiU+bj+73uLZBWA4jiEp0JNIrlsgsDD
Lf3rveRmC7N4P3JlKac5vtcebdl2QNuToYSoOqWcve3t/Om9EhWt+zma9uSU
txDJao/6RUem9qKYYWwsDIZjwcNn11NV8qlecPzakIcvCmSlQxCqXeh/JbC1
PNVEIOLZIC4aSw7dyfQ/X7Ovusflwdc=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG11LE/1qQFpOcNu4tst47Uct7UbTRTZeKtG4otbdQG21OJZDNFX61zo3wMsc0ZfS/yS3SeOFGGaT5Zehx8F8tcBtbBAai3ppZEUXJBZk1wLeeaKq2mSINTdJv+rfFAnInxUiHL6Q6C9y6AN4IQeyNdoEnrRyHrR1gN4ZSCVeBpyeDFiWFWzPofLKq6pQgb+Sb5L8RMD52QW/r2LiOIoM6gzV6LzcSMZh5lSaA63kZyPt34KhOXvHBASs5eX+gCstesCE3b7oPsWPtUTJXAhJTmbWyT8KRXOYByBxmHWclICpCg1RWucojoYbCfRw27hbSFdgA8T2zG0UosbDhaeVhC3qSKHq8iz6apQMn5LlVSETpIaw90zqQtf0u31zZ2Tg5w7nQiFbeB1MEi6nOxCwtFQn62QN3AtbQE9m9ge0dCbDRbsjmERNjRCD/092tJ/gO+x/J1weGj1sIrnENxMTNYFn1Xd5d+YapLs4RuYfsQg8aly/VP8HPqK+g3Waftb+e+SsEViSEcpwVyTJsvir/Bmk8VXC0mSC79KczTtUxLbDF+pmKLFG4LMNoN8F/4vecxy2kQv1Qmj61YblG2PvVqOYmPNw04sqSUaWfWnLhqrPbadcu6ZoKoyxbIBdO2IxOrzVpIsSjy/U9BGr0z+pwxj24CnPjEtJ7ZYlz4MzPu3zQzlokXHRfEGCeHIe/2epCYKHDIUp2xwBH9BMeMV0iNcFYYYhP8ZFsv4C0aPP31/kci8MPupdqt+3mepyoHCc4FbAqggrFxDWC2N6eBezy78"
`endif