// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
U28393XCM4+SnsNv0wcxFP2vQvNHqpwtF3G8wS+9JX7dqMx1yIjIk05f2iH8
UiiB/tQBboWVk6pH8Rsr8XGWgZLWvTE6pT0W2WYDF0lIf6/4UA56gl1BmbbS
4JaXzmy6w599iMs7N0EpD5fX8Uv0i+rAjW6NVoFRPq5cMnWc3maQNU85vMml
Dbb58P7HdE4XBWA6ZLMAzDmQ8hZWdletk720DrdN9YEsjS4xC/vZmnH65+5S
SHH7XuV9/Dl4VozgVWIWdTDwgFyietcVLr7hsowORvry6nlAzoiOtPkAGVhr
88VWaTwAnzB6wG4HSlFVfR7g+EscaEzCKkvtqn+2Kw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WKfqzw9Drd1u75R3Cp/ZENcAygsacsCQZiyuzDJ4F6lMe+/tctqdisqzUuxG
5pghA9k3t6RmgMiWd5Mwolx/e2C2Vwsw1/U/HjdqtB5FDebeISaxrmuF2qsa
3iDigEVMDtfnOVdA6TYV8atNGjujpWZLCr+50gSovS8BtlK7lRQHRGHC4bp1
FAfn7FpYBOZZj/6GcEpLClDmoVr3VuyWf3k+S1A8ShzBV7Aq7Y+snDuJFTCX
iTSnJPcMnUR0MBNXFVrW7o+P0R8rgSpxI0nUYTJ1X5+KCQSkmP90fO8aOX1m
EzriMyZUbBdZdRtBZIk353yT+CnHvaUu/q9PYN2c8A==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
N6kLezdWiQvqWnY15sq81T67NtpOx946lFG6KeNcHnRC2YQbO0HFo9zwDtUQ
KAWiowNPu8nYDAT53cK3l9jbA0ow81Un5xfc9aPRDPD01eA+4Xz2OvgftuSF
/HF4oyT1v9YseSXKFTLvpIR19jZHiQfZCuWediYqwh3sOVla8PqAaNbz7Z/O
0cxMdKm2K7TZcKtNlBL+XbHZ1sIoJGz8BAqgKYUJZcAbRbo2onvdGhOaRHPd
gcoVGCLxiWIVfnJUZFzCT1nNx4k5dRPhA+x+LKl2V69Wk81FU73w/4ht8dk+
vcm5nWf1qt3IqTg+moM22afvJd92H6lkzccqiyH43w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JjxB4/+3kmkhmXcJZWj9vj7bOcQ7ZqhJxh7pXXr9tv2Dxkn5LRAJJjKcWT+g
i9wYjA+C6vzvw0o7wdLAyLxSH8v2h/ePkvWzhHxwC81+uSwIfYRMxsJUZPap
nTJVvfE/77lL7e9im8UooMtwGx29VQs9sKlDIXlKG7JJYtLFv3s=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
OyNiCIVBlDM0zQj7HFP6yPg2HUjwv1Epp6sAKBiOS5VxDd/L1DMB8pTNZjk7
fIokAcbFiJ4sKrFclzKUuE9LqSaDL05UhJsHtTGaVPhg19rg5ko56qe7fPH2
jru32q9M8AKRk1T2iY2btyvjzWBXJDIPge/w6Z5fh/W3FH1tWCO6+Ma0lViW
fHyoIPITv+K8pOlWr2TOYz5ndT0k4tyyFJ4Fcm2JWf1fDBXFEWE8RYXpyh77
71k+yy2uMUN6mnfMRWzo6H/7UQ/JWp3Rhr4WaVoRr4nj/fZm6KRQlIsNwo9L
X5WXJL5xOfWjIRcug70JWXMVry++8opwaP6VJF/4DwS8A1clbEsBjdI3yNBX
h1wpDcgqHDDGik37FAGzAlWwNtLuRY+XMbnUpOFPlD66dEOAAdWONla98D9C
fXVcb2BuCpZOVfkeEV+9a4Ll0vxqwIZ+djpkGM/t38qH76oFKD14wbMHLfVn
pLUWv+amH3TY9sa6obMLRRcQ6cubrJXq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
hq15PMvR5YnfrlnHVJ2DYFu4iGsnlZEKCpcOOqaZhJ0Z78gJ26z1dvd2BoJb
J0aY5gcQH0NEJfAfVTEBqDEEha0l4xXZIPMPUykqFtz4J4aHi7Yi1vEZnrFS
bAIHPFpG3CG26ByARjH5kE3OtVpQ9bclIQO1sOFt48t+QrZS+hU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
B28nwKe57SQm44AUjTDevYNTT7jxaxkNBH0upBQEydDeuF6SSrAIbqFJTT7C
Yqdlx7Y7osvKvDdbOU6cJj+r47m3nNM14yugckI9zJSfYYbzhNOMHx2eCCE7
mbUC0tG3pCAPQeLNr2bgznjoMPNuk8g1yYmzZdG6Ncpwh4e0eLI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 26752)
`pragma protect data_block
/1Ji/LswZF1YwWwxckBHJ5GMw373Q89idi0AcYbgYr71dM8kQynhEPzSw7f3
KW6Ky8tcLfbocmM1/nOqfq/S1Pp8NR91XaUlh97ETTA33rlMCaWauP6qJ2s+
M0uJI1dwFRqUMNhv6Agtmoqt0qJArEgTk5hjMN93UuAdjHfrF0oWOVseI43L
uezjkcPmIOc0OonuwbrkUjbVsapkh24X5UvkTN+M3GObstQ12KyCZDim8eCG
Byq+nT9yYxl9P30IQX2pgFFALPGMhY6jplKZH7vGUYUCIWtBLw9cDqRPdDAj
rTSWx4MZtB6WlJBpkCR4qt6XxNCjReGFqZUmpOPVoUgnswmLhieV+8bYs8lB
gkrNVlAkBIz/NUCxvz3fjirLtNC79i/efPMTvHFrtJ0qXcaivCBwDI1jgZXv
g9homMef/YZ2Ah640GY0bQbJ54qCN7TysT4a6qkMZ7MiJ1fzqbZFBp0kCYOh
kkHdp+pzkXstn6DfRd4u63n2hYXRCVMJ0dU+KfqydOM9YVgfGuDUmmBMKLw1
Jh7JBOfwvL1HW63xXvL9Yh+xp5Pa0pJglIuwSuCjM1HqhevUpHYTdTATu+LI
BhNCeyDuk5QHZBI/WctyG1CJT0T6xfyVPj1NrmmbDf/4IFZdWBiYQUCjqRSx
Eae6Aw8aYbIms7BpHXjvbYgdoRZ55dio5eOVuJ9s8pzFa0Dw2TGirAE4lYzC
vqOrtkFr0/meBkFvEx9GJdd2rTUi8rU5ssNPgcXAAPXc7lsr+1tuz0B5gDoZ
6J5GvSXW84/jECZyBcr0goD2jYlral41qnnPgUW78+UrmjB0Kw9d9Lf6/I9w
4xZXcErWCJub96N0GUbOdh7DWeDU4lUj0/zaaoewiZ3aXnWBrOPS5lSCV/v0
vI8n4Oxfy64Bh/RsAx+uKBFAnKi4E31s6ZF6YFrLVmYG909B4FoKlCzPHi8m
QctjklzazgXiZxj6MXfST3TeCwbB7pGgha/JAYge1UnTr6DnXQv2RKyQndEE
dxPuQSQTRC+HHvVTKCM3X7nWqc5m1o46m9/JLyFPh9hpBiCe80VZqQ5K+ONu
bG/io/kYRibH+4zJi+WT1/Xbqljz2B0LMX91pc0pzTDQ7ZsyeIMagPXFJuWb
DviBKcqirQmFR++nVu/N7cgd9diXSZ/kGWa8rEsMo2Iel3rwNLhRrfJVLdyc
M42R9rj7hpGMZ0nHgEmz0s8KzB2H7q5+++cHxzwdh28t7rtMIJOELpxnGbRW
ZvORrb4tlehkel0ghTdA4pQ0mFcA7Zz1HkDeKsV5rz4TXEdFI/9Sf6IrCG5M
oFGibEIAxsqtOWGkbDycLkkqsC8EgLgS1l6BUB5DsBNn9IJfIMTE0sBwk0M3
dQ4A4p80CK6s5Z/NhcqAP5ti2bp6j7JHsa64aF4GHknp30UqrdDpuV66qX4o
yXFhtorlOFa8npkDbFhLjgJLmguNfdQbJkCmOGDcxCkVqZxr04bkeGh5xz0a
eYRYwjD9J1BdKd7xsIKBsaEn8hNFSLKQZbhtE+TxoNxqBGobkrfoM1Z0VFNS
dodplezhwuC1GtUafQC9yBPs/+uu+7W9NU4x292YxiRJwApeD1+Jkj60e3MH
CVdgN8ZfmuEowZu6Qfs8Qq3978HTQtvRw0WXvYK2QXPXjpkPKjxYKlaq1sV1
pULwIy410NwEUyxt3fJ+TYo2mdWhf0dt62UM9L5ZGex86W36RBQQVVKG/QHg
snJjMi8qs89ldg666+C4vNXAc95+zsF4qvh8Y4XJt1DyNJC0yeG7p9xbpAVM
Gab95bGdRVlf7rg6mS4lfwWcYOdN3qjH9+Y24vGvjeZPS5Oj1y3XwCkjeJ5v
skPxC89TsllN4K+TkPQTH8dDulDA3Mmeuj1Sf1l4msGYMF/UsbeApK52aK3t
zqKDK9Ctv/6XANS2YQWvRXe09t526/2wWZ3gnFmJGX/dpamv3zd1g2X8n5TS
3z2C0Etyt7CO3+mNj8GvBB3kUMTa9nE3Jm/8z0VhLDsJSg17fQyOfN4IH0Jh
Lk71+MRqL9XixPDXuAngbNHATK0W3ACqPhAC3s8UuLXGPWtS0PnSErGVGI/9
sEW5yy+kZHQxJaLfWSbta1X3Njt8/C5k7X0v8F9ycU+tCLO1dkJBDoslBVcT
ds+QNMV+l4LDcU5+ZBkZyaPWenyjfxh1FlqjPvv8kE3MGFkEmWlAT3XDH+dw
ZbPUcaZFYGwanTV3Zdw+wTOvtJ0fkQshlXFQ0xPzMbL0irQiGh6DYUh1eb7k
LlAR8X/UIBxwTuX2MlIvFk099QjKabg1IptX5ESdb65geW7Q5ftRPmw5E4kX
OKm0jdNqS2Ta+/cUwk7w/r7GYD+pf5QIw5eiIlCHP+55Mn3T0bMe1bMZNnTX
FXNxXdu6Uoerw2BcCHvB+wO0mJjTx6LoBAQ02INKyQmkiG9NLz54rrm2/RKy
GjgdubDDRZSF2Tx4HCQMG5cV4+Dq9OJwcpAxhvnjDi9Ayfpm7cXQNHr08bO7
yQzYXy9N4j9FmVzZYTmbzAT4UZRIBQKIHEWuKNn1KgSRqLeITkW4nyUTbPne
OtA95TPv53FhAqKF4B+EjdE/LlnTtP4YNDK1PtBBS/S2eJhfD0+XpMPKCHLe
zj8bSB/DmUxV5TKxZhNGpKH20Jb2uLwtmcZ2jfcSLXhoP3BKl5FfRjVr3O2X
qTnF01S65bOWsV+ByKDnjE8g1+IXE+Ph4NpgUvkqN2lFcsx8GguTdSfYlWj+
P2I5QMglXcxuX+JnSvmDtG5jkAOXnxa65LL8bPkAzLfHBaWgwPkC2SDpsQyh
i8bggpsd6axZvy0GMKaokGkMfkom6GtmvDHA9qoQgTP2b7+gqarCmnI+/kmj
Bb0MajQFwYuIWV2mSM/ksZVIaav2wfVWUZitbmWUHuWZHqWYE+73hNBM4w5X
2MYpau3GCp2djtfJKq5orqCN3RIm0GSe4iVxpae/EDUpemDd/u69KCKq8GsD
Dj6iZjk0wpNLA9n+aNLo2ih9RsHx+Q3LdJdejSQMJZ2VCDtmnsulN7GqDr+4
AdShl3+u6DZMDkQSWKt2Aw0TdJosd0pxzibMP5Thyc6Oje5MFfWbm/3UtXo0
FXf13Nh9dPlFHekqhq8TLOuyB4b+MXT/8RDIu0KjmuRClAbF3y8FvsVkPCsB
wiBFQsbTQP1ViOjpCqVE2SkctkJDtduSibPZnqMy2ALz84sa5BHmfBLT0S4u
FmElwUQTojK0cczOXOa5s3CwSL4vI0d32UFzRdhNHCS7WJyxDxgrLsFrDlT3
b5/6iTfxs3rg5eRcP4t0BlMuifETrMjyBnxwA6EDvmQhUSMaKV/oejCMFN6T
9R0UduRbg5q+S9fg6WKCP2x5u1s5wqMaNeYEDhoBC9c63HSPRZ1KYXK64Lhr
/JvU54SYCdJQ+Zv4f7zKAG2RUS1BYd7kwecxx0PWfwSVkvXSKbQvPvnIBh+n
tWiXeCI3mau0li6LiUGSviXiRlPmh2UPuN00XEuNgvPDxWwmYDy2aEbqxNeA
uxRJRLAYodub0Ax+JDjqvJr/KnWJvtD4D6DL8U+DruIfuU6diXkZb0oKykEF
0bcocuXMJ106yUdcP8Ue64ASPw3FCL8y/+Hrgke4bSk9VYMgkOWOKGFUhmkR
UQU5NTdhRaNnD3m5Iv3t5xD5UitNDjygEqCePZ2FZEux25rtUCR7MJs0Q5zq
gEBLYn4DYO+N6CDa4E9/FGvqyDiKLCllsOv4un2NUT+nN3JmqqBo9jouWxkj
UoNFB7ek0u5/xpT1KPD3z+P9RSHSRVYWvcfTZUaA3IgsTA3g1v/V4z0DDzyV
FKbO+0n5QGi0XE3ignGjYCXZ182/LYaOo237jrBX7TbwY6w5xhHlhaNmKq4S
JNqIkErQ34GxrTkpkQvmMN+OaKzW4nJHKMWbsRob317x0iztFSyftbJhtynn
LXP/3IYj8IrMKvqozjCohYfpoL+jgkQFvi3PH3eTDM82wGb/HqSqw/n/tupJ
fqFN2ODObibykPZU/QXyZIEIQEOKBfM8VQOwyWYOhMtGKONjnsbRGpiKEqXW
emdxnsp5eTz4c74Lx8naPXpK/CqHj3t8EnUjgWxM5iFVAjbtFeOrw7dQspWi
4Shq4a++QHMxCZBKLgAURGBC/kesRTAuLJeU3l0XvTKqiHAI/gq2M7+PouOL
BExw5WPUibzff6lXsYhLj6rzRbDlSNi/4J0WJGOf2Y9bazetPE6BIEoISSaG
0kDUnj8tbGGiFvF1f3xhfkzaaTES5+kpdBsywziswIFTj4azTmeJQlbaNYuG
CI7xMrHzTtBoqYU7G3atLslhrS6t4MmJvaCv1gyuhTMh11qW8RFupXaeGzUW
JyJxo0yPTOXWCk0zHFwxfrb6NSHS5TLlStdQLsUBiDjEiI/B+MbvV5+h0UtU
8guMEwvGNsBwQNp4JkiBBeFFT53Cbq/4sFalhYGFyU9eMzfNMGzC2jnE1WkD
PnY3LmiJm/n6dRSupMIhkTGnghrD3MkSSeMGJXZbjSUzDc7RvuWNcUU1eNNF
1Bp/fA7putqC56Jj7cjz6+NB7aiysklYBewNZT5WbWbLy4wZOQ60NCHvgX2p
PkcOELD4vX/1d6PE7cG6M4IpreHpI/yfPfjWUi/CcE1xlT4Z4XEuHvvYWJC1
MCe3Sb1Zw9/K0OZJdxESM2FJBZa4Bt0g/l5mVvUG1n8VMLamCmhmFhLfRLLB
r+dI+CASJjuoGQFThZyni8JHIQGLsSuZcwhWplEd3FppNk8+ydfDe179pCwu
Zhlor9PHcBVMBBMKma3lOK9yRAgYC8TtWuiXoV//BEi9ip8V1FPsxgpoKm8o
bQJk08fNoplbomjLxy085O9gGWYo6Jyw7K/PUTQNJjFIs2zqaX6UjssBsnJk
bss61eZtoaGgTtLHLwqCMY80Gu9MTvKmF7gusR24Pq5yU2f8BB4OQ5qxzTmm
jwTzsQqTrE0CBokEqYHZlxZcFgOLofoU4bxTnlSdgs8QaJMUnuUhc05NUN78
6pDE14/Bai1LWbFm5NTApz7Q3Z8GlO3i8qtZ+e8SyfnY6As12OYYks0YmnTf
4TCiwRbP7RS8aXsfz/+N9dItiR3IsJHKCIDymndSYDKID9KWdYgRWthuUpol
b+zqW/GlbxVAICjf90VF/fZ3x767Tyv8J5ONciBA+FxvBanJPTsRxxJ1f9c2
co8P6C2TozdtcUz5NUH+Hxeku5IezYFZgg7pBh3nEarR+RPbPr9NXmI8WJDT
lorJoZrD5QVV/0+rfbXTS3MYLF4K5C3AAk5ptrI/u6dcK4Z3Trtl08dQkwZi
WZuI0cijQKNDkt1T8zR0yrSEYfX1019WpBwSF6NgcUjJ7f36fo2M8PqZ0MkD
N3G0vVYsAgQ1TVy04ZByFOHA67yWE5VFbZruS+03HKOMBXPdB0sb7zQUOx0y
6AEkqm/gs6NLMDyFDnIlmDFyVNjokKrx5ubqL21rNDXsqcb6SGpYdd7Vw4HM
7fs8Dc0dw2pN3CXNWCdl+kFIyZe/iExdHiw9SVVbxjPpyQ99OZhiGlFYvoWu
dNMSNiusEoOKD1acilAlXAAXLTX5yyWmIqTVInC38eJnov5TJUQNa3exRhMX
Mry9Vk+bSVyH9IPVX9X1+z88J66/PUYb5Fo6cAWpNNAZ9ektYmWInpXFdnfd
4wEO1V/A4iqZWO2ilqnrI5TOFg9GpHO1ij2XhRLKDffEuvUz++0vJUr8dRb+
gS+at+IRzel58EMxO3CNWxl48XiYXj+BNNz+3BD6IvNFei+DtapNQRc1B1Vx
YuQdoZPKCBU8zOeobqfXFIUYlTKuv/3JcurXkIAaTA23R3NIkdEVhJL1EtAF
G5SAk/rRTQRbDVbRsnDCLN5oADAgV9cBj8cwHFRYN+dKKmXCLfh8atPSwPKs
ef4cf4/mTnaKgTGz4IGWNGVy6N5s7/mb+0gQy+rf2N3BmS6PDr34RKjN7Gee
Tb8Ud/s38TrzUO9tm7LwS8EMgE2GCZ3RigvMd19RLVgw0AfurXmkwNrIpaz0
e9QffD/ZBbhRmgRQQrgG7+RWVf6PVYiCRF6ZrPs5NGZ+74zkdCbZBtcKanmv
VjQlDnEjSRslkD8gSEv7hdFi24T4PUjYE6sEVHNv37FC7na4MvbT82cLE4rS
fbc5kGS51/DfpaO2z2ctEul5SveAznp55BoFgZ27McN2FHQnSV82bSY69LFS
zPCQZXtjPiSnAsw8G2Gv0LB35rnsRZK4cDl5FVP9nnMZQO87q5s8zN6zEpby
kKjMU6qp6HTz9fqt8l0A/XOvzBZcLzbH/R1JGZWKEKcEaCIXKiILEuz3hRiA
PI7pyFErqjZMXapR0j9hEl8OG1r7hcWkyPtPY+Z6XobXPChJEQI/ZmOoSFR0
XvEXQ9IV75V1y+4Hp1cpPiKjTes0tfqbPnQXk87wvkXKL3O6vcI1XkruqKLC
jwZXP7MyuHq4OL1VMwWKEQLfBJXX2EithT3wnosNTcWAwQ2m/YPwWfO08+1U
JodwbuIIJOqtUDsZ/7CsoUHeIRm6VDz1ovsjGCyA4+mzpvPjfLxZDSnR+/8h
bj7pQUJT7SbE3C+gZ4QmoYvOMqPVsT1NHpMmgC7giTovtW4CI0a9lUmpPqHK
6GobNjx0V2K60UOcZ57zC2zUlZ9p0Gckzr5N+VUs69O6nnQKhPXwtTGr/zQ+
XtX/NxxIRa5qhc4jDmLmmUP9JwhGYS+gyZRGv/XAftJcUhEMXGsqreR6XZ5k
gYduFINV8kfNbKo2i1l7Y12y7WUqTCkEvyNVtx97nhYceVaevywpG1pTKPCi
TQ4d6LRwUyiVGKuVU3RRBsb9y/QRjZ/fXhc4ttQdnXLmlUP+S9ez9YZP9ZUW
Yj+TKyowBcGLYinJ3YGui19a8smStOcyT8LgSd5fmZgwvVEigi6vRCO17r9U
UTdbSBa7We6H5peErG86KYvroYXZGt30Q3Kbt+EF//LQqW0N0rI1m4Zs8QXl
3eimkhZOyvuKeS4mL7UjPb+th3Rgg4eN3St5kq20DmuiW2x6P6w4sDgY1pWV
zomlXKXw3ks4xb3WmPWCviRQqbZelavZtq7ZEC3l8B4WF/8fgGEJxLCood23
+E6lOCwOBUGxJrFcixU6Wy/uScpISdXJzwtqgT/p2h1vHzZo5jTfEh5IE0Cr
Rn3SvDqXcjrqCjJTFEQZeyVHxa3cseB0hHH6O4NTSppJYC9ZmXeFKBv7CJJG
+Ad0i597OcBi3a37wAeMKhUpOADGiDlk60GH2tLj9SGxhEWN5YDb5pVx/xE4
WnOs97tPaUVr/BZG233bzKTcagSuEmeiNCyu9h6piEir14ndygn36AO/1/yp
oX5ttuCfBCebkCdGd7A7M63ZizKE1xTBZ7S6zOIWikb3Z7B9QfObqFWM0jzY
u+xBQd4QPzftxJ+e9PoiRqgzoq799aY+Mel/SLStncGjaDnhdIr2aAbaIkYV
teyAzB1JQWCGWw+7d/efYPhSHR/aFBga6XG2V6xQjjhX9wNQsVmbruU3A2LP
n1ZFVfosQAqXaXFO8D/MiFnJjHUm7iph2DqUk1cqu5qPrYaucUcgC/G79S4f
ol7158977WtuULuL9lNrXL0uieJ1BecD85wfwu9T3lPzmQwLflUnEq6OSvfm
a9P+GmYiLAX9vgmPzIp1Ze3ljPwmx5eYDdkyhwJF7+KeBsZjTEVAnviyq4H0
krGEo4L8dQa/28JKpcDns+cL9GTdxUe04G5tikIGq0SPELPvxL+Ir/2dPl4e
R0LYPxWi7YGQ6Yile5rf7FHHTpLhSOXrskH0ZlXUS9Siiieec0BS41b9hMCp
xpntxH0wDrf7nmR3jVExpdt4PNS/+XZFKNPx0e1YKDgQa+hrNpDBQN/id2uo
aAXVunCmKd571gAEYu8J55lWLfu+ooS52dpeQRE37i8jt6B17MWPX4feO8D7
dJvwaYRnfF9D5SbLOZ0gUlJgjVjN9scCOCU+Dm73QpOCWksyfsKkXR0ZPr2R
VCTiI3Jm9fhQSXeiPzEd611hDyMMzcDylQlZtM80OHa6FMxcFK9I8ELcKa7j
FvxU7AOH1cNazUKnsV4pGw4Ep/INKNHgsDJr80bW7mAMMledSYx4ERyd2pcz
XB80mFQj0HeWDyxfN+DH7YNgUApnRE1ed5Vu3KK6NTZiDUEDS5BPIzvwWB+8
g67XkzVK5zZm9W92t37T3Gkomd9m2X7+5EKjw1ioqGrYHMr2m1VCD0MkPdp0
kRO8zzWNlnt6l/JYncW3yUSppsmBkFeZVaGKcCniVkw1nD6f10aroTnkXfkx
3aYTO8Oov7Cij3vbh8vO2AFCEDUGbp3avhtRazd9SshH2RpjbgJQMf1ZbvOq
4KhnmtJtmr9rjisjSaOpyDHIsdFTNpH6YwgI+od2TBI93s7wMfAb5nHs95Yu
O4M8ncsxZdTx1o/kV/Dd5XRHZlzFAKlxyDnmIZwz9AuwAXD50ee47Cjp5imG
FPWvS4K5Qw9ksQxmZfuuHfFDZOFrnUKGIh382HXKq6z/GY/76HsBSVX5bRKY
C//oInFSaSf2IcKWyucvORJy11YvmSbhfqJCqJ/TSI8wG+vUKhmkmKidqVOM
peubD5g10TriIlVs0Tac8i3NaOlj2xym4MeuJ7peq3ALZR/m002DBZGMckbi
Z0il47dfZIUIyrJ7AFdDWKC17ND9hIj1fA2c2NwQNsLyRC+4YxqwtHGDvM/E
jwUQfMOcnPeyXcu5Gpx86jgggBqFCaT9HHNPqvNP+D7PdkpvAxHoqgsfE4ME
4Ld+cD60uLyWrBbuzRMbo56iRYFG3e1ke/wQqg6AqD1eBP/1NeXZ8+7JrY9i
GlQcUlJMgBzgOmSvLB+5AjpUqj4V7NN70touBXXfOfE6IZCZHwSco8pqiCa+
PTqMg4a6HmBMcG52qPGdnO0zmR2IAgLey5KK4yT2xHL6fRuC8ZYZOJwjHfi9
802+D7x/J19gRkjACGM/xMCZRM9/iRn+jQlKm1gNxnGPny6WWMAzGlZ0PBgw
61ot01dRpfz5bJUsfmLuOssGmQnQJTuhPaGUDYBKQAg5WY4tD/GXuirlxpl2
B187NhQH3xkMYWyPfdENlZK2ugRU5lB6+P2tYc2GNGzzLfClQDcU4EoMrYGW
8ZxmwVbUEHjwOaQz3GrHiA4EfIvSir0+omFzQHZxO2fIl7XiqdqoWMeJMA4V
Z74W4siXSVwRp1u1uAtp2zNi9qI0MkSlLzSOzEwkQK+05X2+djX/7yTiY2OZ
Ge2ZRx4cC53CrV41TD/eXBMZCEIRfumSL5RWLuQLnfGaXYapXoA0mswYRHxT
iOeHS1QL6DaC4UtN1VBgmlLfcubkP/zvRs1rTh9MYNO2NXzIWWuiI0cW+NhW
1EoiXmdt1M4w4CTmGid5wHDwOTr8caDUz+HogbTZQro2w+wrdb38yy/tEwlP
Hzy4wNVHBxQ/9DM+sKHp1D8PyZot9TOa8QiwZN3fLyQus6j4uDG3KyKp/jKN
E89R49u6LbafU8usKdNVQhMMpll40YFcUAqaXyDzJ7mdPMkn5dUV96T5JLsa
uxIGbskRBTbX7NqL6IEHY0dK9+EUMN6cjQfHBCEMO6Ttx/vp8mhrUplFmFjM
IVRY1CPjl9tD5EPj3ogi1MkqyqtdVPVMBP5+3kYMwje7bp3nSMWAdEa/dgvW
npwQitMzun3qiVqt47atsQGG1VsjNW6WQ3OXBvcYfoklo49phXqdxg5rih+m
EMmSfChglFbOSpFmyWjsSsaSgLZ6ZvN4cl0EQ7G/dZkuajM8P2cdbEO2VIRJ
MKCMwGi9doCmVmb7fRICPXqCXQGRS2/7WGqL5fyvjjaUUtPaMm6HBubcWDSp
JsBiV8jd8mS7GKVenxRgkwuFy65oxMVaZcSRVYbIfaBCc1WlUmjHRl5FFJym
jrLm6tqnN85CAmXPKcXlLLXQdCjVHa9pOyCQSrJoSgGDBDYNEfdI4QJ3xmzl
pmRYMdt/z5rYGAhRyTo6CV9oQsfOoUN1RC5E5v+tFuaPmiCKCeiI29wOllGw
KwMGOEG1ucEZvOuWM+bW67D/XbdLeH9MH02nGP71wKF8DNOZrnUYSQS61WOv
OLZgDgb79s8/e1anmXH2yVbE5hwnCZaJHvMKjfDFoWfphUkthHOxuyj17zb3
7/twlCzS7goW4l2MVYVo6IZ9mR6XAC7s0F/5tv4RVw4uLhTGt/81BOIrwk+Q
wtuP5hQ9ApL5CCurXmhyeJIwe3wm/xPSMlDHB0uB3CvtdqO5UFihNtXBxmhP
5ODz1mg03RyZOAVeyZOzSEBiOXYE10qYYW1xaaVuWhKtPT9Fh46d0Blg33cw
nElKxuJBzE1uvJR7HO4mLT+9EcdPXzg/YTRUCX81QLE1pMRX2c+ClvWGQPxd
K/R7HJ16O4p/Y66hu8KfRk+weRy+RW3mjVK9Hkf6sJyj68EnU3spLj3pP3c4
JZB7Jyo6mo5txrvoeR38t1nsKPKwrgVDwuFvTfVIzlyNIrJfKzlPD832x35n
gGL/FoNXJpcteoMhJpz99f6Gue2NUdy8QwunfCwaHioGrcP2Xe0M8XY/QCnR
FNtk5jhMA5r3xpIrgcMsnin3vUNjdNmeVcmwjmyM/nNsRhVpSKTnfGBnEfCX
2rZg7cu27jOi7R4s4tdv8alyyPnVBMoZ21HjAT5gBrBOkbGumE/+R65mMPdz
P8BbTsr3d9wjYkfGXDIMCuRS7oPrCqM34snCcWu1FHIc9U2ZcV9VgY5ag9q3
LjkD5n8QILUtlihX4xhjerWq/we0yPVS8l6wIP9gxQgLRgww8oOOb5LYlC24
E+pQ112y7+WoluZV2CfHLL5qFn1Q3EiKkRwvMdzdkQccEsBT08qsF1+lbPI6
cPDKid9FVLHt9L/cy02Vlbh8ITUpge1glhVuHHe8ml8kFxNpDmE0jpo47xrx
fwTvhnCxDN2P9Z/a1SSNNbJcmdu4FHoyxSpLGyDxWEf4/snwi3M10bZtUlQ+
pAI1a9RmX9by3U0He5ZFqRJeCx6HlvSr37dF0xGnkQIeVGc1n1G/aGxkpMsB
j70H3jnoYBqd7HvlR6yWVaUc0LT0LYkn2obuf6YL46i3kzfAnyITHN1Fhkp3
7FYlPi0xUO3BtjZPjM6XrOWZgVwNCD67geZAZQSr4YYrwrzf+2swHFZ2hoAa
TuYLq+6ox46mRLJBNAKq/xOes2Io0YqLUNz85+/L+SUjK7orpL/+xHS59YIw
T1DpX5tbyZUfHDUagtl2kNK2xv62FD686W2Gw9TIzFTAFrPApEKAcZONJ+f4
rr9Yr2DxudCxG399p5Eq4J5g0f5FVxNmkcqo4y4aBPdeL7UK5iQGkjwnqR3g
vn8PheHuB03A+7xNenpiyRcDMLqvvlyf5HHdFSi/MnUQ8oI37ky+5ld3buym
7v+YH/0ExTq6vh0R5x9Us42LZWAzUy1idZwT4cTimylUKeMPsH5VuKpXoYCP
yHpmnk2gy2uUtogCKIgN015lKG5SPmtEnCNcZulhBVHjuedB/6F5SplJzQcR
CmmgMx4UowGeHaiXnWcRR8xKzs+Ya689Y6o2jxBAYOin1Z7Ds47sfZW6UIOb
2QjAL8AsRcW9u/FOqfjHHnD/Lt7ce8ZxfSAcy9Vnbs7PpY3CaHi+LIws2hAS
/43n3TM8eFllW58bhEKxjjG4gKeKXB6kJp8Jfnx/MMRWdJwJfDk6/HgDV8Lo
ftK6Heh50djRCBKdkp0S4QQpesC2K907wDADuHmfMSY2TdwUxpDzxmDYrTt2
hmKaAa7knG54XPmzDEMs63i7P/Jn7D5w3YpayJ8QfX+oeIejOKaLxAPmNmWj
Vyjt2oa048hJSBJRX3iwIEySrYB4XMMcYJrRlnvJmsPhD9Yw+7qcuwl4IZsJ
mNeyLLJ5WO+mx2YcIOZl6+keR6kCLRMOq/hPsPtxljfkUfBU5LS9imD980M4
ljSNjuRe1Sql7CZ34D03riF/xiqQ4P/Nt7h4ZUtD+7fu7SYFkNhazVNoBDmT
ljX2w6pjNQ2AJfspaMdrykr+0jEnUbAgEadmX92PSasJM9j1dtwQSdRljkfg
vjoTXWJvotFA+ehPRYXFh8JSDnl6bml6EtBNWL1lp8nSqacOesJWOsB2/98v
8QwlnP7zppaf6jhW7fECqP+VoaRoyJ8mCOCtQn+CXYgq/8fjGe28+OmsErE/
Q1Ci+4v8LVod9joyHfni1xiCJKDINXbW3c0yBK9+QbSlibdnmAQDrQJc3DSJ
BM1zuUnT+zIKUJTv9RXctTDDUp4QvfO9CDSlJHEFDUPpWRXJF+l/1QVC0A8r
IQrKsWRahleqGHbikFDxAMPJH+e/WVWH1CS9H3To1vdjmJRb1ecOF/Wvqbpg
3+KMORkCZijXC7EOvzEockuej1J+4JDYuxY8LihpyN0CRASKpEa9pDOoAxWu
W7ZPbCF6l9djVvhY269Ci+4jWXcfI3ZZ4e8nH0+Ga3XCk0UDT+W/FhNNTTQc
q7Z3sc3ts34aAbWvDyvsA/2iNn1hZW++KNUiZMo0xm0FE894Y2qOoMHKi6NQ
93ulu0v+/CuWsEaUdxI4h9LFKdZkjHV0Tt4qvXukP++eVUlD+6nEX2CFEB9+
lSH0QnWztMF9GcYShNeY7top7Ol9/TOSdf1D++U67FS5Jfj9VcOTJe+4yZKN
S6xF9eQ4sZGi5K+vheIZT58fwUdxMBxockUcxEoNj6ZTVW4izPFEIYD07mKt
BZFXb7SDJQqRNKMCHXPCkDigmlMUPefbVfSklnUPY5ZpcagkKHy6OpTSrAY6
Pwj0aFYmfpBQuFc35K4etmjgQaS+lcNjqVlQ/9cCfSH/2lCfQDq1hyPdrxcZ
PBuE9fdVjTws+eX0Qg4ljHAdxLh88DI8ETOygIppDsAiA1IidlcpYv4jXtFb
v7l+s+aGNi2dAlFs5Nytf/U7Ioc+Rsb63koWzZYzCE6/f38kXenZb289poml
pY6EF0Riebx/wz9rCWMWKyiPOOh4hOkH1Tpa0P55uBoVRTl9UMhdkvUbv+fM
xzkGN89GUcrFpI92fqX4KkPUnZVAQNjkRRKVxbvMxrgYIP0wNT5xr4NOwPO7
ncsoKQ0WHheN8HT70X3WWE+9lE8cedGdsjHLNGZLK69CIroXqR++Kn5Vyq5H
5UN42JZ3Prltse+oUNkC7iewzvhDJS3KIs+cLhMi9QDM3W3/riHLH6Azi8oj
9+dHnxSH/9tfXJmVf7HJfr2/b/eOtVo2B+HEAoiKFz+XSIfQA2Mn7kO5Ap0W
S45a2Fa8G1dG4oTk8hYasXWsY69fbbnfoRq/X1EnK3PUHaRVOBfoOan1r39v
oOQrpT5sQ6azYeqiLs3F0fNSkzN5WyCsDGvt2+kkn9LudKhN/+39JczBG1EN
Tr4TrcchGFtr45K3Bja1cVKpnNkUBfmIRUn2pBfv7GiI/Rd3UnKl30e99CAi
A5wGDC9TSA6fwAN1ctCFAIBWvyPgRlTT5ToXEr1hdkbk8oi1TtGNja7kjl2B
CRuiecJPkCFw67YMBARK/ZBKxsoInb0hkVFvnfhxYCnO5sDH77I48juU6Fop
3LRul5EMtJ2nDZKx7lIq00ET7jeoBleInk8cVvHPLpCA2XOSHA/VwnrtcTmw
BB8k7LeVU8bzFlPvq5ky4f3rN6WWnARKAI/uXChkZsyTU9soyg9aRu/Yd5wC
XDLDPxTsT7A7xVEg4EZyvdn3LoK05z3xEeVJF5qIMAY+O9O+nDh6RVYw+G3k
7XxbbkLz95cK/qFXxkihmascnWjM6IuGPZ+FyN+36GZvqVCQPHEZ1vXs8eN7
UZbGMAeMNAXVycX/ipj9XBMQxdBQ+WTcnJA9cc/JVqEAe+J5qXGJIceLq1aA
sm5ZxFqDiWQUI8yZIHBMXf/lD3DcXtsh5I+BszoAh8/1QqNij+wa/j2tTe12
thWXA1ub4Yh++cTNlzpv3WX8Au5kP1e2UQ2LGfRmh4EE6Zr4vpnmPAt7mhHL
wwcfwvKUZa0OfisDLlmrdck5AJgINqbsrn8or1ReZSzQ+0jRHUOaKgBIBJe8
xZpnkk8pZyEdQ4Yt+U4odoAonbltYcHEq3kIaGlusQFNNf56g2S40oxPZ88E
xvmqcvSMAtESkRlnFOjMyEf9+qIeJ0TwQoHEfNmF7It2rFPR5/yYgZj3fkA6
iqLG/uh6fEO8e5mbtVzkU/L9U0iovOgJMRUZrl+ApS2Fg8aagLTVYOnMb+fg
yFRcj6Us+Ogvh5osXbWq044EF/iQkeeHjpL+vkY/LUxt8n7EwQXjK2aWQazx
7ExzBqLL7yBXyf1ql+6T+uIUmrYQgKBufp/+iWy7CA9AFCbB/TH5nxXVOngN
fWLjA48hYxUANh9qWoXjUsycFWgHSRfutBjI63s3mV+I68fy1rjmig+KPDWv
/aUTe2GUgNPyp/IK2YFcJNwQmOYyTmhxlebr6Fw+auaiUdNIYtUEskuA+gs1
PVgn66CfwC1Di+gbyPeOi6fB6Ivwe0g8y7kQdq/9xgJHmJZhSwNHr1+j7u6M
Jq7P4Mx6ivUkXudh6Uhznul2RYVy6A4UITYkboV//8rb/viMr6onlGAg7Ppl
/H9cM2yIreo3j287HXEwLof8hWlgDj4s334metiXObmWJEsFdoV/4jkqafQV
g0d01Nv8KjVBIY/z+OBeoPSlvqJ+DT/54QD0lVQ2h4+B/Gep2aV6jrRPYixz
8ja2Xcq5NTVD+7owkjw11eKOSnx3Z+Zd7t8D+alYeOz7b8rFWDFGVK4vRip+
9cvJjDtpbYK49oGe23rfRLTsrhHjQ66StS9iJpBxNVbLKrh7iFxwy1oHvVDz
FVyAlkIs3GBotuIgeIrWxCsfd8ny3k69PvwwhuRMafpWGDdfqIzaSlBr1/tz
X4Fb7+ZLJOS27ob4N4orn8U62U2fnr83qNU9Qh9sLAHl2AHbKqE4Zqx7wDGW
6CMhjoJY3jTxzaNbvq6gPnBGro1gCAX+BTJd95CLSXBMNSz3aX5Gw0CTqZ9C
Rj/g7z0NoCv13U+jrHLyyTy6NiFhaVKzLHWqvQHGB2W+MoFm9UCIQu7tDq5g
j4pz189y5o2cfrK/3TQafF3HjFAX7Ls1gidLC6XmMAC1HIhRlIs7EJDZsJQr
fxBzzxzSETAIGE652Hx8l0BA/p2R+WSzFQ8do8f0ZyjKiQtewxn8L+/wkBch
b4gMILevmznIu+mUTdawMdQQlYKSuBGtyPIx4D0ypS3r6dNKHNDpaFruOKqT
BEg9ob0GxNyjJbcIKLhTyOOt05a2wniTRtBUxZzC25hqyOUp3kfrBSvLJNH+
+KoEriURqUtK9lJo6Kk9dnuFqyN/JxIJc8YO8/wOx5mbjnN6nIjp6SZCL7dK
u4s9akN5b/Gu+Ld5oUNCPkFRDmhCu6F+ma96zxrqRFr9kuWOWo/MUdN5SIkB
5mgQBSXRQr8svKF1fBug0EFDmSlIT0tsjXP1EZD3DQOmMSbC78RSemhONSZm
1SXFM8c8inN3YiNiO4dcxZ88N/wO+y+s+EBmS06TlIsFJ2ooJi1HKXD48vQu
oUSu2ncsDNnPp5S5GGS2LFx/307U0kZP8bXt/RFxO5Erdmpis4TStClIBMG6
nuUc10BJyFC1NWsIMgS3lchBqgiOe/OK3mkuvZF6U3V8vWtg2e1qJ6S+q1mJ
N/h8Y7XME8aowSz/IPdEiFVrmlNIyp1ZCy+5TAJF1c7DJwoVWIG1Z7oQwSXs
P+qAOAXgRXZBSpGFKQEULmZ/J8vEgOby9qqgpxb6wPRie6f1AZM2Nl5TQX8W
7Y/yQ1XNlCuVLAEhb5t1sPkgg04/OFU3uEuDpqZWOX+i/5nPlFfAJWgkw7+l
ljxks3hpvVf6fV3LntnJbUvM3HNBDL4jhDwS/gm9gITYIat5wtbCzPR0p8uD
uwiQnLOQ0g+yEzO4sLderlCb2LohPQsJcWpLungMbaC1bpLH44QSBSuoS6uV
uvbXXB/jnaFx5pfXitnHRd0hvibrA3WjQNmoF/itTvMmY8Ryv8Wz6J6SGETF
TbqKmWLelbgzn6XM+qSJZje1hrLIEv+oiYoGWfHxkcE+ZQZ37TpEHs/DG7lS
hywIeT/5E68tGM1jxKlloLp1wT9f7RiophO35n/UfgR9NhM0YtVzR4oAGGAA
Z8iM5enytZoV7/zXmncd09O92CYJeWUF0N2VBmfFdPT4KcgpiX8DPROOm6wf
ZT0msh1dWq0Agu6UwmbW7ShpFv5TPerqrORpotT1rvjCiEOhN7d7VD06Lh2I
sJNgJ3u3mirVESSpypFsNvakayjd6nGQq78thkWgm6en/UF8Y0/A5GnInfOU
lz2b2rLRK7lPNPqyVS2l60yTdqpH2vXlBEfPxM6rzbLjoFwaSiYKKit0cr5M
8yT6uLeoNTYYdqT/e6Jl5sr+HQQVe79ueZAzs+dOuFjKB2RU/8kblk/y5qt6
GLyWjY8lXWZKaeYsLEiQR3ZoHB4Erb/8NkWPD+TiWFJtK2RdG2Qj1uo30WC8
Wr35WOc91yvGBLVErkMkgA3TzaX/J2hUBObphuJOiIsZDFph/rruKCJHOz4n
8z1XUer34r08flufWL5ma9M0R5du5varQbZ9eLMsbiU3FRn/p8aPTAjpbAxY
ceu/shahR4rsBMnJB5I56sSmEKvo2MR5YrTS2E4Wh648ydm8346s5yY//Zki
EBSKk1LXjc4uqDihKfwVKo/tcqBfyV5FPWmnhRe8XlJp0ej1SiUxbqoDCqEU
w/OIU7etS78mBjzLSyM9g4T86FOWcRy2Q54CUTOK7ht6Klxpkfb4SkrQNp7l
1c4m2rfdQpIoXDPemQNvuQePaxgcg6Q/IsyfWTk0MYgp74G5F452LDk+x6j8
HRa9Ws8GTqcX+gdTB4CEu6GVg15oOAR8IvoEfj/Lh/BLCZoO//JYbRLe/ucd
bwB26dE2qB9VkTzo3Wt3So5ByhkFMY6DJSVvcNGox1JQVECxef5UMgV5DcRJ
64oPQLly5yVMl9LD+jKsmG4D2rty+S9uqHyBlFqT4BLCzxi7pXAkK4F1qIpf
sqPSFy0bJuma+p8N5BLhPpqbQp2GWPttKntRyBiwXK/3SLr/lKk36eEEoazX
Tb62l91EEQxtbUDOzHMgoU69Pvg9R5jmoZQIbh+H7r2TsmQHAmEnniLbZ4AB
2rmPANjGsTc7iZOG2VK+58NwIgE/ntwZPU4PbONPq7CgDDDBlCvSWVPKmqm8
JGgSl04LWsMFzY/khZsaCG/J0vofuDz/bci/uzP4WJDBeqigW6XHhbDVVh4F
RFn1XhjVjI/bT3dpqcVcaQURlcpqTHz/r5rOLSaJTEkrkXiKKsTqlZJ9JviS
epWLXEbkunVT8RIKKgw6tfF0ZXojbqyYTR+Cg2yMuPlAbHAFvwId29BbKzVK
b4yQ0+txtfq6JLyMU8fMiKx7U6upBcGmDDcjlfV7LIqlS3gXmPdPVHRZ5a6m
84/oxU4taab13CJA3musd9oMBQ40KYiIF3cKzRxaCBA0dVHlUDuo9GzLxqLi
xH5CU3E/RhfHNzxgN9EPwuDjyEBUClYMckMy/H4UtldB3uC82yMFIkQjTKin
/JK1szRUKf+rBkEtgoJJr7E416uFD9eGR4fxXloR9pm80Tcc4DVFOf2swTQl
cudJMN4ZwsxQ+xSj/4FYo1+jxpSOzzLahgtEM0Wzbme1rDv9FCP5rtPLj78k
K7Qs406O9NpV9YYvSMkGjOm/V5JAdJa3lzIegJ+XX9Bu7Mn8pYYEU2hYDUL8
3y4IBCBCqxLRoJYNiBD0WJTTPyYkjxVOVKXLpd0cOk45npmtvlvT0dXONXjY
Vm5Qqp7196XfZeYMp2/jHXXISteoWnAW++AMGO95MaJakbf4O0LwMtkcDGgi
ogP7OirvCKBw145w5kBgGn6RO1o3GAIGqTeXsVLl8DAV+XV98SopVZjuNfse
B8rLjEcM4xWC4NaH27z2ixJZ6omg4gQuqTE0KHlbSoZ+fs5FLl4XodPbC9PK
tS6DV5DWozqVle/mtkP/al9xyMo9k8+nxQW/KzsZHJfWbIC37P5Ls2aw2zzM
WTuuQxnvBwcrxoI7LJ5Hs8j5wRiwGRwA76WbHhbcAlz8gxHAeE7zzMKE7dqz
K26DuqqKVXniJZvtp9gC2N/IYNfNzANr1l0ijIaVs6auIletqx8gpgcHYEH0
5RDO+E6McXJ7VlbUbtoSw3NHPsntRDCo6JoF07/6hWEd2o1zT5uZwx2WilIV
UJaIhhoLvkCDVuQHw9wAFDQoeBQB6Vys3Ld/onYV7W/9o32vLgFTctFrRuCu
SMf+IJcX5RxDki4O7apXQgaGuXABq/SHnVDYpourRgOm+N+ZU7wu2sPOQmPl
V+A7iHKpSIqNLSldGGcbe/vhWvp/nKKsZsr+gC0ewMTKOC+C70v+19mC7rU0
t+uL1CtStHiimujV/9USzOxV+jZ7LVePBOqREJ4I+BuzPTxMZsY1fN5Nuf7o
lAOHtIm04NiGd2M/nwgdebykV8nWtWTHcs99+HW+aIEqOJBhAFgfbowebPHT
UmyVG8zvXRy4DgarzkIOuv/FppJvFzKlZ9fbAXm4z7PZXYlVW/nTjWp8i4A+
uy6PsRIiqFjZi+zJwRVNgasnCJu+hUQ3eWKDIkKnH3zGfntEI7rF4IWChRnE
PEwfeD+kSCPmhP8hWXGs6sdt5tC70G1Vs7ZLQ+vpxIHkyytA0R8ZVxPkRYfM
RrcTHH3IpjRdxZp4tGQRmuAHvdI+gHQrfncvV2xcHeG+F7VTMjp6VqGxPMUF
vfkpUyRv3GxiHTCnMJsfyVTc3gXkVxNwVZIUd5kI0x8Wru0/lLdUaLuiI2LJ
niZyDyLfkAyqZMAJ/AZzKeaJfwiHfGYwHba1JCdNJLuVEHliIySPswWch0IN
B2XbHfC7ILFEbH0uMDiWl2gB21R3ccDmtOkBEbKF4SjQvvDV90JctTeyuRxi
oAOQH3aAaVuZiBOXltNuwZ+dhv/Vx4HuuMqV9Gd2Ov55YONtr0A1akM8rqpR
q3Gmilk/ksi24N7qlmvZaMHPOR8Zkem6TMz2MRJsJXMIfBM973F99BJCuHxT
KoVEx2VxdK/GjIWC/beWc8/11tUNGh34h+eMB97iZHkPAWY43zw50nf/tQD4
P/zdd+y3/C/QYshpzMBSlLOwfkYLSFnUTdvWEtgIGxiAliX8F327BSNJYjb+
bijSD99BvCLGNZ+E0qonILbkD+HM9lwrM3xWgJiz+I9getx/6mGzHBV3ZLv6
gJWOzWDFnlPxk2camdG8po8AgQb6648WjE1GYGGGlDnRXxnYajR62inm3JrQ
kQ//3iT6Bx223rrVeXfLMiHkstZ2DJ5trQNRLxXVBzCGMkABa9YpOJ0Xn3iJ
sXxPjKBcUQaa+Dqey7IVP0CvGeNKF+bJrinOAcJJVkAHGRJuswy9GBX2VMD/
h9T+xbOwMJHFZYa5AVY+/nGYLzTmEpcAxuXSrG/wP3j73vt12ZkhUDF4fQIx
tfSUinGOHtdZMUd5eIewdNJzxNtNYRl4vUO0DpCoRJ24tkTdQEsO0HkI4xNm
PMeQZDyG5G+ZyRKCs8qW8UrD1hp01rQ2WUpd25UEn+yOO9WhPTCw4hpCJ688
EH9ZqfD1mbgpKMpgRvYem2z7PrtJcEbpKzN5xbaj5VrETWfRfMEreWnrPghk
Cf39tGfVldsbBxbYT6AXIblVJ1ZY1A96b8kySUQnXa41Mtp8pjtTllI71VHQ
E6fQftgeV8HwVpxCdvnOCVUHBgXTMfr9HcwuoqpOuXnKxQAVSy5JCB5vq59V
9dpKa7RVpqJT4h5gvpuXgi2q9ZCHzayqCqsoYUPTP6zhRgv+UubxafpCwfkJ
TinVUsdt5uW2a+/ObEzNVR1xkrTId93vIsf4RO/nq1B0DMhbpn6E9RCGqTtD
5LBprmAlQgZtjg/V2XHd36Aia7aJi8CEvPH5Ts7HyYCOA5vYpDEHweSU22UY
a0RjvgD7NtHcWyKXsEq3DwGfb9KK/c+HT9JsBIDVZfNaQUpGxYi5ADfCRaEr
+yFnVNt99W1gRdFw68aIosXmpmdaLPfMuLJLIaVynqyroHxx1iWTYojBSANe
wUSH7uo8tt1ThaLqbtBmUxWe7RgI63iCI0EFNKg3qFB3dXMd928bSZ6ZIJhh
nV1RRVniXsnvHruHgD5NeVCWLT8aqIdSvPMWohVOchOnStTqHBDP8A8C3HyI
yZ4NltrGQPkay+YuX3DLaPmUJKkf4k5qny0oh5bIYyPiSq/SUBrJJYT0rkKM
GhCnghyN3J1KTyJ41SKVpr2iXFwEhc5ojweFaakLvIF0fzB4ix/PsFnNAhbu
wMr4JwN4MtOSFpVHRxTFqSg/oRDXCG2SRAm1BKNh4iVgh59Y7w8lFZz2HGof
QbxYvxMpBFnCCypspV+akbLo24eVtC8zzIb8XP6GPXqD/0d05zjXX/w72oOM
ucz4CbtB7IUlskZi9Dlt0c8psv/jkiWTFzwe9ubhVb46kY21UeA6XU4WUc30
/TZfl/5SABrKk7PQx1dNhhWAffat6EnHxdihYQHS3DW0SvqEWSILj79zDc03
IXurPJeLAngAff5OL+RTPUmGjvxkbLOl++qN1+6wGfS8tcvXbB15B5McKgeG
SLIeuz2FMCBNQD+0FZrFebU1ObpGVeln6IdfpRKYi92vsWgtG/1xX3NAx/a/
VvKYTa9Z1EwTf11et/fD2jzwJlkypQeZ9n+4QvXF6ZLihSdcbTV7tn7d120g
ONGaKzoXr2UDUN38oQ26z9+v4P08OIEAQyHzJ4Qv+MlHqGAMtKm4bgShoY08
7JSZ2Z3JAM31e9ZXsIyxMKSCLRogSPxuUtyHzHiIYOP9Jd/yG1pgsDUkFKIn
uO58y22/YNYd98FdF5noYNEqiXK0IPycaFZMK+EdDT0/budPg3Posjcbj/5f
/jZ759IMwIvdeJHp21S3XgmjCyoxTaj1l0RapdeCgE/SnUzZcTh3r+KuBSV5
B5gXno13YUMBLhgiDwG5aAYFh/xB0qx7SzP/XizgiaHGlTTjSf3D1QHHCsD2
HnZyJb51bTXYdaJRu1JfQvaT1VA7WDygm6IgYPnNwnsx+QU2d0rdIA88RzJt
7cGCJCVQJI1/MpzZVeRnRK7jQ6yJwtopnmtplfA2FzuNl87ioLKQ06peWoWp
uxWM3oaFXpKvuVrzx/Vsuuf/v1YPYIVTfVRFChd6QuPsUMfZ+EKrW93KXKVR
yaBbePEznKGaT3AC+28t7lzyGYebrHA3jry//AJ+hpNeFipkjkMLhDF5/mri
PORzCkineIrCYI9hVGHO63Fr5kdF3gixbiZ2VcyPi+nKWfuaK639N57kXrSQ
xVqbqRXTNMBJ0ZKhocTaW5tR3xFRt8QrkNnGPtQwRVsmPLPobbbaicDY87t/
tvK1kMffJdZCaRkklhw7KGh+epJRGhj2Q7OBW16K4pU+TZuG3OtBM9GGaizV
jkj6awSOxpX3PcU1Gnroda/YnTlhFSzN+EeoG7gjII8bPORR0LnKIhhIDowg
ZQkBeb2cFgdFdtGiJdeibR9xOnhxj7S0DEAXoIqCXGbTREkE+SlJN9/fTQJp
EkHBzQmt4++ShWEeq63pQ6qrIXMQDkmUSq8DDR9WRP7n7ucUEQQImfWpCQod
e1aYfMDpLfIBqeW5wbGF8eCYn0/7iBfpQiNWEAX9pNifEpIHTgMi4kCvY5Wm
Guh4WL9xGbXe159c7IpKbCey1HVBTdpyefSk3lwBq+J2c7XiWNd40SgnrQd9
WhdyEzHAqjKyL9Dsq9UVnt/eNOs3r78xqUW9ycneawEY4UX8ozMXiceAiI/j
AWMPhmAzNE2WRQx7ptL8dtsgg/rg0LxuTsV5GlVK/t3jNFnGxbDxYdwTnCZF
zMAno9ZzEwvjTFnMWM1LtrzjWymER/r/asdVRycCqmr2BG5AIzeGJXvM2rJl
HDrrx/Mr/JzxuLGKidcegKFKdD6ceZxalPH6HPxKoDr+PLyKKN/qFU87xrhV
smv5nqNun+BHkajx5Dy8mXSt26GpQDUHu8BFNsAHvIPtA48491KFXzxfvzOV
/4SZawNikz9VTEeo2HzqWWnxbE7QN/T26Bb3rei3kFW3wKQeihv0PCrVCEye
Q5Cr36i1TdUa57/vTS33KF+F44Vm+58UilBLxBFy0LtUb8f3UT07Q/IyRkDi
saNJO15IyrLbuu8ny05mwjhfAeVUZZn6DRhm1rwhO2MRxEYVRy+/tcqtQWbe
V9XlH63S/LV2pvLoOfw1bdhH9AW0sl+G8bidoKwvV8+3rxOe0u86wAjz0Rhu
C+nkSCR1U/1lCJ7n9P4/M1H9AdVdGm5UKMpxrn65f01dkTZq+F0AjGedxxF4
2TSUG08BOEeS2rhGNLlPEkH4TAlDawDwWdJ7UlWbDH5YNH6DEjUwStVgalT1
ZMakEmY/EJ9hGJ0x925PyK2fLq566Ai1QY+qNBgowKP3NNm/bQKB0bYvbiT4
gHTC9/YqFaB2nk8sd8FMB5oWg4fYCsQCx6jKySSNUo/YxqYmQuxJSMwfdown
nI1yFU57kx0g5CzeTrGNs5rRHiUCLQGkBg4ADMO36/Lz2lPDP675A3nqlanP
3LUG44Q8Ua+IVLIWARx2NApOmLu+lyc92q985f4REioxUXi6lHt2WT+sMLii
3PDwUBRcm7uoJVAXPwGeCQMJRci4Q2pKLsQxIU6yU60Lvj/xcnsIxjnEbviu
9cx3EPc5UhkgBVEX5Ww2h3Pe4E3ud8RKVp7sV5qT9i89qOVHPY5ntMQEP7eP
aR9raMRwQLyAEFM2GNDAzxAskwwg1ZKp+VSQiWNZv1ts5bjYIDCKgm8BZ21o
b2SQ/O0LbDSBtftaDGAxyEJHv/fgc/A4ZS3glMzkcEScXLYTtzFz5tPJmlds
XZlBu7i9XW0uHUVMq3EG8vq5OnGbFBdm0VcDSzfRMADVGSRmgFPWnJ4dwzPe
k0wfwT2pMC1CDJjiRVpYNUkkVwnyeRTRUoRm5WBPwPuO/i9xbgGE0Tas7Dhv
hX7B34dFiIhXVaIROXCPYmTiJl+nxhg0FFMFyutnUd807MKM0qxu0E/p+aRB
qFIGDRQtf9VHONmSdV8XCQP/9PmNAAAILbrTz86WXWEljuLrghzAwMNkf+pP
Dotu5F1mMsloxdhib5zj71y1/EGOi8zZs5TMhTLse9dVRiUK+RiDligS9Hp8
AI5ej6HaMmoveXvoS5PFokFNV+5hTNug415W4Aa27B5iPbwr1Q9k6ua/3n0o
78fuDpfrhi1dEOnGotQeAR3Gsd+4PUufJ1CAGewrgVP2vqA+2B811Z6c7QBu
65/DiH+/lRBuftubxSv9R46DV7v6Uho/jrPmE2RgsBKgOLxyt+AY7w6sociK
SCUpPjvuzONsjZy0O3h3joUoPRLimckm6Agj7gkE5HyxZjATW3Sbdq/UGl7d
eHa5o0gGZ6Ou0yCbHSEr/VR89vdMml+ghmTOnt2L9yJdrLfsxB/il28T5CaH
Aiy0jGi3D0QM1z9Q2ycaS0BJzrEEdA1srAYujA2JT2UCjGB1QbeTZIcVx2BQ
8+G7Fw78y+BbS1xtAsj6ndgleFyvbKZeC+BLDAJ/l1FdCQicQjrPr0sXeFP5
61rk9feLg5OXGKpaXT8h5WorsDhzjo9QU4Y51FMgvam9XJAsQtFZ2mnidSl5
HCtx6kHTsj3jEawXU3gFroC8+JK8dw6DaMXwclWZ4AsFZf6kXUPMUFDoJWUF
cjs3/MZrTbDtFjKO24vV+11hPhDd8WA/zRbCRktclDNRSVykrxUyYo7+zm1Z
ptyqGa1keyqGpTt+mLwMUXc4exbEHyCIIzgAC5sOJ8PsfkRbexPmdyDK+5hU
P0Ei1517J0D4DabO6tKqdPvaj58CX7F1ahb3+j23sH/pjI1LjSWrpqRMn2Bq
mny6+URcWOinY5l0rj5rxmHYXVvXRkUIE/1SSsr7C6Ddsu8HWN+ceg4IjhYy
/XaU1Ub2F/f+ErOQVdBxUtdLy6LFP4rcO9D4Us8MuJpHNot+vMKjmcSJIJdv
RUG+0KzVgzCMXC72faku309kyJtlVXgrugySLRC1XjQ2A7UTNGdutq+NCAIF
JSGG6DMnDhl15FmM3hQIoQJa03cEb7n6hcuZ0wpvZYATh2qIy2Ox56j7r7wk
usPQZo1mjvbOAgLkI+817ESR4KAFoH8ze5YIPMF/SLzCwxqU77gH/6Gbu4vw
JytMLDqgQZR8h90zdr0N585R824TE+GSJeXshAXO3FeSHT+yUl557zFztaq+
UUeztiAnCPlzyQ57rhCIx0EfSLOabONTpLg7p09386s0hZuPH32/M3uOf72V
E1bioEJVzvBdU2A6jGVvasNLDFMVKNbUt3W7uibS4nB4Z6hwypvQKe0AwnD8
VIWZ5hOO0QEGL69LZMt7fBxQEJxc3epgS6qatg+qGMyRz0yzwYTPle+ysMAT
kA6j91o3BWxXt4f0PEmmAlXg9rQjcLRjKLUbigVroXYSaDgP+dBthXXf6KWx
NPdcJ0aDqF+toPN6IeX6ldZ1EUItI93N1HdxXOW1K9f+NSkQ/pW4VX5qPkWU
MWFrefEkQfCjpPuc7QGV0G+UKZlL9p6LPOyQbVdoCiJlkLXEeoFcWXdLSTrc
6zw1UrBBcLmwiNJweT0aNKKoKa5Nx8U7hx6plv2uAhNfPq82QjffdSzAC2Bn
MckbdPHOEXxpEfVJYlW5euN9QGne+OQ6rpjk7duWauiEoGiBQLYHR5Kdfxsg
vnECRIrpf7K/q+kg0nLDIMVbkvCqsSuv1jLdlmR9/u8fRBaSVHtz8lBNjE7m
M4wJfX/8gtAX4MoTIBQFjc8b6QCpfhLjUVKi/bVciYVaFghGXfNRlGHWGY95
4T9JMgtNEPczy+YiXmp9oStHam689Q/OheMU+HhnaD63j3oARTAazi7IyltD
Itcly/nmZbgrqP9a7uGilXYRWmeyKubt71fFYrA7gXUc9Ac9aC8IzBAw+GlJ
lESu9kq88KWtNtRYb9oe7Wet+j8RTe2133INwqlmfI5xRLWvisR/4ve/e7F5
ghxOaCPX8VtgaPq1lzmQddymlxKBkF2SG0fhs31WaxIijYdH0h+W98j+p5AX
Wp48wQuwjLwjdNugP1UwgnSteQGgZ9Jed2N4Coqd7nW6InEd/0khNb4u7p+8
yuO/0Kg5AXKZGB1z6hbtyfGr3szugcdPHcT5NRmtLDHlX1Iptwv8Y09UJEhb
/EpSXKH5LyjjKPCzkti+vy8a9XbS50XLzKXbkCY8C4K3tENApffH1+hv2XjY
k9pcB4M/cNFEWOr0PEtmrtW9vMZv6zCfgFmcXxCHGXo2Dy8I1Iqt8YPsU6WI
jVXoVQRdzrMNnMtN5TokyvO0liUBUIbZqj1FS3yyjo64AZAxUb+hc/VdfxMf
Rdo5SRZwlJykVB82AGUUFDCrd1MIqgbj1R9w1UIxR8Wtj0TQvs8EproQX7no
+rHAVwG7/yBa9U+CfcywA2Dli9HEVyT68r5kYQ/IwKRDurj6PgWpGCqARQGu
TGs/sXj/7MDlzvtZ04Gh9hqOBl9ic9qDuUGK8KtnFTAu63dcXRVzOjPZlpTI
1a4Q5dOyfZDTRdk/4H4zoUnE6HXUTapofhTu9hCIa9PV3k8b+srCigkKwuwR
qLwXjO199z1DuMsqDqkbTaXCJg9btx6ifYKMoO1K9K7cfNmqwHMjwGlYcmY9
vKijyfnohDd5mE6EUyCD2916Ddfx0MMK1xKdEbGUxCCGdlNXWN9G7A4E3Pho
xaAeZfOmOqJ8RW7hnthJCL1qpV4I8tnns3yqwXBLjDZldulCuuthdYYBfWco
VGEgAsHwJXKmcludzR5f4EFxrt/JEmPTLBzeB6x3CVOBDOy9P62fEVs5H3KC
PqRJ9WKFyIQwGrYQ0jVn0dG521ku79iiymcsrqdfQuQ63FL+4B9IgauMT5Fp
OVkS/9CwuRgEOCtmHSe+8eGU3Acbmqs8A/krM2sbMQoCoFK4ihd+uku4jlsJ
rGxtXyQwzLYh8JKS46u9cPVS/axjdNgz+lE/m0QbLwwdOSD4xM/D5ctHNjTb
kchEyyaOxwTcHtEI3RKNB4MYmkQFVbhP6de9bK2R0vWzOy2G5cEgGeQpjLSM
qO7ZIzTQJC9j7B4IVlg8KYYxb8oD9x6IJOzmOHWQVksTUyHOV3hSdjUOcpN7
byMrYMeagAxs7OLhEFgSMEnJLs+1QGEKyXjQi3hm9L1iAa27a9UbmLvX2Rb/
+dM42u0EjOeCFG9ijRkUEUtjWPhOpdehp0vTalhwJ2OcNPF3Af8uzh9yyxKN
amQXQq729jHVOWT2lXWkvYHQ56zPDCh+mDNaueIAVPO3mQCiGQ4rkBOhMV6Y
nZLYyFbwHaVXh2P6rkHpIgDwXjHAJFd9m5f1jkmmVh+f4L6t9AZxTfkaen2R
7zyNwuRw8Nxi862A2LdHAGqCjmICZgAs/uECIsXqEUo7X4Fu67Mnurn1MwdT
lTZmYAJbYBs6IEPI8A1EEfvLXi0d1Oj7ayZFRvopWTm/XEQSUqNGIGDBLWMu
k5oyVsV7SoieLJ3skPpqJXjxcWD17EZm0WHqUYUUowNjaGpD81T6tf6niCCf
Q1/WnH+uFQOSFYjr9GEC8SbPrTWhOrlaBl/naEJ3dTqY7CFHoxzMTXwMjMTh
ClVLTITG29z0XdE3lOW1iW3CL4bHbO9BlEq5TDnNujEF69LsxVW9ytEuDyAg
7wIm2ZGk2CTMXhvT4mlgNKJ6v7e7aTYt6wx7RZAu+gnYL1sIXPKGhK0tfkyq
c0pC9w1NyplEiBCptXvRNNYqP256eStz4jM2xgJsTVf1QnAKoX0Nr8AvcC0M
PxplnbIQYwZON8cdxbZVg/qw3+/H0tFEVseChMpZU+2Go5Bbkketo/3IR04i
zgdzYTDUGr8374ZV420sgQquilDcslbC0uxtVaXj+UxF2bKUFKs5l4S+G/4N
EzbdXZlIA/hsqtDh6U9xaaTAw2Kx0rS4h1+NGh8v+pUV/zt1LnShiVwmM6Hu
WUKIWyjDDIEkhHHrc2JyY0j3tNUlHuC+Btr1fE0ci4gy/ah4b7driTonM8Zs
Q0d2NUDRyva1yEloKgws1YO2qeFnqyWj51D7h/Lh7jn6jpoGKaL3c6PYl7/U
XleS7YlbnmvZeMY+z39+vhx7PRblqfIQer7bjOGoH2tb6JQllt3nb09+bg2t
XiypB7znu0I6D2ntMTcVIp1onTGn+KqOlKQLB0eWHvcaT3dtgRrDcatRD0nY
1Vj7jrBe2B+g2iUSEE2fM0HNF4RTONR1n9bEEXnVn1V1lWytC9+AHmmZED+V
UrONwhUkeehecwkNECflc8NFWdCARCbU73lkCSmVvPsqPEloLP6fZTIdayYg
xlLWKrQzoPY9eavCuDLVNqTTdV0iy7jMLi4dxPUUiAe0haV6V0pCQpW8peXY
oEnvLeKaa9l9by64emnoeXubvE3YMuvgFHx+3gvQAU0SsvTuOj/BZ1sW1UHQ
fG+TPmhc0jO6E9XciI/1VT81XFhHiyjbcSEzBYKHAe83MJrO917iKTU7OkHs
eOGar2nhacGXqfiJlmz3WfB9Am+enpyr7PDd2wyM5C4tE0sWn0ayr2qeZx6F
rY+HwOnTMIeFrEUlXxWQFDviaCDo4A5Hbl0hcNjr7zWH4o5lps6gjrDY2OXr
u6wDj+CDoFQAQH/5X2c0+Pv2uf0E8MHvr+gG+nAZR8V1HZKoFgNvlpyb1bXu
nEQu9A5lTHi33p6Yxh+a0sFnc/QhNTXjVd/HMULTR28n4DwObspUE/sajjGx
7+v8THYvawNQ/TAw83qgCOGTJL+N8kvuKpaN+WOv5RQMEGIlMnqbZB7x98o/
0RXAdygTVHbkfgatLJa2Y55isJ+8MxUkA7M5ueJN63VgGi7GK8l765f1PxFw
gCswMDHO7tVMhIH8WFoTzcUBpTn8BnoPGSzIAX7iQKpii4MtHTRqVAuqluQv
tObTwnARXklLDJkKejUzjMTxzrIYH0fbZjooP686crJWFPrYgRR6ae24umAM
pxYkVFSeDKMRSFmKV5nPqnxgybwlgWATvbmjZDkcbNPfB55gnKU0vTVC+VLG
2gqW7IZlBkSjUsdSmH+EZxj/81D7idlrTlRyJdLkzCnxk4m3b46zwun3oDd/
jx9Tsp04aOssh2gJb0pwAGAeSbkbATgI0dfVErYzY0tn0ykm2QlsnfB+PUBC
1iQUwj1IviZREZQ4vwu2eHyvDMGv8WRFmyGvQBI0FP0cN+aLmsOcS5co/nqv
7Z+Qz42TZhn6s9lmpb2r3hk/QMHpHazMCHoXN2afVGPGRarGTUi6NPnyckHx
BoUqK/NoOND8UT4Ji5EBKmp1CVZcfuY0H7pIGz0YvEiHIspuyHWr4zrlEuVT
Kd/545HOGoJqUxGcor5iuI64pPX+jHj4JPSkfRbnvWY75XPPIJ9k4AQXCAs0
NQx6Fg3NdctA/Z9GQWRYQ282FNe8A+GjtgKN/0e+moUmMa3xTkt6Jur2DTsX
Btjo7F7XxbxR1C6b5BzdAILzb9POa39HpCzv5AsKdjtSfdAlAJ5DqjoioAon
O3P8ZSUtZmrZ+HTBlJqU+5dD95NXAMOfE3OTt9+UD+/D1WRQ5tBYpIpGeg8M
oXgtAa7xK3yOOTPywCYT0O8cc/BTLPo/ZBu5oIzVSqW2wwHfD9Eq7QT3cv/K
dipJAOaIb3rJAwMN5VNkFCfQ6DhqIhB1HJSAn5gZHKKERvhDmnowvgVrotsV
3sqVmphZ514xuzwcgp1zgN7e+AC2FJtgZICsvPjT1KuDEewEAnKSBzo7AKL9
cIN+dwpQDmmq8mf/tv+hnQ6L1SWYESTSEuGuBWV+M7pSsBCCa7+n7qU8PIOV
sNY4CZAe9GFpIMtty+Mj7zPyCQ72ZgfSQCHeEvAQSabSNWxac0xogKgHFRcY
9S+gnKybxeeKNWOOwebg0gNTErF9B+Af44dHlgOcGp7FfTvuhcndcrBVzIyT
qrpe5ILi6T3+MrattlMcXUlktckmczaAB9rKYOswAO8qB978zzuaFyfUSOz1
bYtPtI5TriGuwATI6EOsCGRTHg/zL/GRIZ5ALI45+ZFr3LHKekXSGYpPsk1O
gPRld+xxD8zLr2i8WaxsInsBsxy/FwTsphVzQcibpAa0VYPwJhHuQ9c489A3
io30V0frmVAq5gJl3W8OvTWyA7vaU63Ji38piulhA9L/XPFcHcm4l6Rv1oJF
vdjA5StD32HhX08r0ifxdBRlhoer1X78Jm+ebwFKplBG/5gFGfkZbUdrmwk+
jO+5xFbef0Lqcmqraayj1i55tbcOXlYcHI4xR81xD3vN248WGu6lipBOhJKy
6FwdhycqN/rj3gA34hFTqoAcCPlFKJTgeNJ13FU973EQdpFkZ4XabJPH6fZj
cp2QyEOmZq1rD5z/tMYw9/8EfY9KRdXb5f7seuvgSZ1hmtwhrQdaLGSNV6of
iqNapTRDfZJt1SAmbsBzboRQI/l009YYcNINPZgWEzYGDc4oEM/Rk2TgvJKJ
0h3Vsfq8ImhHrvEOlvlkF+CCGFee6Hyaj6NbMIa7zlvs/sFQG1ZZg8wpY0VG
5pTjtA9ugRzbhVd4AqzGeyCJRHqVy8Tn7taQ9esIaXUSvmUOW48be9/rRS73
hZ+xgk54lgWjYIB/sgj10nMtM8afKfpTqxuO/OGjfouedbcHbsPxRH3/ri/o
9pIA43DFuTcZvbze00JSmgAhlLQymUi1JIdJGDQe34LwxwGF3CxXoRAIR2Z1
dd7ypHoFB49ozfzKbAGBbW66x0kJSBT3IL0tCGnLEIho8+pqtj9cbybXHLmA
i5q3STx3Ha2gxbGI71RtbtFCilRpewLWRH8dVgGpmX/nvaZvUGvsvtLLGMRc
9O1+TzAWK8ZK3DEDwdeQkm9T+LwjhcfizF9iD63qQfCjjcmJjKQhrZ2Vn+3K
KrtHiLnqv9AIUqZ6gnh6b0t6avKqML53OB5iRthatFMw3X8mSHjNCm9dJFWl
WILayU7u+QN1M+ec9hbt7MgLvbFCphnRy4/0mHSpBfNJuSquWhbjiMSRH1tY
Ab/UiDXZDAJJYM9PBfdqshz5FM6wxkwNg285vJ8nyKa74N0qwWeWj+kpkVJV
lvANQNXRfDLRr5JPIO1zWFqYgIaxlh/ram4gHanCwmrCQPp9G95gEuDBJEqp
8WQMeFD+f48uoEa1YqZ+kbAvKSXfZ7Ji1RPs1iwCmuW2KnVj/OQNsEdJMI+v
EmZdZiXHYMw4arbAffB1T4IH4PPaLd6mHHq3hxnN7fwKEbj1rj9ERp5BFZ8+
7laZ3dhfB8EC/gpIxicfhCyare2fKNGy3NkGmKtPq60I5gqKzYUruNjoah1a
npS72gQK93dyJq8L0DaP/Eo6SEX/mELg7jciUcYeuB/ROo44gZn2xoyYGNdY
rUeFQWCnin2YhZ/6frxDH/M2hmBCf3BGflGHAqK+ls28thcu1+TK0vPDZK3D
cmV+ntmaRNfM2WIA/4KeCkEKT0T7BVYChNsr+rPbHQ7MOhA7P9/+YZNvxTIG
juQDKYjyFWaiOY/WEPlCS07vuj+BLzJWLc1VUgQSNKn1r8WNFVtUQ9lOT/Kv
3FhzDuPj4Wc1kXyxkLh3i8GTu8zmeNNYgZdDXBg0FCg8e4CBE5/m/wSjThfn
t/hp3OEMrDo0OCDJlBvgixV9Jna6YLon2gNcCWNpYeIXfrZjP6JiwBgKiDxy
b9ckxFvqxeYauGGwRfUGHf5XzYPtO2/XU8/2SN3QJ7u3LtbxZ9rSK3nWNM5N
HH+94Vtdf8YlDKYhmObJEjEUZDYVt99DLyM/Q6aOwiPksz0QLpL9m48wl+L+
i+6he7CE63h/GMDO5z0g5rk1uLxh8JVna5nUENkzOwqpe4ymUSvx19s7lsU7
nSlbeGKBgIhANyeCxAwXWXSoPK9z985dx4hxvRIUjcwh+afsRYPPv+UyjLZA
/gRugGYK8cGUYV8A3haAVvpA29W5Z2JeJPWupkVw6x2AMWKXJIw1R5Jz1oCR
A+4jTwqGgDtqqvweukVB0L4jckRhlyK1vT5hBLZcyygdjhZ0pTuizmFg7Osc
gb8A0i9jRK/AYaPcLS6+9IIi1PP7hEseTyKGvKwTXZuer3pNDgyK6LrygIPj
y+MRoHnO9nj2toovgAMlwvQ9rbvZcPih+Oe9JT/DRXrhiXtCXFlleeoosGlt
tUxp0BIV/IjZPz0MSrAbwg3dIDo/m3PWNXgxq13rZXQEeDMOFN6iVY0jnU/f
Tj1DTCkGXwrX5qbmFChwpO3Hflw3LDwUSnkS5CAdP7uMRWjbu64+f6eo6DKn
Dgb4lC5WuvPOZpXS8p1NMlFN8tirqEb7uYwHGfFOMEcMRMz9++A/ofHSwnWA
yTPp6VZK+ATsuC7ShgQAAZGhBGT65G6VC/efr7fWzl3R+uOBX+LOLr27ynN2
odCShAh2/pPrT7Ejm37A+K577kmaZIRVMSD9hHmpZobusUH7tDvaw7KGdJpn
PXSGrYBOGRnMnG6HM5285hW3hFWWzBkU21PrwMJHDeMWarOQ97kjGsTBN1ej
8CneAG2ExmMCoF6Z2VjGZG0UUDj2kej65d3kHDOOT93vDRXH+/hUzJgkTJmJ
muQrG3OgIZ9hKQoFfYe4AaY/cnWg+hlTr2MiTxB953/X6dGWt7yzH/Oi26mI
OFWS1o93cKVml0GunOQ+9FzIfxfaAGd6/FsnWJXZQpdT8CZhup0hoMQXapC+
VfC89m2g1Gi9AaLOOxNg4lWtGq2KnfpOURkkWcFujkTQScktvotaP0tr8Z7H
n6Csop4uKD32S8g7/7NYzdetgtd2tqQXXWtaHSFe/W48kEp7zgPjPpXmdHZa
RGD4oO2PLMACN7LgrGrUuklY3EmSeJfe2EuvtyGnzjP1DHs+yIecsY0cP5b2
JpVgHGzqhGChJ33dZak8V8kkqjcETTEx7NaX3M+eMLuV+K5PXY1Rgq0IRdy5
K1EZC1GTaYBEuQT0HAezeWtPA60In0z3P25xCa/wNAZDVI6OPfZVOH1gYy4n
RsWm0lZg+UAE0V6M/g64MeYMN9wxHmFsaknLdM7QUixrcWb2vyc651ldm1eR
qMqm81El/KXAMjV2QDv1qZ/pVmM33OYpNtHeZ3DwNJNOjolTCAVMISvhYJy5
epf+Nh9594dh2vvySGI3y9EVd6FKi1b7Sa3bJJf2Zy2edmD2twHS6VBGpYdG
Pb6ASHjq1uNt5VFESuup059VO+L0AVRq8FbaF3TM10gWnjF54xCJ/5q73wCP
v/zQPgBnxiGXWdGfdzQMhi2f+cPvBtOQZLh4Bv5Puzrvlh/lUVaUlfc6LZB1
xf+2BifGQqZMBTRaNCmmavd5PDfQY5Dh/qNsCTaI3dAVFB2ZnY+Sy3q5SSqY
O1LR+S6Oyctm/FKUz3bWgjssYxbynfYmk7rpeL+VximmvMAOVO3TVWU8fW1d
Q+Xb5DjYpluyYKqZ2coFsY4ntNBVF1Jy2tSj/ew2SBxFVk9LTXjT6yxxsDlm
Ladjwc8H2cYmrQgXh/DbHIplYnvHO5puodPaVq4CnemsvUx/6a5w9wqNxbKM
0QbTMMpr+mYcpNjq8wSW+AN25pR6sDv6tFHl980Q2kjZO51Se9NycOtdIF4V
QvDSHXT+bpUYyk70DpNMHIkg6e6hSAWah2R9NLb8BNB/m+zHb3NK4h3uf/B+
FBYayRBtj02Fxisfu5HB5NSSpfTpUujW88AZW3qY6cy171xgFOyPzoEU+z8A
fU9NNARWLgIxTJWMYyYil16UpRTTciDcrSiP6YVZ6MGLdJr7eIla0INSGwar
O9m81Klfczeuwb2LpzSDs1qfqvUYtbwom6QD5+Pl5AF56jzEKNao1xwzbe9F
Xj1c9xQOOxqwlDCbYlguuTlZn/Yd4+ghkM5SQTJWk5yCuATHmNDe1hx6NsiX
n01XMebmIPRZsfx4pmcf8mfG6WbfCxyf1u0YImJ5Cpdy9Rr7GHcyEPzz2VPU
/IoaApGkFnctVssYfiM5wCqNOFb6SgYCjdwYPAcsjzNSFLzuP+iFw59hluXC
0zLI8ybkANu6tESaZjnFCupgfwXX9DxmlKWqIOpi28QL9BNN40PFhdpIPAqP
M7MzOpTv8kg5oPyRz5+Mb9Z2oH4UOqTtQuAQL0aGjPBMDSiiMqOI8WANujPr
qw46fUFfBvQdHsdx40B/Du6XRdY/9qmq9nPhua+GJaMf/gu0cmIz1o4TYx8p
CmZcA8DZ8XwGvJ/quaZxr+YtgJB46TOvlQ/6oggN7ySCHg5t31saB36I8hEQ
CCNvJ2BLIrY9iKHI4wwA5/ttsg9nHGPspySVAhcH+ZRsJJR963APXcjwxUJ3
EZM2vCTptAXmHw9VnQ/dZ8H5cCvagtRZIR5B8hAhv5pRP6hq0UTffcMD3HeP
bmwPfdKn7mH68gTHEb9P1L7e2/HNtUnmYBKhXECz9WS6AoP7l4ABwf0m4R4V
R2kdFv3dJIsriEtihdfbsoHfofX6HjDBfJjBol2NxhnWG+d7g8gyKXRRdjPl
iqh0VvNNU9wpfNoaILU735pd3qSqyeOUNc7Rl+e9P7Y1kem402oiAo3xE26w
D6DVSt3ngnE3RzSeB1teDNv1aoKt14eGBzhaJXcDJ9zIK9ZVK3CoerrCiUq8
uw9oRjMs36ngew/yzuyPDyQCfT5vtcjQzOKxuEMct5Xdz5jBvVQx/+KVoDL0
A2KyGbp7MU3bF5MJxAi/nKLtHrWrj+ARR9k8jd1G2p6Ae0ehXKHa4wYI1bhZ
9EexWcJD/QrLYzNvRepRUlEX2I5GRm5GPw+deCFDYdADAViI01Vku7sONwdf
Lw2ZrF5N0KdFUJ9y/Vf5i9boeJzrftzzIarbznqMa79G+O7h3UFAzcX58sy2
Eg+o7xlAXXntGouEhQliGLWb34SBfsb90OIzCozBMb+62n6MAaDfrHfesh1A
GiwM5zCDFRMXxZfGuuSCGIgmagxl7VaXqQPz68uXUKDTDOgXnuMhe14ck1oS
jStSSb6LK1WgwJc4IxJRoor+n2WvfdjkXi/FmwceeEBPbMA0L8Gt7q3KwVWo
N6TnUOFxPQCmhOB4Ufo1845CPHLuaGRlTVPbC4M+hgiuTrArXpgBan3y3aZp
Byr/U2m9h9GlNyTrQoAFBlrmwGMNxVm7KJVaHRw9E2m8hiUdu4/f9NHf4kGt
xm2N8REtekhtU/DAp4D5xgKF9mKfC4pIp7kwroOS8wjPuP7XFclL/QCdN5jD
BIjC2YGA+RkdMxrFB2ukMukO6eP+6NZYjBVlvQBGYtj0/LuM1zJ70+f6jpIA
YO7H/Pdy/3+UT5bghqMaNcnfQr5HEXdfz9d/NQuMKco3OVR5ptxEfPQxReSY
r1CY1D7xlZo9zFpNHMF1A4s9FnTu2VKVX+DiAu80Rv6NTsxrU2y/UyKyn8zO
QGvlZBYI5Ev2U/ag0igvVFVhRzjqsUJbdhYf14yo5ZpsK8TT6TwtQt/dbJaX
hS0TiwOy8dJhdxSBn88/BEmERjBGu8AA4sb5AjBniUGaFdckFTUngsTUxZyz
VNCdXjwueke1kAJdiONe4Lbo5gx99zaABoAsKzxRTerFpayDV+qtiUVVU+VD
wSVMpq3fc1h6l9MANFmkWeaNnM0iNJBggSFeuJMPgTUh+BCO9vZ64l7hHKqp
cEpJVWgnYB5jnaFqXEL5hVxh3HV7YiiXkawg8VCN6k5ObMC5sEKJQ/QG4/nZ
7QlO2EaI7MwCX7Np92AKEdw+REWM2gSSapNUFUI9WRAfkxG25fsoC82Y/2EC
UfpFLOYn11l89b5UF7WQtk2KaMxqSLdLYuDCTysZgX5D/zOlR7TocxAdFyEQ
WEsuVhxTci5nk4qSlJaydgHpOkVmhxRO+hDYp8L/vrKURaP6CYCbr2e5bGiW
DhCGdSzsUNC5QmKvVPtA3kAnXo/NHKF28gb4vA/ue0WOWru+gQxbfn0aisYR
wrZFG3MFCPKYnLQCUc73QzIS4wyMwZaq8Uxnlf1QJIW1HhP2WmlxrlJqip5R
mCwG1KAtpmVcOlOrarvO1y95SZiDJ85TL5jRX7cVcbN+GfIbE39nowmyQcR5
ZL4M8DAg293ZXjeCaX47SXCvn8vHpj7xyG1RdpShv7v1LxE3jQ5G/WFti1pz
xra/woW6NpTVQQlWp6ZucLzyt1jdb0R/+h2WMuVgnAVNAuUEVXtRcKyQ1B5P
eCoj+cucf/BNoWZiIxx5TBHNa1mGBasiKP0p9xHkmJ5EnnmjPV+un/OU1PSK
+gkKW88TMnxoeL7IMK+Vg+lbKkkgamUVxpTj/w+OzV0I6sGlwpirFFrUjisT
Sgu7HJyPOuO6ujIF2jRn3q25YkjqNy1HY4fJK/T/ZOl+G9BCJvRKsT9YUMPX
/GMwfJgTVeb6gl0pDFuu9lnMExvo6v5vuhTT9+TNibidosjj/sK5WQQo9YOZ
pCUy5W/1fnJ1c6va2lz72YR/d7Q0hnEgn7b8JBZrgJ7lh4Ir892sXxqR9cuz
RHzj/1vUw15HXcgnqz7lLWWrsOwHHg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfRtKWiwLrFELBoWZAFZCKZAVTGBqi5v7btnQDRPnvoZaKlOaEN3V0cLM89F/MlnV6H0W6F1pyKDgUpBOgwMu8rTLdYZnnEUCfZsufC32H8C3ShpauB5vCY2BbJTi3/6F3LggqKb3TtKq+yGi3GNPPvjOjQ9S23nQzVC4Gm3DXdQkAUSNhFYUg1/2BjwMkGSx/5bzJ5+Sd3A3TxJ3vtv10/ClBJdgC51FIdwgF6RVUbM3mLB8/PfBtMg2NjZR1uJni4kdq+qigUNadLVJ6LdJnlfwVIMfxWsWGQRPti5QWpjiw/IjF8mH9I/GqhdLLw2/SFX+4ypBpE3DEBU76AdS3IHvtd1NvYl/b2Wt2rvqRSEeruqbWXT9Lu9IgRtneWve8wAsjyi7OB8sec4ymXsbDL+vboZDCG2SvJht5DwPQoCIF5sG8yhN7NJMXBh/RW7Dkh1Jls7gBOaWd8p7HUuAAk0bJCT77+G51l1skCAIeIjdGH0TOhDEGQTDn/tbJLjTiGgJhCZ8vankWi8SgFP/QtOozLDTyDFoGa+o7Jo/Rh+1rPZy8CNLDidpe24ZaaNZu2kknRsUE8haE0RLcqiTvpwo5+0p2NLazPYTaFHKVN8Thmih9sziBGVCNklzIeb+jJqHONyGdiOUnpjZXKHfJaozUXiU/jk0s0bWOdX+GJDp6oRaE+IQdcq03maPTcHn8wsNdXY5WMcvi+tVBfckt3HTXyjk/yijjwPCrOKkis3TwktpA1ot/dIp1MEzUl6/yRucCu6hq+XZRp1rOtmuWvq"
`endif