//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YcHSy1iMomjibiwQswtQzUl6asrdIRwTYnCKZD0ArPNVru8VODCup56SNhkp
/EA/Yq2oOMjFk6WRI8fHWnqB8M+YN865jIYLeCW96FM3urCGZnx6PNA6DH6f
66NePbX4uyfNyPLhE9OpzHJ0gxsWqB75qAtWihBUTVO/9EK8NzK4WC862Hpq
TPpRHJ6y+GBuGElfL8pubYn6us9DotUZWOeJokVtUsDzI3xwGnfr0jPjSpsn
WtXQrxL1lHg+iymVWNS64j50sLLCmH/P1YCWqnOdypK+xCy5wHF7Qt0mL/bT
wdxp0vtAGO7DEEDqBkzFNW9SbtGARNF2xzhUpOhgNg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mAio3XpgwJu1o6/1KtFnQDvD2aMclVnl5hD49qf0wVoOG0IO0du5BNHD2LSG
njmRaf5JLLYDp0VH7C1ODAJfLzbXBevjK2axRlIbbV6ULG7R4Qxf/CUlsa0N
nKXT4JxETKvKtugV0iNeYaQx/X0rFAnFUv8BT9q1RGvRw3UkSJ9Lg8t6hSAA
SLnLpCl4SwpuoN6AKC+dWpw65ataTiRF5atMUD8ErorT4nN1uzs3tbV/DQbs
pqGg/j3cz9bPmoWkBi/TdcEmrtrRX0elLseh7JT0NQp9SmAy9UQecqJaqQdn
57aYBgksXsP0JIMawvZH6kZRibtN7xsFzTjWFMWoVg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
dsHiP01/DN+waqQi4RC1cZF1VBcNCq9/9Az8h+6iJ4tYMmdBXZmYdJYKsoV0
WW72mizpcQeGwFLFSIxaXONnGW6IZOG/bN/Lhn1Ohy1RrnuC4dD3M1BZSIVv
EntEYcEA5M/ytMOx7VCxJGwcSOjUbK77CZFmsVLaEQJMco+7VmigRZsdELlZ
gdRVmY9zgex4UqxqlASecdICUnJz4EnUvvRHIjW4yErsZpqW0VmWeRn90Z1F
Du062EnWkOSi0J6QzKnRloGArb9UKAPBkhrMrP6sN6DsI7Pc7yDt4r3idW1y
cU/Khfj3rQQXjj/PWD/OipHnzS4j1pggnNUQbNibWA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gczc0bqV31tAo+QV5ubAm3oVZynxaZoPLBpiCAivM1HkkVE5IOWpvjDkRvgU
LHwQcyZ23Ta77Mtt6+i4BQ4sjFZrz85+xA21fSwjgqNWVzdhN8JOzQnfQ70S
z76o/FrhmOcS31i9iReWXpg+fM/2he+j5LXw/GAGs9pGOU5lBfg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
IH0Chv3oCxeORLZgJwiH7dcAL788Ei0uBuyXxjVyxh04n3OpaVkwkcsXr9iz
NXLJb2dsKbrIOPggR3YgsF9gXVLeoHe7/LLAku0xyUaSdQC1OhMlVA4CSI6f
0ojcRaxMI4eu/GjNMfG2jJh8rUJ5iAGmEpAhGGLaH2DIPFb/Sie0InWGljVL
GKrZjQijm7WXH4O05HU6sgxrRA4BGz+ZBGnmM/tmPlqhImX2bEuDL5Vyn/jn
3KMSrVjxgaPnRX/VdWdfQoHmXjrAzR3kzXToFfoTj/757rAJ1WkIDKoUzCHZ
x0oPzxWOUppcb7KOYe5Tl8dtDRGeZ+ZUkl2pXjKVY/5tSvaWXsMAQzjsoNdS
SR1ZONkfetn20XGHi3dCFSx0K43fT2m60TL/KZIDhhy60GffpeJn/TkkTRYe
93ecF1GLFUod2GQs4v+m0n5dNen/kSmhS48BPuFurQ3yqaX5uhs6nP/yOuy6
M9u0aT/YOPB4f8DGghV0OJbksZsKUpxq


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MAOrKTwmRXQU9OGiCCzkRQSdS9BoAeGxhpcq03cfslZg/CqyuE2a5D+CR0Sw
wHTytuaIOnNw5EcTl4Zw0HpKNZaK8PoOpzh282UK7APiYD23W3STs7VeFtr0
1p26NCeE8kfgi/5UtnvTgOQEDo5FenuTR8NIDz7er6Mx3LB0WeE=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Yx2ohqdpxvHC+Y+sbW4bjfYiRQc56ZmPgs5ZM3fhWtUH4sczhncxTbdXVnlF
o16IB3ql4T3mSHgppgyCwareFOm1zTH3sKggdHyK//14K6GqIc+hPAHrJfao
7N0AoemAL/dj1TritRgxCOzHlCX3MfiN0/cgr8IKMkoakHdU6OA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4912)
`pragma protect data_block
sCvLKHy3jl4hbDJ78VWw0eceVdglQDUdeD+OvmIhECJ/BZE2oAnJR5ADc+no
ZmQd8UVBjzQ4SFwhv5LkH8lCE1B0KdC1DNscN8aY/NNP0GsLp9kUavtG7B12
4QZeuz9DKAaN3VP3n3l9JwLc+/zQROh4jVftyPW7f0/IIOuLAQ83cndSViUQ
L9crKIkIkBZNij1Tm5MfKvTFs1FTzF1FaugNqnzN3lkxtSxnSeas2Dv8uAXg
FPBY+vsqwVQZKU+XuCaR2fb1s6VNUcLtArtcIy26WZ2I4DYaxTsH1dHFVOna
eSQnqxUHgVRI7XonF1RtnYsmfkGUsPZIIh5rpQgytvDXhURiCfgqVo4SNR5X
70DFlmmJxcH7fkQUVvAbI9GaM6v2yvHATHze0ikVjs5wfEr7VqYG72cgwsxk
HeRE4yM3/o6Zz3AjzonPW/BFNfLLi7avjXR7Kfk9/4Cw3WGNy3jFKwSmZ72h
cvVUsekPWe3jHCMiE5lWWGcyYYGqgczGgvPWCyUDPPgnlyY15/i08Lkp0ffY
IOPN7pHzsG494z1LpvGWEb4GZzRA4I+hX0H2LDjeyMIyyRmuu21+vK0CmOwA
IR6cybzGvNFIwctzffI41tbKX/wVYY5duRhez8z+wGQivMZhH5urT1Ukx8+g
lAWjKCXSXQvtTksfrxv/AGawyFeu4/uOvgKb0rjaJ55/pZ4iAo0GSYvpUjSv
U1flmYIWGetLGhVMJJEsoM4e1U1lwpEVoHQG7vBXUBCQ6r74ll2YOueSoiL4
ginzc9Od11ia6Awj5olEnQ4Ei3248eRB9q7nRkxaJvTR/GiLNx4HLujn42PH
na0LwbNOXylcdNgi3iq/7RHKxZpZJjrROeI/szHRNJTM2GkDV68CMR/Ov0Pl
hXeGGr04pNvjxI5LLT2+sDBJL4gPaVWiXo04eQPaOXbEpbgac/mNYS2sVm7j
GG4QesBpVc9FzNFWWpfPlyIhg1wkQy++uowqKBLyxnQoXxWFqSSs9sMKz2O5
xFQvZPLRSFVbo5h18Zft+0VQWTI0CuAMEBXx/wZ+WsESm+4Ac6crXmQtf2TA
N/49Uu1vaDNeei7jiBddMbwp2Djk+z7e1u0Sk27r9MS1K/IdpEFg9mwzuW3o
QAGaXjRudXxsij6dltLs4+hsy5kG9NxjSKwo9vjerDBcY68lj10Eq2af8zNr
oKF7YPOh5WE6r6BoAWYTWb6Ls5YU2AVmy1BYs3kV78AU9ml9OuUU38cBn4w/
KaXPjOzx+9CK6DTzX122X8+uXudT0M61LWob02fUYlWqQ/eqxFx/vrBp3Nen
y35FdtUmMeti7rreksIPQijY4b6tbnrkUtPmQCLNpQrwGgKNhoI0tmaNS1jW
uVbsQP4fbfvw2ZWRk/cF9rFCH3nrLwLgJEbsF2falV/b/qmJAf+EwtX2blfl
yAtlOLZlvllRCts+kbTw7j89rTN/p4paHXX/7mj+QL1quRRliyKQs4T9HGq+
AXNGGukEznu9m/iSFCdZdZlFvrOL248qMHSp/FvWuOzNX8NN8mo0+z7Cskzw
Dwy5lu2j6hUEHWGosFsUho4rjrlyMyZr4ra9GOx/k8xu+368FAoXC7yJ//dj
gvImWVdVkEK+Q8zhCo/uhctJ0wN/r1RBESNMTr8hMt/mv01LCTE0RVr4LazS
Iiq2U1zF1aL4kuT5pn20bxc2qn7JnTgcYDDho2FEWpHRpgfmH6jKw6hwvDx+
yen48sUp2gGmHRLAj6ZvzmMtU7KJktXC5Rkw2OQ7Is0RIjDiQ3gEtB6jTC+k
AHasIsP98ptsvJdxhcrQJmi9lcO2pG1jcqkzgxRWRNDbGdW9iXPIRP/kMl0i
FFKsObYJlANZqEbHjhmrhUou8rupVn50iptNdEeHpULk/JwzzmYelBti7EYs
dJOBUqnxPUsXfJV2gMO4PZwMSUyTjaJGc2bAWH+pxhAZjEg/6u/HjrEPA7lQ
RZTnYV4eP+jdsWyXnVqvyMVeOxP9FW1F34IYXhzDPOTkQVYRuxMPc2SkJgZJ
9kNQYsi3sbyReNGsaFbaDMnL/1kWdORhtnmRlLIf+w0n5Cbh/JSSHthkGr4s
zPJ81l7S8oz1CRFl9hDJ7NWFvP+uAu8OWnaWNU8u6bUnraMsz8jneeSS2ZWy
5p4qj8n6EkjHRV//CCUk0biwhXhH4KajFcU8CcF+LqkCCCcnWnC/OVkWl89f
H2PkjQEHn9URaEcHWyGSoFzXu6UzcW6M4HmIc6POAqlc4DnjapAPidOSkfw1
N1e6DQn3fiq9lrCCbVpp/ieuG7+VO73CdAKHxutkl/kHTKTz0jvKMvgFOBXH
1HFXlTbIU5pHMs2DkqbiMQT1UR6Y4aIRKH4qqAVZ7DhQBCKQr+hLETJyt1eB
v8O11hN9pe409od/2o36te37KJm0D39CJMIWS+qsqpfUvBWmOgUyFtEjs3Yz
3J9aBToYPvEOokLJY1oGTCI9rEHZTQ2JaZyUFPjOkRr4jDR07mCW92+45QwO
LC/s/3JrPTTiFch/V7gXCVh+GgTwYfW25Bj541ZDYnyBW4L/ZftdBMMrsW0I
29Iq1YBaFo/z2q5RWJsWyvrmpP56DjlEXxW5jOd6bvuPCA5igKcq3CMImINQ
2fh0EzUPLJW0rvCRYjLzrZDM4afqID2U2Bw4xcTJmjvhwNZ+daQl/x/8/h/Q
tIRJ5e3FlP9QIfFB9Heq0u2rCjAyPovwt/fKk950ZrMAUtmLAtEm3hx2DBJD
y3R4QV/e7flLGE7eSURD5P7BAiHUiRYsdfRQkw3spac549gap+foC4nr0+yO
TEDnvfKLlPI8zT0HthNYEFvWP/qWju/gof1C+kyQ26gPPV5b6HU8bS/nxS6H
8nlkiGOe4Ha/zXDE4ookpggIatQJ7EAGb7zYMDBP0tZJSBIisSGgmJjJUKpV
MpgF/YMWvlE6IzBxaicJpy/dbu11vagNOhJ8DQDpna3Zz7YLSHOh2DAr+izt
UJe4yLLX6KvmE8MBttFvyLPkbh0GJcKxgc9yUDr4nGVkeQMMyNyd98ysxOH9
jtrqna+uLb4DnfeBDz9zEkFKt/VL7Vk6QuJhJHX5JIGNyZ6LPeg6k/zXV1el
gJ3d0kmcgYsSGPHbW9iD/flUt9m9LPIJxl6yDFtf4dAYjhLxmzAh+ztkO+pM
Ds7WCpm1DIAaNt0vTsE4mGsHc1iJ6E/jcrHEyVLgV6R/o10QUvH8eXWtPpNB
ybfhxAl2gS5g/gTEiVE++pHYKZbZl3g7J1E+LZIaxkkrm/eT6Ai8w9QzMSL1
Fq0p4nUop3IJnliRJLRRSWCyon+c90kzuRsOe0psRSnAF/q5+vzqddZue/t7
IHJkBuOM5MisfnPEIjYwcwUCQiJHAnJJIa2y69roL+ubYLb6WI0Us/G1eTvy
mfPlrsZ25v5c1lBvf/QrGZJe3+p/lpZ3vF+/Qo9jEXhKrWPxcBwGFuKgE35Y
CAzOu28d2f5JBjQtSKpyJNWE0U9wGpEKelwk0dpkNtpwEtqy41+Xgy2KjemG
EpgMADQYV0xbPTvI5sm1hsUno1lF4seCxSwlfsZ7S+seGvgPsf+auT2d3+Ps
jS0qvxUmezJx+rvUZYkb9lZjsVSDiwGnsCFWBdJfxMKoIOsjgg7Jng90s02B
rKCM5Ivb1j94IbP+OIxbWWsOuOCJM7ZhSUPbtBa8uI8TJuYPN3xf2PUUT2Pt
YurVPIN/84RO3S0qe0RUQLbjLIHkCUSAt5RIN7zLxJUo9ttBCWgtfiYWb0K0
SI7ZL/DI06K/Dtm0PsI+kHIllkbpPxuhamGQ/LFRvo1UJz8dIwpzmuzLtM1d
LUdZEz4qhhgsrQ1c/oyJHAogsAd0VMtUNael1UeksDZ6fpPJPI93qsKkWEep
IYEzXZHUI9lD9orvrSuQFqjMDxt6dB0gq5Pc0W0JnEOnlWy/t3gQTdRPDiNJ
yqHjjYAz4MKbz2DmmRRtU/htgO6GiFjgrlmie1Rw4OMsNEnmUOpnyhZ/Mb2N
VyGGloFpENXNNdChwtsJq2rQR3v2ZK7IfwahDF2iBDrADeuuLIynOoo3naIM
VxxzKBtMyTAjxlwSYvcPXiRj0eNnXPAi8x6UuiothZuFjHuEY12tBm9JO1Ft
eMWtcCDGw2ZRNF3Ah5ZP1KSQnay8hVj/VRyfwMAszA3InwN9cTubhjNh+Gkp
PafxHw7kZdZYC00+OxrZ+xnDCgRozkpFcFGEC9oDJr6SzESr7F/Hzd03Gw+E
pTu1SFLMiSBIykXuIc7BHpf7b6h9B+Cyjn7yefPpKKfh3AhO9y5Pn3L74Rwi
K/VwWncYLHbHiaFr7tXr7GJFzRm8It00UBhW6ycBSD7jmzo0jUX76OWYbfvS
BZtRCCciuQpvh5PE+I0Y0ErV3r+orz3ofY++CRV46xxXvZfWq2AX84QBkTEg
rp0XWrttAm+luMo+8pEnEinlvfCtCUuSWR3IPSTllBHVZ4R4gcDHziyjJvYw
rM1xzu2hYViSiMZfq1gK29YiRnobxFd74/Za6U7SGmh+97f7rAYmRBN9B3z0
kIgQqJl2mkqRnOv5Zg79X3plW+fQRAQ0ZjpOwKBvus6MZu1S0I3uYwUIwUBF
9XiGkjsmfXok/GRPvQad/PrdVVShbdta9Dyj/zbKru0JRR3EgblN9K4lR06P
Ecy2Cx/K08Ly5QbyP18KO6b8Q0GdhA6jmyv8GVIeDB7uPxPGPZx1P0aY5q1V
Ys6FLDJBqeIqflaXh56c3NbYnKTIFiJvl5X0uCoYg1zUxzQWvCd0boKMduiM
fP1Vv42Kxj+Tf9viFn8zKjK4/W/7ASdTjlPfhMrLcxjmnyiWOqUuS0eQsh5t
JDv1jw/G8zhbPNBW7xLJExpm7nghxpa6wgx3fhpEo3PCK3YH8CJJxYhS/RjB
OiNHxS8TJBLrxCT/io1HxMw3lmWsWRE8FSkp+RPMCpDxjIphLEKLyEISXB9H
CeFrU0zT79LJlIntg6/B27NC4mNQg78pP/vdrlKzsF7bTdVXzAsZY8+JixeE
n+23OnadlxxYnA7GXjMakfPjQJQf+kK98Y2xywqcdRGBagPplsYRSXzkplBC
Klo0yWrZHPjXiUUtYc91f6jeL1ECJNP4wOGM5fpvE/T2Csu8PMkO4VpnVRk7
waAQKwzrFduwipr/dZU36KT63c7TrpSZNtuFk940uziFM18zMMP97UWtZ4Q5
gQ5GMI8YwsDvo0kAi+59HvMtQKVH7ShVQwek1ugSZ4MCaPT/pPi22EEaaeML
wNnU6oy/0ZIWCA/BoCDzyALgWtu6oojAzgGSOMHzc9YFjCffMPAUV5aM4PwI
XGlWYcMmhW+CDV1fDYnZphEdQ1RYXVeUImAT98SIouIccg3PH8EzEQ/eGCTs
LvL3+p1DW/2oeCLm1spkUgCxY6OSziIkEUgN8z0zz4xO8j9q7821Hb9ho6N8
tlkJ/UBX2GrycnSEzBDlSBLLbF1F2XlgojD4CStPNVkBPAuIlqyKdEnwDbZ8
7SucvffZqnxQxX9/NtvBsTTNA2G4HJ4o5dWb9aVOTBLhMjKJixEUCGTOstp2
cMe6VKVH5+Ykef28GEn5qVyTUrEE2yVdx3ncC5ctM2vqESFaxVL8j64cLROM
tMBAoiqgj2rMnG1K+Mhg+r4/Q5D4iGIZ8K0iyhV9ytXAdCM+vSE07ucAO5oJ
iMWGpimf7YhyoYHM18LOjdHi09dujbi/ikUVKg4DBhYjqwaCvEtJhUcgIKRI
evWPZ5VDHGJE0/d3m3MnCkCkEJjER+Dr28+BXZx/mDBEoa1sojSr06Hq5Wis
keHvTb2VsQd/1BwtA+Hl2l0cPZxmP01BmJFWt6KRu6YKtVEtE295biatAV1o
VDphVd5nHmNnMBC2TXAFy+l8/p6+yT+x57mXV2NUxfQ+/L7sx3/V06FgvTTs
kKRZT9Uu5GbhTuBWQ9MXn7kx6aSYqP3/lRBSX6m2g5uW0nKJa/9Z5J9Lvkz/
VOGC2RdV7lVXuCXyW5tw/WypQiejTYC9FtXM/QHD9D/y81pp9xCGtiqfDv61
GZYuECE5y4rnyqrg2gQWk2CePSn1LqGc2Jn3YFz0o+uc7+3ey8SPCdqR04Gm
t1FOdFJMaU83CdX8sqtCriKLpaV5TM67GeD8DbhOWSMd8CWggsxPPJ2/B18+
Yyk7NTUEOzhFbHjlBUjWvORubcsjxMXqqb+XN/GgkH5JbIRyxwu9dAF+IkT1
6dE9ErUF5X57etn8+i+QNLhNnbJIA0QB0mICa1XQA1PM07NHqCl896qERHK7
H6qcucJKshCJm6SNlDMX/ZckLWpi9HWvJiHiF8XsXANl01+O5t9lvlh2xn/F
KMQ2JLE1dWufy/tl4SDCqgkpt/HxwZJWBCGVOYstPCUrr+Wz2M6eDP9LR7W9
PiAAz266GnJ9MLPvq2Zuuu+jxX2bPIqt8IqxSTAio9DGdtEFvvnAb2ale5Iq
5+Gg2bpH+pHLu4OShZsdHPzUCwQMQHxPGsDv/SyJyobeYZzlvF2QaJoMWo31
DfDauuuI6Q==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+kzxBBDen7oxgPd0cWx2j46LjER3nnxhzAThlK0Eou8rfosOWP1D5UpzBd9qKUMPWr6h7oLvgzs5Epj2lej+2eXtICCjaYpogCt9/0l7SoNtzVjwh6Vll9KNmhO0bUK2CWwtCRuTJvOQ/LJ0phrlRKEt/OmuKPgjrLd2k7CM+emwmS8Wxf58G2jqicmJHjR5oAZSEvmXffZ6ssbZVrNiRvUKNVkk7/A2MfVKSeShYdi1SU8d8yQTVpMWhopTsvT+53lMSWRwSxonN9jeDN+MvCQMikGhtPDJMmRCSaQf/snOC6LgTC8UffdUzrp8aBo2ucCoBT7wDncQJ6E7neC+6k3jAOpzYyN869hb5QRH9MmojnjQms5f5l9zErq9xASWMIqZG++hO6xyvFvoz2CW3p65JeJdoStI2JwXIYgSaFq7Zk802I4buXMGNcJdkvJRaj7Ez+k4Mmoc8aoUYPy2Q4ZyUp78Lb6zqZ6HUTzKvbEwdZWfAUh/Ixj4IGeW1vToE6EzX+VqoD5Z8XBwlbOueZ+rCjm8538w8yofdPO/p8V0p2y9vZmRJyPQ7L8cq1og3LVvX41lc6A9v4yOQPEkmJjCKhg2I4ymD8YKc+PvVbmQVdd9orBxbJ6XsIV9bEXKZQo1/BjNnp4uL4aL0s4t2uAPtjlce7exJecxOw0inibnMp8ZAcGPLnc3gZWE+EIs2aHBLIhK8wz5BWyBKKD3AERzbxh80MzD2orh0bJyJW3CvbLghUxvsCUPms1yk0nVQxxXTt1dBqNpCuJeMtHo7yW"
`endif