// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XdgcI0VJ/wNuYWPr8is19BCA6pDeAZieokxFVrqcIozujiLXeNmNorD/N++N
y+1iq99M/IfKqtWMJvJAb/AKNyYLOwDloeVF+mIJsJuRU0Xsl1kDN2Kil5gv
GIFGUKAm5KhTcgf9Qzs52nn3AR+//BzhaJjMXzgSs8/7tJv84BodyPkSGe0x
Mrq5tdS9qkhqWmhd71Qjoyata37E86AoM8X6WhFfpW19+iky/3KDJbWB4QRw
65aIL9aB2vOgvtQfEC0GikuvWZ8aLIHt2cN0VeCJoQWMm/+HmNfaq37qjwsD
BiIslazyppsRq9ZkOMYmgxK7eCfjysxzjHkmJMIsaw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
ahDZLf/hDxkUD1arFR5LJwBN5r3yYaoCBgyWZeJ51PPCAIFHyQXU3Z2M7HMW
qgdOIWxjRTx85lF373A7jGUaY64vOEHnM5PByWb4joRAPlmwNH2IZiWacvrm
TshicUz7nTVtK6ETeFs0o1A64QTC8x7aKGvNDlhGudCgP+iYUPri2lPulemU
uwB/AHpy6uRdJm9d7X2qOajcJnPsg3GULMSBQAiuJh/lX1lpTSNi1Bqh7DP/
L88XsEc2YGYFFadu3TlmvodDQo30Zs+zePSdWoqaZ8e+gDIFiT8iuErmUAg3
+O2QWKDH5tk4dGvFAz+aenaca0JHmOG6FCWMii0WPA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Hs3iHP92hTQo7GYMCUIohroivLkxyiDaegLDfu/4yuYPl6VJCiq9hybipz5c
PhLWMwwRufE4QXWlIR7dze8CR82N+RXJk23nZWbEl2RV3CORr05gk0VMx64b
NTmilMktaC4La2sfqs7d1NJWF6Iq8O2xvRAXBW13QaIRGPdsYn0Gd05ydAKo
6g0Ji9+WZDsiDLJ56DqxH6SbuB1XK/QfYHN8ta5uKLFIPKs7vUu5VDxvY0ir
WcMwvVaOSkd4V0jmjoQgA0endgrbvmNlhaUzXa5A3MMqfiDxXho0XgcZ/76h
IfBpM56HKh1jnhGroVAGp/p2G0i3b62ilW0XoP9rnw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NvLXehv/tTatTUjc+uGE9k7u0lh5YxIqNLWvADFXAlm5n3oCHAEdKrMDICdZ
lHh+5WJwLj1Yns6GdSoneWZM8qkA9RWWYA8Dpm5Ect4DcJEHgVhDAWf/lDxi
iKf1uDHx3mWWRUdAEFD8xp4reBWCPUa79nI794eXMMBPOF8gQBk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eeUw2dfxIFqnLEHhh12woT/YBgvh04TPtbTOnaWz6Q+Wg8wTwwIebjW2yirH
v5Pzwxsp4ZRN4KOhruF0rrMzaao6jrTCC/OJUR300LwD/EdNiJ0XS161KTgr
W2nCdmoBnNeoUNIChUqPyW9gIfVqdzBsqr1MFakGNUaEtU4oWkiH/P82scYB
RXGF8rcm4ILongiPNLgr739E8s2YVHZojDN7R3MThlvz3+0nrXlIgvkBqYu2
UAvISnnPZbw4bYBRUXvW9r+hKihZl2SO/3+Oby38WXNpU4KoUYSY3oDw27RQ
Iwi78XtR66ciIwVjQctg+Y30WBXAd+vjSz02ZwnWEZMKwiOV1fj7peVzsLTF
QW0/+JO7MfSJHY+7iImOk7b/aDmymdjshICelj6+sM4Hso1Ul1H8jNVMubsp
gRti00yWTAR0/etZ+KkVtm1TywWwwZJMjyCcZmgE5teUJOaAAy2ogzBLo2Cm
GrKEXoreEiUYwo9bPJXy0c8l3kb1bRwn


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FHeNLs/Mzm6WvXsPBZlGHm4VYnELJOrFaXXU8p/eTsofKlfKzUc2qjYZ/Ikw
y0rAsRKU/BNAJagNXqP26ABYz22T9yWkP5Hm4WN9x4foY/ELAwPbxEJfTVvS
encAjq33UlK0lA7UonoK8JGiRe5K09M5JiyJotRFPDJqtGzAsmQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
IeznJjDn2orhEj3elEUIecLVeSlKgwasSbpqJpw1NCdEOWwETbD2DTSfmDHn
PcP7Xji7p7nmRV5BZcsrjWCOydOlKeUY3LtZiqPXq1dliuQ/pVlRcMbPb6sn
i1bsYHh2RW1l4NBa6vg+PwmgxuYXmPhrFoG/s5pIZYQ90gKn3+k=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 153680)
`pragma protect data_block
4GlrZOOMNALS82G40qYN5kwlt6j5haLdngBFK9d55j7v/hMv0itKFeMcMIfh
8m0o9SUZkg7JKAIvGYRcpk10RneHurTHmEfrhBro8pjiULI34evwDmt1gJVd
6d6hUjS5S+O1eW+awWWHgJvYAwLfwbdM3niV+aSGjnBT+n+4Jpay6HShoUeb
0hYPseTx7ih4i/ku8NLFee/Y8//dNu6v79kFO5jcDCCEtc6hVOehaybvNUVy
zZeeN4SXGsFq96DxFLgMv74qU0QpmRxLKVQeN8+KdhdQspedWcXWQCVGkvEQ
vygTJN5Jdn5oRpAkhw+GPLQHaokppJPcuOy7gCb/3Lr3RO64bHS6W+oZb8i7
GfZwfvMFRqvAhJYycOshI95tpXrJu86NZj+UZ+lDxt69MJIhgukppNoZHu85
4zaLXNNh+T8rvgmCSLUhWr0TUq3+GjJXlkz57byfu51SVaUJ2s4rwlVQaPcI
RSJxJMoHPmijSGvke0tjB0RFeitoic9j7+5AYYjX5q3FCraJo34D9slkX2/J
m3qkjrSrSCnQCnYGEd50HCEJ9ZmuZ+/cjxAFfqa+bjpf8S4MbbvRwkTRqcvu
8ZmQHjDwhKcKivj0UyC2OiJvzUcuIJnMzYuAeASL23MI2+yTwAC1sQls0Tsl
rVRmE2hG4qhdRb6GS4RLhsjmAVopc1Gl1ooEGAzptQmcKqDCAJoGMcWg110g
k/H6ZCCD14rm8GLfB4z/GxkbhUIENQWzB5j622ax+TVMLtobdqjL+f2gUyZI
CAqlfQ9al3cKTOszTyMAx+YVV19I/llJznnsm/qMSKp8eRUL0mCcbhzmMyhe
qmv4lXPfQrFtcYD/75uD9FFEWZ85ksZntggOMS4hraXem970rW+shl1ur0tW
aCvVRzcXsIf9b/+JHvy/FMrjZMk88rL4tDl/QtBHlPRPJ9N1ntl9Cv2LNIbj
4bqHg6pzD6whkvQYnQ9rRfUbQU5FKZBsj22PAUZWLaC+EltdpD2FJpyaExTH
yX5BGesOsrslOeWe1OiQBl7q/HERDJ3YOo1RsKuWx3oBjw0KnYbuHgfkaYl2
7hxBsPC0ayQrcuKaDptceGGTsAtcnsYQ1a6uFbJLv2hGa7HdEYAE7rp3+VpF
bW2mMeeq5Elb35lItjyaTrSzXbaEYkHERedFEideC+FAHM01+pnrW9XFtUbp
UEbgFsPNCTmSPIqNnoj22O6mFypNaiyXiAoc9cEtaCs3bhgOGEvPv5pk9Ok3
rpu2AMFlbgQ+a+yVVVRMZovMIl0d9dzsDn5/vEJxeE8BFqErx+kAoKkxhz84
MkbOARIXrHZeZVT3WuBeHZrwUt1M+qn/CgGM4bRF1TgOfqDazBDdtBy6mWXz
dovECNaWsmrBZ9SX3Ard3BBNbkVQGwGmuGi7FiPgEL08bPEeokfQSB9wYfic
vs2TIytqpL7FLDFtjyh5GC9ldJ3w2qZmqTDW8wURmd+NBUjLhqyRuBdDPwEf
dgpeHKSGC6fYacdeP+GTT1SzX3iyIBazVxYrsnpBMPYejxmp2PpvHdwExIF/
wCEuMgm8fGWMQttOsrxN0u84mWT1slw8/9jHVDELFEtavPCR4o/28lRyJ2CB
8t81/fjCBQ5zo0JALO8QyqG7U5u0vqQMt51mLHc/psYPEbEQ8+/T6GwvzbcY
yvxTUehJj4U5DO1vSaRXHJNqc3YslFeJHBBjQAuTCjR+B0GUa4ZG3m27Up8t
a1KZRJREMRgFzp+WGRmzF7lp0a5vbvg7dp1/owqit3txQY5rM9biBXB0btqQ
BxOmCvQB/OjqZNvbLfTBWq70f80B/ed7Pkx2vYv6u+bOjcRNIXDBs4y04QJu
GNYCjq8ErYLoLuCCXqpD63Mut3baDHgB3MbJwkWViht8LVrqa4xkgnYjfLPq
GSgGo7Rkpfr7aC3KRCvfN+3ozEsVMdFJ9WiuNqMUrnyYgme76UGtqqsYrMYu
Laz/aU3VZrUim5jAUew4PACG5ULnCbJoSli+IcSevP8XThqIkoI/kt9oqBrh
YGJ7BZW6ahqTtBhNuZTyueHLk4uG6kDMn9Vf8WY+ZWW4ZatDZskEt1wacPCM
8ubNI7FJ7l4B19qdL5c6lTgomDvYpBB9UUXsjNXpPFD58kYWcyOLiEvaflk+
lWGpkBqy79x7YwcYAez12nKH7VRXKYvCl2pcJB/aj7bfYGdcSA+dz34xfXym
pVm0mf2ULDWdpdpUQ5fTr9bLYHtbHbfssTi/Oh34Kqp8prFVG/dyxBvpMpLV
kWn9my62YevzIO0FKkcYkrhzZPRHYZeLdREs/M9nVSHtjjlsGxpFhqfThV+L
QPrG6ydBQ3UKPmkdMdEbeBVqIqAh7cjXNiQPd5GfZUraKHZjwfY/o9d2KX7D
ii4EXlLkSaUU45jtminR9nLJ6D4V2+pGPYHFL5Ab7F7Cfm7W2J8jd/FDQejm
PJbZ9MXxb4rDmC2sFjegHN4GFt3mU3WkrGY2YeKOoOVVs+3PHFHJHFaIiA5f
T6Vh6GWfiQn7bhns1seBfbs83dkIi2ckJEV0s2wyslppnJgRWuZNGIt/Ddr4
3zhuK8e8ns9GDGNJ0phOnqXf7HCbcuSCgHoUkHu0L9mjA/BuviBtGwDP3FeL
HetzZDJIeylfquTqN11UDk50sKww1awV+E455sOmxnX5ltPL+nIjZnJW8XwV
QIJv83bjQOVFXiCmnSEYpIYPvmuWJka0hb3aGONHceS+KB4X9IGQFPp3P2bc
Jprp9PczUWvv46fX+VT6hfVLSC/enxfGzalvNhMytVIoTAHpYSag6GJH5pcz
hRw6qIbQBgqJriFt2urP+UYsADdffgYycmd5EYySrftMyxrvgds61DcA0I4k
pPFuBTF1CzKX8H3TCTB21QRmq4t2D66MZW4UEPS9xcPtV+C0ETIta+Q3MHyt
0LiIkIBuf388grMKxCxMs8j2ElBd2ReYpcaecCH/3aknc+zDg5qcqu9Hurtv
LiuiZ4S/TVC+KG4wxN5pGZnkKOT7U07Hc0D7EGX9Z4S3oXFwYDafABDXhJuD
QtEa7KfHQigrVxwwKpLxhUDtBpItGHy2Z4LFlIOUnOXTMkyimOEggBW7GAf5
gxrn6cuBFWQAKW6VtG93G+Kt8nu5YyS/l90bZB0dd8dlJ2giCBXeaRvY40Ew
qj+X1CSeHdFTvQMqDT3WhakdS8y+O3FiuNjKreuzHKPcsdH/JefJLten9y6S
G9qnDpcffcW+fygHs7qua5Bl1Xpj3cyG5yHHkDf3v40QyanofVj12XFuiAwN
kCx2C7yrcIkxWGsCGztfFKuYXUme1DahXSyN4G1gjymiYaX39yNWLn1/Ufp2
pQYBfBTpH2L25MAhYXWUNwrXjJCvACOPFhHLRvgDXFjaaKL7gS2l/q6HKpAa
K24+ab98tRjBkLwhatR+ruIT5ztKMemoO5s6nTipk3MmveoFsYaUbKmH+fRp
8tICaK36zL7aoQeAaFyGeLB0LyOZmEf/9IFsa2Z1TtPAY/W/wDyII4or8wnT
oXSLZLGM5bjXahYLWkYnmAdtLiD7tVIios0emx+nqTyVSNsDQGj1sPTOuRF9
RMPVOW6kM9eQPjIE2WTYOTSxF+r/SI2Myhx3ODu01CUoTQpPFvd2vKQkmAEP
VzgIxx7Te+rdMIPWKV0QQULtQUlkruzCJ1PNwOaNiveNgk3npUmSWMpwmcLt
0sOnOexffD0TZ6qAWmlm3SoWRIER7Jl4rXLB/QArfW3egNJ+Ef6xvh2hV5GH
K0Ls3FotLFDzHI36/p2qTMkOpTA3k2wf2mikEBPaPQ1V4Cx9Yqu798q1B8Tj
tBpI6TzY/xII0Cbpv/LkorxTxjteZrD/eXsfzb22e6sChO1sCwCj2zVVBGCt
vyuqEV9IWgJjOmAsxixXyM5nekWHey/8LQ0NrlDll3GRRHp4MsjD1Wr6Fe25
HgUw+5bpR1xXrh/CrnsnNcsYt2MKJESX1Xa24fjobx3EycbC3MfY1Vn8H8ng
/8Ozgb6SYhlgvTwUTfnpF2CBARHhSen20D+2T18pQvnErMNbUXG5IQwm/BjZ
eSrvP89BPhLSvg4bZGYQh2s23K0a/3mswrway/foXaymtUG4vVFNy0AGDR3X
+2RDjjKFK6lmtXzscdhW3VKGxDXVvL0354JfA+SufqTxvAsJnpwYjXRAB8i7
9fCejI5sFswtD9GVXvACKxiRCu7EAC7o2gCCyoD4JsSoIB1P/r/vdjDflgyC
NYIwbngha2APdrkHNY7WW7xQPauhcCF90IiokmrnvfR7BdHwT1qAvBFcNtXH
jw1PWlZo2V0C/zW0jYrqvqWesWP3Nnl/mXa2/LCgDg8yQV4CQu1AlE0wXbfB
NkXLA3Knue0GmbTI9OS2lOM21glm4Z8lOmMxnZZxqZMH9RohnhjCcfwKdLCE
WW6DxHNPEbsRaGZcZXWmt0N02FMQ26vnAA+s1/qlcUyiIJSrDs4NDHbZctp0
gw0EJxK+ryE3dX/noo830hiP4krSmt59Dj5TWeVKizYOKBo5UahObn5Y+r9i
HsQJOi+SqtGYa0zfannvsYQPjmUJbYUS95z4Nob1iRSBI/JfhC6QpuVfV6gt
e/2v74dKHGPoTHX9H2wzNnyrd3J2VmolI5Bt1lb8+nf0G53s4P079stzv8Cm
JTYqaTsx9atalqnfiqiEfVjBFbevr5Uo0gpS4fWTqP5rUfA2ot1Pm4fj/3Z8
SvG6JO+A75Pe6KKm+tKrUWL5B48NOgPKOAg0QY6dULD58zObBeop5KzR9yK4
m7crt0zhNIWhA8ASBmtr446B9yO2iWUFkloc2TxMT01SKZK39eDvdZuvV23E
HE874MTXyz9P7FCX+Ui9BbDF5ipNe1CsI5Li2DvdgQ+20p4BrtD7cKtzNTz7
5w8rXs+DHtyDaACKZytSLRO+V6bEy10z5/avh9OKWCFPINh+qAIJTCRJZ3UT
44nSHZFvOvvqGEC2jh9YqHA45Oj+uvlzrc5jAJr4h5smPhA/oPeNMELTxaM3
5usR1jVmbBavKmwTMFi5ZLd8LBZ1CanQ43FOoWxEST/Hbpvg155iAuifYPcO
uMXHDEqcRphgXobwTcc+vDCvrMMQouEEqUmXXh5Y94dKCgypBCQtrDokKsVu
YJ1SPbI/bHLTYGXJtVm26NvpzV4ZTIpM2RkURriUCv7Vx+Go27CcLV34bFGS
upys8+NdkhDIDrJ9xBzJi3yz7xjhtxnN/GWBIQPkEWpLcDnqH02Ors/JC5Mn
ObZPsesbxZM1P9XYvqJWDLqBIRQmZn6Qh2xlWDvhNIGPL1wKUHIWscKcq1qC
PiNzUJHIBTa6LoWucmqLD1V4tjwvgPEUMt/nIiIS4RSBt4begMnhJRyxAfyk
lchBbbU0+WAa9tXsEgm/6WsvFCoTnLEMlTELzxhEq8NtO+bAbutq69tiVXkN
vysjYtFXpqazbUrwULWcJqIVpJFikaltOC/YNi8sC+yhlYQhg77htwr5nMul
7ZnE8INOwpJPvd370SdX71RRIwDOqHhXMSQxrSq3qMtn0SOSDfCJQtX41PSZ
fhRIQfehzjOdBmso7vWJ97JRIulLidD2G6v9fHlpAqBVWtVXiZ/QNX4ozNVd
WyeBXSCcSfIqzllinsqt/GyCdU9vMphDlNhL+xON8ILKOqQ99GKYAkb+xPvz
5mrk2vWXI+XA4dYv1U+u6GrNWXo0SgpV9II/OJTCzFsFUoTnsUDRswySCoxe
Cd1d6cC4cmT0d11ToeUsYO9c6C22A8lwpyer/rGMa9gH5+vmr4IWlMRdy8Ya
U5smC6lN/15h5F+HUFx/70YXmw2vlbdBUYZpxAJqyXW3ki2x4LYze+7F7qHC
Vh9HUwgzJ0dTE+4TcChoW2YaROcTe4FEeJFi5Pvk6qUI/hA4QpBaCz9x0mql
P1t+pxbags5BceEX75+fTLpwuSnoT02XuuVFVfNHhe7ixFPJngOsnUZRNzWC
RlgeSbEz+tm4Kl2RtzxNwJZCyb5pitgkbEY2tQ6qx4WSxCA2PwP8GWvjhB9X
31u+PPn5h7T7yRk7881JS6D/P5O5BrHBL86VZ+A8c8rIwYfvK77OS1SDGJn5
UE7q3WL6fGbRU8fcwcQ72h2kvfctlZ8SjpF+DrIRcOFqnulUKd51TLy7kzgp
a9uVyoE2QgxezZ+GyojFpsBuIRnRn2pQzrB6blIBNujPLB3wUxrS1yeL/eRE
3b44UVUVSaysz/PB39S1Cz27zldszbuEg7SkbMQ1hoOHAmXlYjd2T+2QuuT/
sR7x/6bWYKV+xV28iXEP9w1cmeYX6aWjXEYDAnqw3gg7EacClLpMmD4qyv+U
pvMjE/E8/KkkW3PAhZvVFcfHnHpTAX1Ey/YeZf1DTpTNovajCR/rlPS32Csj
g6+zNHLAY9U+U1w/rae+0LqO/6Ad10RMvW9A7/ZMNKaAVMzRTBQO7C9rS2lA
fAi8kNgILVsXWhh4juSeboiyVEyJRzXNanQokpmSaqQ44VSrcq3u73q77NqV
BmQ209+Th53mU2hyFvcQr1ls6jOYMUhhn37liT++f9xajinA+aB0OqFWxAQ9
wAJxIRNNGm2sqb4HCcQh2I6LxJGOZEzwmhFDVXLGcc2gBuHFIR6Mh/pzpBoP
zP1a+VwjrPSxZPZ07nGwoXescMnHO2TsT+7pxgsX53SquR48tCxXBPrEPFU8
TGyaaatO7ALFQ9JvHCbnMjUxCkJuLBl38Hze1fUtHGl+IRwOOXSL61xaYoOC
uOXl6PJrX9RPPlKK76zrvx75ebcnGXxLvTaUX58i29sMMY4KeUrd3Z0BHgiL
krcBbz6OL+SZn7cobjSPS7O0e/qcoh79ZsjICh7y0vEDjhcU1+7vmXwruf5K
j19VwDdlF5VzFV+vTR+cOZ/bUJDCqoDiEPQDl2QcZ4lsJNFFeUr43zOekwJ/
fKYXyNJ9lEuDjD1A3Yp1l7SFdO/fXTGNSX3llSxE40OcvMq17GFTf/6E1WR+
dwTRRGwnxyfvoXCqykjWDSq335hKSfsB641Eua9qH7THGGuU3sMMOY37XD2d
HAbtkhUrwnYC4RRzsIQK7ryQNl8FTWk8FhsjLOp7KgAkOAh+mZS+6kJ8WEW8
erAdG8YkmHAsrz5kgGRWrw7TKsg4MDZPh9MqKBl6z/a/17qmE3OJeZLSPZjh
QoxTJpxiDMsBzHhADrGp7BMY3Lkvi7u9TUd0d9htF+AQBPoCw9PLKxTdd7Cv
9YtQSMSLu7mEbMdI6aaHbdmOvSNnFCOFJFLjJEMNns+o0mCSAI6P6s289ZdX
tiq6WOlP5h92LrDfXpKfrLFimnm5TnN9Kioy/B3FL06CozzydOQnFpSNqObI
CCLfzSkh7VZVn9DKtGiuQO+tVMg2yyx/dodzkfWJFR/SOyxyMk4nGlQRR9xZ
Cn72HsoOwltlcmaQC8+2Ik+EHrNtwFIn2GXqAF9/GmsK7xLht4jchQt2iPuc
GmvfUrSFya9j7caREE0X/6pFCXbeUYKTAQCuF372O89e03PbKS4Oga8UcIho
0kBKAzgGo9x7ZG4IkQxIFZTUBbsrKCvkzkh/W/V1+Tia6pM8DaR0G5KIIASQ
9RL+9mExp4LWjKEzI44T5OENQ43d6EG7FjAcUzSHDAaAhagldyyvpqaEbjVG
QIoBrysSb9RDMgr+WOmFDO7cxo+Jlk0IJRAVi+w8Tt+bXY/gE1MVA0R0vEJN
/gIa0vGA3YxqkG3HyAJzI9Y9e08DGk5nHr+NB/8eRlP3daY+CSiG+WgDMtoa
uok3gRaoynY3PNPB00GG001imW3/zS8osGdmRVCmHI12Oc+/EOS6Cyt0o1e0
FOKJgz4W/rWvyNa2OIsSAS9EXshXaO8rvfNBn2XbQ2K24mxq5emC5MRZmwhH
kCnzKYcKw3VIvB8lfCCPDZhlMCNArnELljgEy5B391byk/1Zxrcz9gESLjZd
3fFXJldd0OOIJfvjoi2sKAdGh4sTpxjGa+L7A09PshE9tTeB+OVnEFdYm3un
SXXuKiSJdB+GVXSYX1CxV+nluxP4i7akAK135eEP+hM5qz1n79R01b4i78r8
Sq35JR4SoE0TWsN2Tjqnfm8hJNgb35KhlciqS/hVd2OrBNAcC6OsdfznU9/D
TdXc4iC6hL1xtNn8Qws1DTOp076LziQOfBUr6YLUKtj3UyqQTpMinAnnXBJH
8oudy6i5l+YttosPJ1CwTiTSjArdU258100z1nRF+uc29GQ4CpME3ZFGgBh+
Ph6stpLXmRnEvs3fZ8JoZmNYsrkuYoocVrxAzLOOTKjLN0r/TyjBjAq2mgri
cSTue5Pmor+zoTLO7jZl4huEcP5mgzVSZKhQZ3ZcbBjo0ZukYV7ij+0t2HDk
OpBUVQhroFI6LHYx0fOuoapAXA17XOhKBqNed1WKi3N/ju4NR6H3iXgHcrsw
ba8hucpR+9aOaTiX0C/oOxiW9lAYcs0rnqOSlhm+b6ooaGlRuXKzFQSOClfz
c0/q40a4QGmeC/vDB0MgocuiAqmCSUdVA55PIal466RVcgMcQ89m/VAv8MS6
3w8yD5FfCBr1slzmvSDkeZpGti+Dg62sj2YnOUz4uXZNUB028KyD8baGByT+
P4z6uWyw2d0BUWz0fWMxD6+4/Q5P8JewoJ453sB56g/GupsEZtueqSJPIE1j
a1BWnVK8byWYsHHRY+G0Khxo4Gz1pPeaoxsG5i2+dj/BFNGaPmebHwjtbLfn
6u+9cvMGguCezjc/ndS42BU4MX+dGI+tGDeMJBYWOWUyBu/avx4Pxfzse9g5
aOERY65ss/Wwa09Lwn6AqaJn7BCTuwq7vGKUNyCeYcJxWzVBW/TPsqn+30rq
ONHXLeBCbaj138rv2id4rCF6xD2N9+Ik8WLowour2gNSXBs4oaVDn8IhOEO6
+zaKxOM/0WmI9Lhb+BlCc00dK+W4sGz3s8zCAy8CLhXIR0m+cYrzpFdzSQJl
0EuJE5n/iY5lbC51KzuDKqSu/qMg4EItuZuLGEsukzV07a+i5+84+cKF5TzI
h4IWExasGM8y8ZTZHe1ovvPZeq/8qPF4M67lx8D6SBD/7qnbYdQPLC7jWHOQ
Yowo1TxJy10xTdFHElQy/9LnvKqtAnuiD+CJ0uabOJsozxvZYHcMw988Z0O/
bKDlR/ruK6XxlIHP/KiigBMYB/4l3PcSbeSslWcf3Zm2z2n+moCR3E0gR6eG
SqlARYrkvJrR06r5H/cmi6XIlDsyceEGUTJKre/J0pfo5GlWV3fKS4GkTco2
MRoT2N/0i6uvgZpOiwxTJl34UrySojsj+dDd4XKe5iy5pDk1vTVursq5kpaa
BZ/yq9CbYb1evi8MQLclX8SJlV5wMqj8UbR0T2Pmv/jtZo88z6ix068u1ayI
gt4CqsJeQWI+oc9lbsgnuMizaj/p+YYvfjXof8ljUeC7r8AZmeeHRDX4zp0Z
FvRiIpvyNFqS/MFxH0QzHq0RweWyOVou6owR/O1OneKjVLVYfixITsOJiYgD
s2jy73SMcEGempdOIHFyTXi7B2YtAzVkRXjl2WBTG3U8X4z/SzIZFzgPtljl
tv77vjGQ2/PbPoF8YJy5ebVWduF5bd4dJQxMcgTgou8tF8oRDS6nkuv+9AMw
hIS970IJpRr6wliNdmJ7nTzywSP30ge4JxpTXqJbm+SWZ8XWWoTNbKqYCC9L
/F9mA9I9ltBHbqmVApAFoesONEEXHr8bk2vQtyIaLmTtuC2KG1rcIV5p1Kek
d3/DLr1hm69mSQUXrzqNf4PPz9FvaqWONg3ub4qyQUZAsdXIjBjhgI2YfGUT
zvG1J+XcW4/Q9zsVZwQOj1t5SP2vHC5Z37PwzqvV7yWhvF2CeQoXRYwOyPRM
FfAJn7L19WtkYLLXjnxYPMa7G3sUTWy7VV9KymzNYO6/y/1Q3fOvy0f1UW3J
HMmqZbg/GN8DBnU8sPGNkD+r6iUAEbkkv4Ts4IX2mqbi02asX6cp8SLF5oiQ
jmAeGH2LPnYTnfgQ1Y2HfYzZ3DjVwf5+OaXD7opkVi3y9Xa08QBr4+AmjZZs
GKxoMm63kIH8DI2NwRCCI+JnNKV9PWdFjoliY9MJnNwsI9RKzN/MDUcphGEs
ahetqf/soiERMZNE3XByoCuO+CPmXOpgsTN99aMkkDdaYXVTwVwZ2vkWbx67
XQKYibe1VyDrmmj0GAoc4kfnmoCAmHqUM+Rs3pXGeDQlUHLsr3jBt8TClHbq
G8zW1edmNlv4J8s6fz31+67qeVHvy/hgzzUfF3fRPRQz8Ugfa2sISiO/tvck
HFnXRpkMRezzU/TULTMzQzQCBCFFf6oTE6qplP7ZREpY6re8KnwaCU0/plxH
iHiul+PEUgaGJWkageQhqkD8DKDGXwcSOmOF1zasRsAZTV6KCIDPtCy/+/Ky
2EdjMt/LyXG9UenQR9+jqrIEdSsyMU6sQXW7/wdlxnwBc1Dk82EubraKmByi
6wDlLXr6gROwdC3GfKtGG8NjWydqfk4quwwM1lTzJ4c0+EPU0PXTDScafDyQ
sDKNLlsl7xMXbF+Zm7yVlhd4G7U1mcyFjqT/thwg00nUmA8qHcNH1WHsV7b/
Sf2t1GROpM4aeLBtnYK3zeNftXoeU1owtcz5F2UNEN3KZy0IV7suWTI3TPWY
dUafEs8FTffxE3DDFM3VpZK01LAcHyUa0q3qTpfUT96tsXxA6FGdItgMpO0u
LEpuofgFac2lh9VbDLI5xNnvqYosPi/HsQ4S0hYwPd8WVwiuWIVxzrP6V/kG
TwKNrYZ0dTBSgF0PIjhWlB7rNVgQsgncvtSFxRE0uv+Zaf6tzb29yBJk84yX
MEl7edC6OefBT9urXcXxpeJK40Tm6dqFxX7JHAXnlkZ9/ECpTdcsQCNpZVhK
jkjkxjOsqSmOhOEI4EhnMQU5UUUrJpus6RwXStgWpjxiw9usfZnEgobmccQR
YHSxfifaeNGSoYvi+722fDBG43hHl9WQ1tARPBJj+XKyZLcglKd8HaFldGwD
N5QafyDhmSz0JbS7dJqNA6Ne5CWEfl/F81V1Z/ycT2vlPwpk4jno1SvRnqKt
Rp5JXM0g/2iMlpoV/dFq3WWSH3ZjDyZmG++AzJQqBKCGjKTmgvQOgk/s92lE
n7XCXDRE/q5JrtprwzunOcNXQyuj5bB57WUKU+O+9maLGky68Vza84nv6z1f
RZKKIeuJ/9gnzzpHpq84zoxSWEkEH+0bYbtJhiDv3DwAKgdDDlH/l+ueq70e
Z5uVms3f4nPQU+iBZzaMnEUs7Cv/Qm/xYaMiiMkB+TJ+B/WZumE+on6subLr
K85x3XA+XnlnDQGXzzQIqLVluCBQ10g/IIgPSYqTGAh2jNz8Y1IhnW/otvQS
1daM35zVAISeBONeLrUporykfGCsm4y8beFA1NaJpXP9a3/GQVLb1TlsEhuJ
RcfR8kPD9UY3KYpLJZv+KL7gIS7wGsDzsDUAAfjDBmeXfnQGT2NRQ2y7ZKF1
3bBF5WnTlNtRm9ni8OE2Sa3wLSZCuEX8qlpL4qspwhQYiyEWjurfx1Ha/1HP
2lLDg2DHVpzbOXp/Lgl+ozaYFfyLgF+0efoBrdXXugWDfASAcf/Xhis6XxRU
iCBFLvoPVIkj9OElukHb+S+Li4nZ3b7546Ual5MDhSEDxBehwFXkPLXQidOq
BFJIaePkbF37LPYSPIx7F2kzEi+33ducOm2gvG1YixKldH2wIXIKg9hYV2Wp
FEoYNiJdKB/MDaJ3CMqz2svL8fDqIrmFReMi2sLAQmAYOE1U6/LolQAxWEVo
hAmfED8gX/6+er3wH12Ux98WdI10FEk63sHzO1Jv91AuiwH3HdcYwPVqdk42
LoMOsgM/Ncmedk8h/4pssKBHidHRvu6Z6BGzvpwCQfjb5e+lCMot4ldFLbkE
UVJlLtQ7Ty2eSPaaEVADkweLhyxuX+t7bzIQuwC9NpP6W4XMgiZDy02Y/ynq
xn9OsOOPuqLMKkNG5rZWC9NlmOCo3379jCGVcfpmxej5SrCGHJLferVTRorO
+9c/vOZiKxZx+tu7M9sV5TDcMVf4GHD1y/whvkfxSlssD2Ijf29HBDsXmTBT
kzPb5M+oLXhKZnbVbGoa6EnuPbWEv0zcvf56zpq9GgcgxGwT33lvKB+C/SVu
5DIEEEGdmaQjVr6e13inxHKKRYzt5ud2V4fvBRz4wY4JxQa4eYp/z1ROexw+
iE0csXq1VuWD5Wn3hk+U046WmldJ52xWvBGcVTtggo5MgB5nJlyQG0E5CNrx
DWyCfBs5YmyEO5XW+3jh6Yj5ujtdVj40WUO1Xq1kDTdVGTWT6NpiIu21mjrr
jPziWQQNVHa+G21JBI2IL3DjSXknZXYB+UxkFqmxkou4v6T0e5H3upsI3mAs
k5eIhUuGipFQG+uXtnvUjigi01aUipgvfPKpjFyQCrhM5sNaMvdSduqKAWWB
FnMn8CRYVCiQ/vXeYiv/QWx7tW21z12ZdX/xbwzRAvFMW1rNp8CzN+wn3qKc
tkGXvdfyXZi+cBesfq0KPEmf6fxV7fr79cD1eChYILmQFXR+BgH4sC1hR1VE
TbmS9Ks7qH9Pq9fdXGLAAq0jHGSNYv97gbTdOlix8AdBlPZw8GWB76SPmDSF
IQx1gYTtvobn0h+yrBSzkMHf2BGQfPR8G7DWLpahIU6/iZFZlNuZtXDJoy0s
A00S05LbS3Hayn7QyAm1lWMC8ADVwjv+UouyqB3mq6U9DmnzleIDuJDUaQIm
1MBYw3nJB6+u058jqTo1j1yG/5YSZSY+MFNyDM/JuZgelxImfZwyikeyqhiG
jLEg6dhypVFyZksXChVlcjuYR4K8CGVscTdzzNNDz9c+1TZz+S3KFbiOZA5c
OkPHizw9vQP/MsB6m4o9yVdEaKKY0g4bUvq3JIVDOMd6dghnXanNg/gi/Pqb
klOmDiC0qeU16hcM4PLtro7e/CZRoUEyHlw1tOb5BzGeHskYKOQVewjRLQLV
O45Y+EfhwObWEUEiGJbewHwJLiJPINeVh0N6bi+/WomMycbnZ4k3EUQ6sAMZ
+ux0RZUUaLu+TCe2ViEZJmRCdh2uZkE5YANPTDcEJrNLVWxmX40O6X27jtFM
S+pM4iPpONa+IND+00X0YU2tkEpwEwMVnLy62lbgkvTuRufgjxONki3EAn8V
Md4Z56Usf+mFatb5tFyxoxmxPLuPOnd2lBT3SM6vwNMmz1AzPMXAz803b/MA
5S0Cu/BcShMNNAaVTznZyLuluh5uDl+NFVQTnFbJV7Kqa17lGWntq+Ruw+rB
K9Ph1/6Vhc+ClfG41H//NffH+pQ/jmqUsI7/QOB6owmLKVgc+TP6HXzyMtqf
1JtB47xPs+/+mjqIWyDYZcO5mVjDh+6cLAwaByE3BbMIaz/mXgp+Mawg04q0
O0VFD1qJcj8Ybxs5TpJw2iweUpT+ZY9lltqMYdA7VaW9kbzFmM259nJOC0Ur
5cLCOoCiV5YROOxYW0194wUpLN+Og173KdxRl9Z2l4UtaoNQpoFbc2jbHTP6
8Y6bxw6p/G+qv7ka8Jm7abSZ24swXwS4vpQiAtILIAwJGs4GCpNtvXuQOyRb
G7byWQ+gIQPQmWgChq6Ont8KevvnIAkfSIgyxMekpkFzGSF4wWUiW/jR8U8a
2NBrDC8ZRriCbNYOhsj0ECJgtDoas6fqwW/PSt7OjmBuWMr1Gc7PA4HQTF6z
rFiHa2QPI2eN2TaV19CJ+ugPrV5FWgVYruvPa258RrzXib7rQ5sGINXD/6yK
LidFl45TCmi5r7YaQvl77/YNZzSBsacYe/3AWHvf/w6qWHunEfQ0YsIUsZhq
+b6vwRVhTJl+wIVDazu/ueTkU+eiE+VK+Q8oM3r8T+kh0TDeONwBJLCDAj6Z
1TMq1N4YigKgot3nENeba6VUALW10mv3euOxHKTJ+PB4+4LJTphHsXPeQCEz
of1VskZEt/afXBb9j1mqR2d6AcBGFdPuoUZv60bJI75uEJj1Ul+qbx2bIa7V
OyOT4GANMuJ927vx75jQjIzjMljgxsFOEoWy7OVM+khXFy71QG7DOchZEg2l
DRkPrjTGpsEDoBvq+cYpYjUA0mrr0BmsKmOH0SM+E4BCPr/A3qG0/fP1MbZF
6ShMjFrPK+z/mh9zZJlvjkpeuw9BZdA5ir3Yf5uET8akSNKnDkAqBPHGnG5R
rxAyfwJlmtMMwAtc0228csJYYN5O06xjs1RrjDrFlzHCnhSeljm4SQwItMaz
lYdzi6p9Wvcw25wgaOJbtXrJrHqUAY4OuW/f9W6dyyn1FMbB2emvuNlbbE2v
8fntOcOUWqsksj2eMEihcD3nZIK9d3M261ckx9/8f8yT1wBMWFUxxD2IXPo/
y8mURh+5sRERSiuke8aeoMV18AeUfTq68DkYFgB8RbAj3891/yzlSfrl6bJy
ixMHBgmELMdMnGEyW0SIt+2sQAEdQFvEpgNpHYYnYeyzaWBKHY7JMqsXe1DL
qB0M5huSiMikxkf6B8JMVG57EKV+DaT0pfxZYes0MtQzXTjm3zgE+AOiAiRh
A4bKtqcsS6HzgVx0NVb/0TsHH71s6t7fCR/wc9c263+Q/xgeYFl4I9zl0JtB
SB3R+5pYFRdkxzBVEIhAo8m0WoL95QrFiX3mcLyhIfjYnflYLBjJQd4E5LM3
jhXLfAfXFrJ0dnuE3Mk02e64YhH+aYtQNXyFLui8rKOGZvnEHuyMXWpL4Tmo
414svsQrpiw9ByUdkPnPLUQnQx01kNubUlJxUNEhTvB3LX3gYpNl/JApIw9j
GUHPoPluzDCoBc1Bi8ZI9bv9T6Hw7XWIxCS6fR7pU3CyEi5QlNY1XC84B4wc
BL3Oy2+hW1JZYQf2MnC3h2D1PaPGPBnrNh8xr3CH3FCQ9Uw/EieXA71JZtMP
gTSlPKdzkei5rilq9frfA5XGkWEtUD7AXLpZQT05BiGzJFdTpg5WC6Y3qKw9
O//iyw0t3v8tarTNyy6IleEP610vuEh4JcPzJ/9aSrRQ9fxGrXyDMZntVnh1
qdqtCf/ZPEhwnwA4wvMl81lR4UpYjB9oUJrOVzgzSKL0Nm3mQSBOORR3zyn5
dugwYJDjN0uQYzZA4tIP/N80tHjvSgUyGR9wy04JErhrtfJ78NGreWeh9JLG
ewZGoyE43ND07KfVMKzSNX3KBGDZJ1Qorl5mtP0t+A8KvJpcEnGsNT/DWuUq
+nXF5I2RceqSQQURCBngICkgBe/GmlDYXdFR81brduA0ePn92UkwBJcRzBCg
iacyCDwBaACLHkplJDHscQPLZkj11b37m6XMN7KfwrmrQSKs6f9kM5tGjw87
7Sc+eeAo0P9dzEYgnf48wQpffIlPref8GXztf6IYqCGONQR/REzWaN86dJQE
DgH/1KKOrhMQhLJ4r6/UKCbWBqvy9k0BcTd9peclAJLc6S+z+UC1/NNO3G4E
iH1UtaPCIWpWZopTWSdXzvz89RHPJdEhfU8CiUzuDw7QoTu1gHJVa2u6UFl0
2S7bjcdqKk/tw2GaUTlSbWwNsfx0irgQOEVBoRQNO9NAnEQ0TcgDyiCPlkqW
OqjycrCidtFzHIAj9wObmqI9HyFnZIgmJzLeml4CIqNOyi7M9tuhobnC7p+L
+VPSsztTBfN/ts5NTocK+zi8ZPPQJlMknflx2WIJweXBbcnRvCPBU0tzjtDC
VI0dgBqrBI1BANkm9eVrhzcud2+G8GovJNcHY3hUDSxX1zRQzEaU1jkMXysl
cU643Ww4u+XYm/8B1ntRhc5cOiYs2XokiNwxdSqXe8dIBtscs46EYZdUrz8+
ztcmgSJdUD+S6pcbTB6W5TzDZIgZUYXpC+BGnsdP8O1WFCiBAVY+NKXgBGZy
GlHXL32XstM3QPF1FqAuXblaGxxjE3h3AN2wrQ1FeNjpKhmm6khD3Ashw+G9
dyfbCXQrsHdjeFLjpkLiySDq0l8R7kIoehEp43eETF3ZN2R89ZfK+MU/OJTb
dfoWZ5VdTkvlYY5F67zrr2pWRzsX1gYO2BuVNaZ7J65K8jsO+wQELJ0lzEQz
xonKRLDvgQ5RAjnzn8pR1aj1aEX6+WPd6RpjOXnVwSzSiRiRMHN3sVDbbiPi
knl5ZA+EUIYT59ulC1/M+F4r18Xk69n8arNLiG9VIJGFtFT7f1H058G/PztV
sm7Ac207JXp3JxdX8SlsWWUnkjeUcnmrWUY6GPdJOfSS7yIzcssEDniTNO90
cNvIinMu3vbAR5nUwreccBlZ/uQx6QrFlRGcRWPFCPK7nWreFV9xyA+V62Bz
UFfjBeYXlE78yDvLe9FL4FH46A7eK5FBz4tm36sSPHmMjGKLmKi15GbhHSYv
gtkR5nsrOdLJh3nBq46TE16yz8ja0OxrXFDSNAF+dV6ugaeulWxzczqfKcOi
IPBlt2MwPIGHuJhRgcvfZR5K/6CEnFHBZB3+SkBj0AfAcPFXUrDf6LIIlcxE
RsruY7YsebRr4LzSENzcFEFXsbIW0IIaaF2ECWi21sMdmSKXRgnoUO3KSeKR
s8WDhZVvALxBnDR9xnBIf7QObFThTcKXYtiMmuCfky5fLvFHlyg4DTH7Hv0z
Xk4MemjD4T2EEto8vskgAv3M4eZLrvssqvgfiXE8Y0RdGS8+0oeJ1Q2+lXpL
iOii320O4r98bwZujFZfau2Z6o+eqWinfPh+BB8SexB+t6gyM9VM4BmsSnFF
y6583ZvRwF15c/oq/9aJfBgIR1+I4V1+In2Vnyr/jQJqD1Ew+3kZ41HSCtC5
i5w6ESnHdvMfDk3k3GdVRZ6JNdOU0Tx27fIyhwfaIO/Bm16w/1jWvADs7Nyh
SHN6HCWApdUfxNOGJmwqhqVs2SXnnJdgojHa+ApK2H1GJi7u2nGQ28dc+3Sw
7zHVwY7sjZqOZkAvP7jVL0CMaFSKZoqh00VSsGzO5uU585W8mT2bFfM6uKci
WTCbOY1JARE8VDy+GYdgHwnJZHPls85myREqviG9dB1FaL/VpkiGbDoC1CrC
Omfnea4IUWSZHYsnFhiwujJV6VO/KYHMeTvdSCNLDgbk/iE0CMok4xCufFOL
mZObCxih6P7DQW0FR8t/r54qx2gpu9MDtkhWfSCHFgcPXCDIA0OokZbpt6o5
3Lw53TW4268lMRmZDeMkM6Bfoc3ohfC4uFH0IXpG0aqMZkZCwNTZmFkJTt9K
iC8dnh1PpLvUlLkcjHZLo5HJvVwXXYxHiT65RKqdPmbCnGRbGpSe2U8c5VbB
O5Z6BlbaG30eiFJpTeQDxqxrzV3vL2Xt4KsrufOdA2yL6uJvi6eVOnqviWTr
XcN1x5VURgZHEn2G0POTNYwhivF7ZFVhizThVP0EURGUtwAB6otwtF4Hy4MF
BKW22WKymbDbMymScuNVFHmSC1QKohyh4siCJpEH/pYuNGXWEhcP7p4AdQwL
z3AtHhUAnZ21Gz3WVWXdQP7FaIFEE9cBz26fGM38O5KVirURWPyEOMFwstvG
FWb5C3spp5v5NIUzvv4sxXLSosnq5lYXCyd6atRqPSN07edeAjrlLA779TWd
SZXoc9nby8NgRP8LeWQGqKq9DV2SVifFSnFKjtcdBwIRcpofBAICt0DmtV0g
Ab7uHj6BWiPdAcnIDppjTZQN/1XjHFFAAuYKtkBP8Axa+lrHGZXkiONsTVeY
9Ev5/KPyU6ngdhX7i8WWQsIZbMWDQMaw8aARE+Q9Nz/4Wz+XkBPYPe5OIItH
A8vW9vKF1w5FkL19qQ1GxwtwgTrLZWV4UhUGB2nlxzHfy3r97G4zffQEVX5M
7EoeBD8ne8thpeYGIIP2QP3EE9PZHoagD2VWZjvja/P1wf+t4MBGjDGWWO1D
c9j1Hn8w3LwIGBRJrMsMxMIgevMqKQTYGYy/IwXPiFAx7EEjId+N9P+bPYur
1o33s1gvvwjR8687az8oST9/M91xUlDMic/+vv3NlVEqJJg1RGBPxHbypLQp
7ma0oKoSS8DhlffIQMilS3yizQ2ek349Or9190xblt15kni2QfgRui6a5QIU
jS295+Byw4awR/+6KGMgFYzkH9adCQr6v5ts2nSJk2RRSpivfCXqkiRTN9Fw
SpI63bgS1CvMbLvR9+b+Q0d7KWrmXoh04vYQ1TfO5wKFYOO7YpgZvd1ugaBI
qki4gF7KIxp+Y7qqLCv6ibgdLEYkdQCuXVr6JC9Tx8aqqMlcVmi0Tp6X0WfH
3W2vOTAJbpNyu6ThtUmFDHIrxwwEcPBryB/kuHw/OvXFzP/fJuDOK54AUHUH
MNOCipCW4cZMmo0P7+BsbJTJW4x2QE0Y3MqPD7GKoQ7KAb2BL/muOgcMSLut
wS+4VGCG38wz+yJHElSwPLw4oZVc1fMG9FsrOOEzfsYbgbyM8t89jJlcrh4s
x2Tf7rMY4Ghd2LNWZsuaGb+1HMaxniZ9v1Ux2ErQfDFl+dXbqhIogOXaEttY
8MWX3bsJ23Bad0WrROykrN4JaMOnKp1YJIe00mjPGo3m5uxUVRGKq2UDgGWQ
uDmqZJovxi/unQDBFOY08bojQcOTqvSh7VFiGeDmCN1nGQUGI2QkYpzWmffP
MdVILc3RFQzTWVWdfx0zRK1i5X1IcdXqdnEyJq3LI1kbhsChWX925VmvBZA4
hPbxDTp71jvmQQdQaEX4CzFErzIRm8Ph54MKR8EjLb3o4vzfp/2cm1axr4GI
uih8ZzHBbyEHGx9oHsWHQFF/+F93libDxENLrFGLLX3eze5hszJz4Wrqg7/A
iplmiJip5Xnrn+TysQ3hzMZ32gDScIobB7+25JcIgDJDAc686dqj3hoMDxrf
wZVYG3jDRa4UgkEV2xQDSc4C0LSNPc94shFkNh1XKykIuiyToGLTGQmV/14c
/EAHwgO6ytPBKQ5GildLT5GpREOkobUXb2CLm8PMmCo40tA/iGwYWgwsHXSr
zIv712XjyfkySrDtJc10/hOkREZzF4pjYJqEAOhpTy/cZeOsocEoMjaOb+mb
QAuJZuCKAXjV147/OW2Gq0XGCZ3DsZgqmd2zxlBHBFs2Hy1byYQrF1uQ3aij
akmGdg4347uDjBpwpqF/1989VMI4syvx8Fnpr4ccXtyBdpAyMDJzbTIA2tH2
qA0QS+JSYiP5jKnzMfv7Dm3k1isumsoQGPXzyUoz5z1D70ci/tns8+8/JU5U
c5bhBCYTcOfGlsrX3ZwXao/4sR9yAiNsK69DWGfT2luyQKapSW9DJu21f/Lw
EJx7Se7EvnRP61m3+9Ksrbp1Uy4YJQVuR4pj9R79VLONS9nNLbswkLKLa2i2
q6AL9Lk0GClzxLGsEoaHVicsZz71iECqhlrAQEzq1VdxhkjJ3+4wjhIr1r6b
KfbQXUQwjUIonzvmeWIlwXFXFUWdi3ByaQMEIfrXfEcrvagLHrfsmM8x3CZ3
uKpAYWMZl6EFrVS3+F26lnIGb+p5VIJb+oGEZgDIHaoaESDhm+ulwiWPcA48
fkOwh/B6ZIUPhUipqLZ9Sdt1kKvB+XQ6vziMw9C1Hu018oHExJEuDCfA8ryv
UH3sKalthRiO4YDVqXk6TlVogLD9tmH1RQOD3DZsfTz1SYd81RM3tu2cig0F
kYh13WU69YK2VFJHECu+LXo50hqpHfmmNT0qzHvfIP+pBzV8J+l+z1ZpkBC5
9VL8tlSgoJAF5ztW8CAvY8VO66l6O4zIo+dvTi2VT03rXg6Hb4X2GhUDZqH7
iywYg1+XEuvEEvSo+5wsrQMTUy7AHP5SyRzBLrk/UpUCr75/X/yH5XQZsFTM
p/Ehe5X59cMX0o+FQGHRAwIoU0rthP1ev7Y6LaQ8qQlsYPW9bWlRiOwzRq5z
baMY1Zin9Fr6uKE6+IxHykuP40AmVNlS149OJLBYGM/FCfH5kgF70k8BEwdM
ZCCGu4zwvtmeNfYxGi/TXZZsOMh75+6tvUXV6PfThQgUkc9D8zPNTkn8FH4V
M00Hn5i3Y3vGaTbOHHqrodc5fvhtYU3qCNJRLgZKcVsRXwdJ2V2M88Fip80k
W3f0ti+E5Z3h30/Hl3j3h61VXejIQYqycZkG9AWQJ1+hwkpWfAwp1gZ6+6No
jfcqSNm6NeqrZ6kj4P6EcCihbx2rs1BlEKL1B4a+3Nbfnw2b5EPcaL7g5fpM
VHGKyxoQDkw508tx00Se8Q4UaT7fr1J//lYvOjybnziXNppg0KSBP5NjAOq7
z7+WgE926oWiQjUFYhUI4qNDYb2/u9r212xNybNKPQhQQgzGTjkSeW0mTxS5
0mPmQlo9VdG0ObwdGcyuUXhaHUqzMaZOnhgm1kIlMwxFl6k78e8FlANDWoVI
VdYrP/HvwoLd0t23BRmiMHpnOwQjZHJDX/sDDysAxPhF1aVO/nUPBemdnxrq
dNnMxG84HiPxCpFulKTPIT8KbC7CKo1u2VCDfVCRpZZLFkp5/pCbvKbyYaTS
jli2nBMgLqjM1uXC55eBpbKT/xQrAES35Qu1GMckI5zmRf1HDKYh2atEf7GV
SYzukVs1kobcCBoChhLjjarWbU+D1lUdigDfJEnUsdIwQXdBQcOeMrsGclJ1
mUB+FrU0fJXsbiRLiR366hxv9Q03sbe4C//ksRn+GyLlTWyUTdfIYILuF7XH
XnSTUcVLi8L/vnpX8GykDyl6Fc2USnoMKMHIOORv051PK/FfI/pEXQvBTYir
A6QEUAdwz01I1h7ulFPyTIkgxQeNTeh5j+aGXn0wTcgRURR3j/l9UWq/jKTQ
VhmV6zqRT9GwbfwyUkJsCyCzw+HcT5Xdc/3BkjgsEWWGdBzahj+0Vv/AUQkz
F5LeHQ4LFa+rWkAtjgCx+9W+gLxxINOh9FX44cAuv2U2UtEJ8gIlbQPcInca
TqxLZ2PjA/kE3/AiDuxvnk1rnts/m8ftUR3o0gNV9ueIYJwWAkpiT+5sqn9j
mBvfNHXqZUSGAFBij+UlISg+AqrZjkEvQ43B77h5qbEhGtgnhKVuSK8ufC33
+KYdtpx+hVCalaBS/4rjjQefOoHH9AnJyuliyR6/cbuJTixj8hH3sWCYjDw2
FJJhwCbyoo3i2xCZdG2QXYGq4etolBb+CPZsC6xlP1rYrWlQypEbglFYFJ/f
pA11l+hAtXl+uIvku0YqJzB4TG2U2qLQA1EeooyJ0o0Z0sdm6/ytwHIh5q6c
U8KIB99CGh9TFpYJQynO/qCVlD6LQAdKnm2v6Pn0dm48c0VI18MHztjNdUu3
1V0NquCdqs6xQZ6gsjqXBSZ0OI7vR5WmrfdvM/t8b7lHIeLucnPBwp41gw7/
6D6//ZL+PnxsWA28cA/dupD2neoZjuEWkoMBhL/8GR2Gi92dIMAQ4BFVt7Fq
L1qFMmbh/UX1kXx6DYRZmSJUHxZGhCOZoWgDvhfGMqmCRYpDHykSZUjYcy/A
K4d5nWwBn6HenBl2X4zS2ovAGiTgndYprkLxATILZOvPfKMq6URH31s+mxKY
gU7yH76ezZtbGpoVHw+REN5hMv2xlmn3f0eKip7SE6jwjZ2q179IIdamFpPl
qZwZuDO9V0EW7neIBQAGoEOWK5OU4YgpWhbAmVxhvJ8Zn/mwb/n7DBU1eKQU
fT+AVgygEo+TIiaLzWzJtHmnh/Fd2E3SYc74zKndCptyQToKnhqo8UYfxZor
UdXBhq7PbhO+QvnbR8KGZ9GWjiOrQlTmDrLUGkAlYDV4DnyfP5mHFyMpwVPz
hn/zU13exE1wj0tmA/gRSOnxfghc/b8gUE5Y7RQbQ7c7PvXdh/3SlwHSjIRI
stMU7mQE6IfBC2OKBw4j8LAbFUkWEX5YWsq09BvXMFTNobmjbpobWFahP4I/
l2zR4N7FXQr+qmoWvtX48cJgiPQFpFnx/HhL/hesG3yIPYWji28b3cNx7CoR
QdOkKu+tTUCJtBH/f023yfKknNway0/yqZ87r+COrqQ28A/Pb/h5oh7RnWrX
Z9i1VjWbxzcryyAXwH4SXVUvrQkEgHS9QXbxrGvzbS73jiOZV0GHd2u0GG9t
afIBSn9e6JOf4UFagwGa2QibpDZZgiKqtzC6jw3APlEk5Oh+/d0qUCsG7RX4
cA8JejQTC+SVs85NkWktSM1fv+aChXQC3Aw9or8FmnjA79exRzSuqlDsdump
lXYvWilLD8GEaldRHiRp4gsxzdd4LQcqzg/mRRnCUWk7NA7ce7EcOHdM63Qk
CEZFHP+K2dluM4d9pWp7u6uxj2DAAM5SobPz+d3LveoNq9BgWhyeyvkPxr+x
j5LlPU57GMKQRTfZz26YgSfbL2mEywV0fVZjxnVsaYlqO+nH4AbIzb29efPx
4exgu1i+82OgA6J7fN+8WyUy2E/QqkBEqItRZ1NabZzjVfaQLkJil2bjBPJW
fA1EZQ99g5lCaU9AqdULHzQJ7kSQsBOTYLoOmgO3TDMtWWJlMO2dfK0/EgYM
pncENfoXrB23bmPsDWANjb4Q7JXHjQk7SQr81QVqEzUDli7DtHWOJ2qiCO2z
osKRBBHUWdUByll52FJvX22HLNW+7AHFwdVe+aIaQePYm2+UjN3U8BQaUty9
jDXNnNgJ5zyuIddAKsGxSNzbsB3imo6vqagHZtsXVMgFOE4GDDQqaxcX50KV
AkDObBMsiTa7fyFyog9F1FdrN5A185I05iX9FLzigOCVNaOwPrZ074jSbLzS
I5zsBjPew3QMrd1nmIZTZkFv2wo+SsQSjAyLycNe/htZgMJrNUAwm2NdPG+E
mPQ6FvZutVEePr9Cmb/gKe9eZhdD/VCCrQ1B6i2pOlK4U5tE8nUFzNqgwDcj
2fNlXBrVuTxv0FL73y7dk4wTHx9aVjAUqiXX49gP9w3GI3dO4jUu3MQfYWsN
KbD0wLixGMGcRbKy3PmqgN7trYwn7nIe6iDzPclSKHVhLqAhurEkLE8f/iBb
ZC4SraO/Xr4CnWt8LmSD3ZlfCgWPmN8Ipw/sw78vZwsFzy9SpZFoqsnS74qX
4ELiQ4an1SpZoq67qcDK1E8N1HKhjVFNVkCR81MJjE0nghe8hYY+/l/NGzFF
W7RYe0yueWgijKMOQKET3WQPyHq3kTff7zGAiuJQ2TCwG3btJc/x/tuKhbHR
9q2Ix8m6FyjoSxiAzLxY4mPQqccepmbsL1wgJ50Ri0szLEczJZsXzNfV/jzk
ZNUkJtBGBTk9BuHIW/BZDsfZeBuP12+Xg8slPYv0fqzHP0rDTjWw8GjlYYmv
Na553vt6qLvnDS6ETtCYZgJ5nMnG3yYfxVH5oirwqg3b+wQ6iNhu4oT6SeCW
BhkDgaT/61/ZSYqiLNIbs0kDYNKM1mDTF3FQ2HpSndkos3FGpUrKgp/NrbVg
QvzXXU9mjfmIle/wPq89dJMrh2ugQayvd/iTso6sMGjXLmvW+omgHRc5FPIv
63AOLQwup+m7kQvala8iOUzixDrsHeRMPena7u3q8GEne3Y1olx0SSfn1gV1
2Z5FoBljcO0WiCG7+NkXFCNNL19ukjEPvPXb8BShTkQb35xwCrV/TSWadHvX
hYjWd+TbNbQ9dkPxXBN+2zo1SzHxmOWgGBd10aI3kYGAZatrZeSmYf1Isyx2
vcL06iYzVZnPYsR0VqYxWg6LEUOjyBeFBvEZ24249TZeMPGX2NDC4ODJCvYt
ZYQjmgeT4Z4Nn5E0elxgdxChNSH/LV3BOKLWDDvXSwdO9ZNU8h8sjoEyVF7H
bHVUtXZiNpjU1htHdQt/fGU0UyzI8BynT/ExPNr3bvD6p53Ut/XhO0hHU9rO
H0D3VD4N4mMZk8w7yVPLP6ORjCF/CZI2fbb/T3c/JGPsLb92ZOOij03GNx2l
OBvoXtompa+zqjfcPtevewuVJ9QpiPb+0oHnVUKwngIOu0xJrMcA1gILT3ZN
lZHzBZZWIAQxs1WiEDd2S5fzli43Fflip2h2Qgc64RS9MpR5NTgrPCp9ViJA
hIkUEbLVXyzjCKRmFqxgaA2xZ2yvtiP/2OUPlSnzAaXHBG36rxllJZe4tQrK
AAWH08dBkZ2jo+VNB2rYcouovxc91TdRWafK0dmyt+edba/9zcPTMCJsWkVq
qOYc8imsRtJDC+OHL8h0/rJOunF9d06ejxlE2NJRGyXQxPQJDWnfssOZHJMl
tTnPWlNF3UPqA7sIrFph8JTw7/389hFyTIhiOjNnA7s8EHhik57x4zkoYvMk
YFlZye5icVa7qSS/rLOfN0MCNwXkovPZnUiSE8h/WcmYM8Bl7YpgyrP0SSt8
T2n+gE9GcIPAzWU5/vFDX8MCAD7HqIHX1/xdlHqsQB9nBOED6SAhkTsBLWXO
t6UyEuadknvSDaQlfYwuz7tz+1dejUusxewFfhAYsgoZcGk021szg7OCbW9X
XgozyDmZZvIVz+C3fxkNxjP2tG6pMBz9Ew6wCgDjmS27LG8iHt/7Yg7pPr6y
2kYCSfAV3siBA690swogakfp7LRStihLjUKcS/MvzVNm++YLezs9ZAB2RIPE
J9DQ89PmyZZy6Ey9a33ZZtQ6FPY0j8SteQ6RRNtXvOqPMWod5oy05pGz662K
CZbyPzhAfoC4pEKvCNYKml9uwD39udqOlW8P4TlnAgZN2Dr24qlgMNpIglcD
57W5rkN5sOyr8e6ckWJaSK+F0UiC2eRwMaGDcFfXZU9lyI6JuJ99BkB0e7lM
vStGuLv66OLNi0D1wZG+6nQFzT579JHfzjG2MPRlNDkAFUh83uIyxesEK8q4
M0tZetH337wenf1udfSq4ABV24y8RW+AFC/RrmVQxtP0a/v+GZPENV3TVSWQ
E6KNLuOaIelQpI+oPMDIEJL+soRyVRe1t/0StCgfVe4PyUhoaJnD0HiE22+i
5Lb2SFiX7RUpxxdCHJgLVIjS+CweImt17/VHqoaZTBu8MwM6uXMh6FWoZLxk
q8eGzrFq9VHfr1Wk4VUTVmQMB8e35Kz+sr2mLnib25wHYV8q0GG2VVQQXHu1
F3esaoXTDJBrBqqhp7+Sp8nfhxKJb0bCxIkc2i2VCx4Zu4SisZFRTzCdAq6N
AZr7HHQPasmO2eyMDwHTQlwNJraqA+bw0kOLd/eOh1lgEBoynVcxtCt5pbYl
zxHU1QASzwaekq4b0BvhPJsV/B6BTYOaz7a/k7kFGUSw2xhTebaP/U52qoOX
NpUY/ugKZi/EiRVhA/+8H/MKOHbuUBg+PPZR8oDxiAuerJR9HHiZr5eeeu/o
q75/rDvNAA5BE5jgkR6I2vyLnoafOejJ2pvcNomBqBkahhUWEW/9VaEzwHW1
Gt//NGDGCLEJDVh66xit/5m9BZgcNaXhUKbRrI4uBpkmLskpGNNWh+32aCky
HhRSX51ThXcNonh7gjZZ0sVGa7LIN//tKRLiWtNgZ0CkLLW+nBaoBHsaaRcm
eJd6aCCOfZYeas8Rs/y1FP4gIiSX1pmxj2ggJRMvwfpUnlH9H0GJlIUiN6hr
ifFArto9sL0KX4THGVNYIF8ul/WCyaY/eZikSul5MZ25AvK52VMiOEs9oQmx
pd+MkTc5lMSTEAMMRL3jdbyKvUT0qPMninfrrDdI6x1Y5JnXwKaqM7Yo1LO9
8y7Y1J1FIksA0r0Us9xIj9ycgqTFxPDayDEfxG4974Op9h7v5vzqyk0VYffV
fiVlKUvB00uR5OLP3BV1eS9tri4ch8HNUQ3ojeSXIXgIHS1hFwfr0ipGQLQ3
Fepn6z3+mjPflAuvp63grm0XRwRkf4hhvI7Utsa5aVFtFn097OlNewemIsOt
JkdCXDFGx2CB4wcRiRIym9KfRFf8wcHEA7DB51nyeAGdFaX3XDFG/sVpX5cq
KZas2pSn95dxI+e7Pl9UPbca3XpPWkVBG/AfEoo917D67hKeOYbjtu4PXJa9
2tylZPPp/rVNQCnq/l1Fff3H2DQtLf+5KwTJSEoWHDch84F/U8RUNkXqfwxW
tsHwCZg4oYDE5mGt5Mxgqz+vYi07Oeb5QhhqFz1iIjHaFtF6Di9blWn+uJC6
r5ntHpkNfkfymQmjQBhKdoijoUf63En3MXsKMaA6QS5h8ARM7Qpo/2IdOOaC
E6EgOBphKv/tf8Vg+9IwESmW83WT1TxiYGMcKgX9qdaCobApRMyEQBn3wMiw
rGOFXPyNqLhtJzPPnVAo796pbFPSsdKmIbObS+gqon67K2FSMyC4rqhdaVwx
6U1uEuXdHAn6sUCkumu3zKZbB5Od8ZFZSLEu/Any9K2btYfv2IepgVu1zVjM
4/tcnjRqUMPSWhcyx7w7tAsxRLyCot1ihS/WG8lSDcPrqHd6X5dl2WeP3VzR
zdeTUVXpT5SAUiKi+gRE4w28TFMc/pJC+aFayjudak0cVPvTi830UzVkzIxd
/+99EWIyFlQA5BXBidsLudDmZcePvrUOwVcHhZZX/383KCuGBw098VLBl3Ui
QQ+ggMJTr9XSrPSv4efUNbx931ZTQDxJm/BVxiJWgN8uhOfWIJI4EaZ7ccL3
B7hF0hCIwL7pWNlzojBaeuVTU1O7k0n3dblzWMdBNU9gpSVcTAmBMG+zuy2I
14Wgvu99qcH2Dz/rkoFOe/7lRhFvrKtZ0JBWM6BoUuFPkPf60bMj06qczKg7
8NkaguhFLWt6Bf5Q/Lf9PtbYbz4xfLasijYd0B1Ezju1ELO5HDp6pfGkw5iB
eV+A+wMZqZCKIExXAAjrBU0aWkLzqDrV0KnOsGiETUGakzsIHxmXz+tRBvLe
ZTttk3SdEsNygx47moQ1SvTlln/r8HZoagNb4kj1zMlGMNk+xizArva7yzvF
0ys5Ln/F0kvK2CKUeRBJoFSC6ZcVvWhdaVGSKty2hN+Z0/ahWnVVHroKD3y7
JLrRMfR7kCprA0U0PgU/oEBRN43CjaieDQ6A6CvhrM4oPRkMSe9ip1tLT4a3
cELfuOeEqJopuSJmLwjxePzcc8VynSaHjEfeK+3QL5tKKmvjAE41mM7PymCm
chp46CM6NSZv7x2nzwWfPapjy6wLWH+X9q6EiKJjzFrIinciDWXFfHkVJFVN
k5JJucw2U3Ejk5oTTZ1xG40Xmrk/b8rs5h1wAU3NYmAm+RRerWvM5d9DSQoj
eV023w2RxwiA0SDS9VLZQWCPG81s19FXzIP4/EMwaUFv/tlWXWMB6w75AqnT
7Vxy89tjr5Fu1MyBsmkrAHn7d7AZ+D7sCk4VE+OypBd2jM3HvkdG8mKWo4m4
juC4rutxIzDCK/XfbtA27Vf9Gc9e0Ew6psnmvyu13dIGaU/yfudeJzePfYbg
q0YWgKmxe0xWEs+hcq4SepceaiCDMJ7bvxGKPCFLQjmTZSsUbNxF5DjCajLU
axD94XWkdGeU62d4jiyZe5EUNx/zNrbgtEkl+pnYYP1edo1XLf4CX+y+i5t+
M75TKjrJj7nI3W2PynCD7d4NQ4TUJKk9GUbpnj6JXItK0jhHwiIORKMFxBlg
FSCpahp2KHTOrXJ79dRbzAD+1NvJ5jPRPAm8fIPeG+DINg4frSpuutncJwhI
bZdVURp73qSmkw7mGGnjufc2soaUoArWTx5zwmkntuybii7ORMNAZy16/ABD
jQkJEh5gEeyE3cxh1IFGvKtUwVyI6YrDaSTbHlUJVWJ/IIeDx7yHdivpio8D
+WqfZKkMEnrjLTUbS90S94i9J5DjGlalZX2dlojDdn6FfjKiUINYrVqZrI2G
iDKtrxtYZxrYHDze8dVoZa5VyLVsu+Z9iCJ5QZn3MeMUpLW6jh+W+y2a1Hvs
fH4rk18MZ6YywV9Gsvhn7muLR+cvjFCre77f1+xhdutEaW+6F8auLIZ7YwB7
Ch4TpVRd4K9TWGrk1eGTlO46HGw2Sau8MUg0Gu6ivB5ZYvgZnsZJa0O7B0dU
/igS0Sd12F5yM2UW2dZ4iogZQEc91bdG8PtQ72ni89d40bV+7ImxBrzgm9q0
tTwBM57sAEiWZzbuJ3nqidmsIesK24nDl8O/LxIod4ODI1cKyU9yOBxQyWcZ
rdTUuuR8pCNpqaTCaXV+M8X4+sypGgE9z/bCX2iY2npiR6/uozlm/50bjMQ6
PmWSBaAvcmN/Z8F0p4MHsZfrdWxjvjaBF1jzFRiWMSz0gqd8aapT/V/xO9Rr
zUgmksFXwuVfUAVhMNh74Hm8BUxowJ5CY8KNyWaVdsO5245WPN4VV4UsMI2F
D8J+DxgslhdSpYlIdxmDZBK03ZkXZVnDoP8qjkPgfrBVgQoziinqVty29X07
PYjt8n8bO9YMZzQl1a5wTa2lL2zEyKOpYja/xnM+mBid2c0gyPdThj4CM7Ak
YEcuGF50MnA2TkE+XJd8WqNB1cufce4oHlNJE4u3jHeHIYOJf2JS/bvtCYBD
e5RbbmYsDVw7PnfKa6tOpEFFKoqUhXQvj2qexhdEijgNAhiMcsdQzGQMljK0
9PtSFgr4SS779cDFBd8vOBb+m/zCYtasfVOxOM7ttJVRII2xDrDxQCJRFlfe
GGRAfSf39IUclMHCPJzrfdTI+G/CDlP/7nglTigUzOmgQEWGn9GNVXMsS9Km
v/BtdbOqoJ1dxOw2c6cB1zlVdk1KGrKK8Zxkhj+zYS4HrH0VdmZxxffL51FH
yWmHxu0X2Xj6oW+yCYGYUwoDQ3yJDnhIgStD+gfluUs/AjM3b/xhs49DFs/4
Y4NWD4UeYACoY2sDp8BUOpto6idviDY6P8jt7n47EVuFJtwcKx4I1VG/E5Qt
NiKOaWF3DM7IDOy4PbjNkXWSmyP0LVso32boFjGJ3gLOrKD+CLLNKLtOWINP
mP641uBJvO094EYasI5xFnGDGaReL5x+U06Iux33gN2xuNkVyAGTvBcH5npA
a7SnEA0QUr41qv159cHMAy/Qbm7C4VONxwqLqQEMNW0+9Eprj6X09590I5a3
lFdQcFJ7pK61mnYuZBBtCmxJxR6eod7vG4zE4PEJ+XFvJGV5QzlaIqzSbTC4
mjql48aPZ+UBmyLunB6k6oGHYuaAk5gHbNMQdDemI38zoZxz/0s80t9bQAKa
h5rVVOJ6BFw46KwtkMThL1Mh4fBA00uHfO7pUPyJbjr5LY/GoGFnG9V7TdJr
36tmC3t+HK7BUoDebNv/WgbhdFnPF4wDrOuPvOYydFt/CrprkSnZTjwqiFVG
JjY6YzprED+h37NYAcWpG47TTGnlVLrVRM8s44eWi3i1y/4azy3ZlNCep2zL
QOYONJOT3A66FjMzaF8U9zQZShkwgVfDmfjt2Q0W9y7GxPfVmfSFSJ/oZuKy
eoswql+6ggxx0N9xC7LYUjCtlL/GuFqV+XlOcy+pxGm1nGFGKmYv+le1uRNj
4iSxt6lO8iVkGf+5Z6KhHoL4EH3h43bUXa9RKQ2b40gzC7aziP2NVdn731ro
Te5I9Q3P+ARhGDFmcHgYq80l3PYeq1F3XCtbuAeOxveweGpxECGLz+KDKqFE
5b8gwJ4kK5j9HD7eKtvpWHr8lUW0wB1YybUowP91UFxKilhBHUMpBDqgf0vQ
tj41X8gU00r3Qj8ngfkHotKQMtzdDI/sWwtPqO19UnSp+UikxJl6+2grWnhc
SqGjuzr4ZPrnN35xJqxgd4gPTYlFkKChQ6kZ+0W1hCtbqVqeY0MCF/N2BPbI
YP+5tabpzcwKTSX+fiHi1ox8zTf4Do7nGN2Ubn27Y4Z71CqAWrNCF6DKtF09
4C4DSOWhf88UwEnYTvISkDOeJ3UGSGBXufYbhs+AmqzrsYDjvbBg1ncEJlvX
c3/Ws4yrZlFdCTlG9Xd06XUrU9qbkUVauutKtewwRo3wUdnyXewzETE4bwwL
F5NPamcOg23tgpIY4n5kdRdWS0sJIQJhkOH5qfb+tB5HiYlpnB0FuAMNkJTc
qHQrI/kQSOM9PSKMgu79cIaXg81LqO1C75Jre/PPvw5zm9d7/eAyDFW0cRyK
+5bo1Az4qhJTwAFt8CsLm9dpIlZFCQJgok7/pXOSbDczKVq5XQ5DYz9CCcYs
arlxioCdKot7swGxMqb8kLq8YlkZjbU9aVVIFVrGrdBtkSWTz5sfhCz2j4Tz
cke3Rd/kJo6D0+YPSBZL9aQJyr8FhNUmcpu3tm/EyozQ4wmTCatxHpOhJ0HP
F+/k/N6ZsTqO0k/MSrm6V+shHEnRmWG7FmsqUKMPeqwhRMiPi5Y91l9VHvAP
xzAI0zzLS3+pTvaN34AZZJbaDUTAV3f0pIg4/Ws4zZ7kdjNm0jlrtdp9lvCF
IPZ7QhvjiKaZX/gU21BlOgN70qjdDG+tfzA2uUky1tOAdeAKkAcvWkkHu1VU
jMSCzD0xLFYJnHz5IijtEzHsnXLOjr8sEqdDMzCOQFtZ0xJbqOJoJ6zg0Xtl
8AQ0ocN75thIPHYQidoYojOuR4eFpifuPoLAEXybq0tmOey3P7m50eO7UxQi
o9noLJ1hJUg8XWjjl2//iaRr41QAbYn9SxLf6z/B6I0ZKVkUocdpWeA1ozET
/9IutOOCz4ClCmQCwiePIryMGEUBgR036W3b/nlAmCAG1CDvo82IDb5Wod34
WErE0TCQo5P7FDKj6VbNx/kANTi6tEnQXNYNp76JxowwI1Z3iBV9CxAaxeNW
3fn5WHGw64y8zoLzpXgW5Zw/8YMtUhEMz+kg8Xf6hJdvAQPWlXYGXS6BVnc/
f0QlX22+dbQRTtluStklJzwNJEq6uTvExeBkmB4QaUnljQNRAKvlY6PB6lPx
vyxmOQ1Nchp61Ijji7Y/fA7PtA4IrGk4J73rRDRdYu6jecDK2Nb7c44CQbrM
iM6xedvy9iLInX9l0VGAEPe2LRAS31mBeMGtsG9uPCXiaZNtSw3EeRG1SUOA
JbtVDkUm//7x7aE+msbEUZNVqLja5EcBMpO86BOH1p+eEKWzHCFldAKZYENP
kxindwWRmD2K5nHJiK301OS40Hkac1IuFeHcSnPZgCNgqnaFZqhWX0+q8lK9
pMlbdeuz1ul+jUklrqBMoaG17dtCYkbwt7t+xRWF5wYoSZZNIwTL+k3e6iie
EOrZzZjbYIl68LWJq/nX7gUdaO0HJTTKCqU8k05q3BlERKxJ2mgMja5RfBCw
jLMpj7Rf7fDc0XWFh1wI2snc2n/4yfFuNq2yZlN5aRl+wziRrYH3ZS2lZ6Ek
B1oUfbWEVjZoY7Nc++PNLUkiHKGeJcOoJHRHtsRieHQ6Ibta+CHMMzinyTE6
bCspQo1q02apeNSQ/fgdlYtBqlxufDnD6vPunY+vr2/bdrgeHn5lQVp6hG5h
c3zGVN3dBO0eyAZ577wskr6x7O25vi0k5Hxzv3OTjSFIQZ07ztG0ICE+gQZV
IHslUh6slFPNvIqJXPtJeAFx6K/vvBxPonp3b+CAZV8Ly91vzcE5MPnmgy1i
0VcHwBmfHVlQ5Cl6CSom7LIBzQNj8PjI+pR4U71zJMEZRNasJkkRAck6oboA
Uk8Dede4HsdLVvJrnbxZdn8gzyyrc+DqMPX1YZvf4NjkirQy/rhivHacFhXV
i/hVyXwvkwbZQWpn4SF2ViF100amvIebine+8xtgkxE+VtsYBueEYMpLn4I7
X6gLpL2SPcHu2IiB3v5s421k8k/WeDur6XubRs2NEZGEhNIJKo0dH0eElYv/
aTgaNl0oP5DUZPW7cXTZSQ8dZD++HAIdpgEcLmdynS9qOet9rgrcBBJgvbLL
PnizFARe1zYyjxGPGVGWD5BGYnHdLgaD5X3k/GjJXp8eCGQM5ZXplg9pz7NP
OHJBzep2O5mo7NFNoqm6jhA4QK13gC9Kb2+ydHTVk2si2wttPiNX5si+Yu6U
X3lp3ivV1JjnXWroCHqfe2swxjcNzoLx999sw4bt42QKcQFHpVzB3h57hIDh
pWXDSRTFUKdN4mq3T0eWwooPmyvCycTsgo1hN6h7Y8oQfTIIzER1PW8tolgI
EJ5HZr7LOUPj3vxkqIE4JTOdcvukBQ3Ub0s0GFeg9YHlePnt4moCWQZi9ErU
C1g6ScsxDKjFVfQ/+x6STeyqotUjfAYQU15yOhTdg8hf/E8IQIFjCQI1CBEz
gKBVBJUKCzru74a1q4PG8fKniJzBm5f/K5hwMrCo+n8Mkc8x5eHyuv/Zg4pr
zcrLi8y8LBUv6ZfQSg9F0PEZl1R0xGMNXLvvNp9UL61j2ui9SLL1oTRw0cht
mOk+BFOKy9ji5BaG79NoF4JWJindcBAW0Cvx+FdlWANTX6wLTrRdeXTvxV+0
LjjRE3H+k/5EOwfE4bfxaRIUpmQl6sJTAHdNCIeCpnrWT1dtCKwouuTHcGkR
FXGr5i30+KeKMqvbPYI/Jp1gKJzihv2p+pqljH6yII8w12CIyVpf+vhp7HL8
59yZCDy3l6MRpWNnOKbyrnbp9PWaB3onJ82WvESu6HXvNWBmvj61NbkfIR9V
vn8cXR89aVH1Om+ogYOPQTox0FK4zMtKqEhontWOMapuMjQ6knrzUNXVruKS
1CcdQQhqH7WYmm1cnyjx4c7Yt/xa/5l2HPjkUESdtxf/BMS44BCNmICmZFd2
I+llNL+n1xA+1SQ09hlJDkr0XQ0+BcytKYMfiTkG4SPRKxGS345LQnRHr8F/
DYW0794pjO2loCo2Z3F+vk5Ftoq1QwX+7GD6iFiYH1l1wyKXGdwrt+cs8N0J
iq4XcPulNigsMIMLHc0NMdT7cfOQYQrTb3AwsjT9RAwCpDsL8N0jS0KDmp8E
sWiGziMLQ17eAmYVlyCKQzuEMDwy2FCKUN+GDlCbxIYr+elmXPzwWZi74DGF
WmS0YbkqTjK8HxW2yWMGbS+I/Vu1406di85Ik4/HV/K071K+3LTQXBZiXAA4
aTW/EMNoVg9M2SiBa3m4WrXDjZnmPdLNhhRilWIUQnfa7xP+SMU/6vQqCV1x
r7vvf5lhsUzFc338L8OfnkdxnolajOo0G0+SrI1ICKWCpq9hq0jKjfNGlbWF
UverFkfjEHr2EI7TNgj+aasTmLL2coGgRyeCHF4Fmes11QdHG1c810BNf62s
INSvvohJn1MqN5wObBhJmjBomktW4eum8/xkqMZTZsG42sTtVsQz8aT4eUe8
yN6mG0SvraxVtuI/Oly6w+23BmYPjsobiIXvoSwcb53IAG5dOq/v5JaN3UVN
pz8hLX+KETb4PwaoVFHPgp0CoWXlww+7KQuM5Uhr6KqEK8JjOV9P4c6n884v
kOs/BoeIicVRvrfjOhN2r5sIq18Q8l90IeZPsDeN6Z0KWk6Y4ODLR1vSQDpP
XL2TNGUA/M0BpJ+IozOKU0ipNWaNcSkDe0QjGt2fVedUdOHjCupAUheRH175
pMq8VLqc/fNJq9vYfz6yXL5H3WQEbWk8HJ2QUGKZ3WUetkNITHvzJw9Te0En
hGeawXlnomAIe2HdFuovoZNAaclJionzHcZ2f5W3P6eTOAkSudE886OaRdt6
+usKrotfLEoq0W/SyWNJqZQgQsUmSHG4bnbBXwhH55ujwQxg9SK16VkAArdL
vHPJ4NZZlSqOKkDLJmNfGRQ0BNtUH8ZLVt1UGAZMtHjF3E55OoOJVqd7Tc6Q
DMhEGShb46Q3cgevlrsAuqhkO5hdOxRDJXkQW583DkBXZvElKMBit6AHoNcY
+JkluV5nDgbrPvWIv9Uxl1oVKaVWMRY/pLsLpnKo3HPcxz46pFbOkIJIVU4t
1YKRzjZys08B3ImhHZuumajBu3QYs/DKQcLRwQZKruy154dRCflaS8wrratL
QnTkK/ETOPZJJQrRlOV/Mbf82L+UKqGt5/70rlcFUdDBfbVAwHErV/5grOHo
iJ5UlqseRzlqRMT0dF553cQKqbRd6lnRxrSTs4J1cFfrHO5lwSCWywEWyg0r
0mcFUCy5Q29Tv5HJdg4ZLPVhwA5Uegyc+fFGePPoxoX334T0qfGEjXoeVl+l
uTCIt886mlx4GbJ1VReUv5eJaVpFmQdZko2kRz/awAFXB41QaQr0VB46uy8u
2bWCdXJ521I/weZoZ91xtFrpBSJnLNzA7Akx8yyfN/rKuAmAt8MeCi0E2P4x
/oufAOiVYhe6BZ0BEgZlGc5qz/WfWGqS+NXzcIe4oee1WF2leN6jKK6gYumr
BU76lHcPvPTcsvmu/blt4qtcT4Vas2jI4zrx5CfBTzkSAZuBuSVI7fgYp81X
0mWUOmVAJOHUIONutm1MT7tMylWFmIyQgda9NQbL4uW18hhO0Mwje1HHWHae
et3KxexAXLPa6siYNya0iZvoWwMkxjZ5smDPyRp9o5YZXbthcz0juAJnIpLi
jtCQP/h9UTpubebexpvx5mt3VxKEnBSS0Jg803c1302t60jmWvaa5tOf0Z64
7bNx+215+wujPQPfu2k0ae9DXxAaTKDX1fssZQSrhp+8hccRX7CgOudV2mSY
bSPJn+JOyBMXnFAeZxeV4IuF3bHWikZvwZnDBzs5BELBkCzu8ldDHmdIasy7
JOGcKbilDxAIx+Z67QCSufUpPeCbTRn6zEH9Fe16ez3tvV/GkxoxSX9DuK9O
0wgiv5rvlXmd6pqYPL9C8z7SnZglGAPLTke+Q1gxlaJsikblGA13/+J5hqhT
sLbVRHaSZZMWKdTlUq/Mps0xBk4t+djQcJFIBal9Sf1IJY2emqhf+TCQxS+M
LxHGZYl4DebnkPIYMBZ3aQlkvpgLE/rrBIGrngNUW96kU7h7pLJun4daNe9u
qEhI5oWd81d1fko7chyAxTaxYv0pwgQvpEhZ5abo1LICeKOKAfVgo3g+BAtH
WKU4xVMYPwnLrVnHtBWWX9tpSyS9g8uF89MocUNg5VBzYw6ueX6M2897FbB9
uguCWJLo82U0olQlzt/+fwMDdgMGvqyzXYfs5Ca3VZn54fcXcafVFOwDVCJD
xouCLDGhPQtqWQYnmXL6dCvmudKr+U9ZJ1l9+OgY2PaYBL7e1RXA6XsJFGD2
aSrJp3WYcfYq7yoeoTg+OXT0E7+I5RMgezc0n7l9J9yWWzTiFcKovEkGgYF2
lkiG0o0JZsCGCBCNH7Q/DQ1s5/W7ls+9PF4tBcGC6O8JrGwQCpdoXj86SoP6
4dQEazPJfU2QkBVD6+D6+Abmr1byxUZcfhMX1OTM4jFfhVBI7zeCdaNvsF3C
ifgHgGq2xlyW7PIJb+H0PWMISan9wwdyO3l0/f/hVIB8oOtgNVHUXlxycmkC
nhKwWIfyIB8+4XgRZIdIMwSGGtSfGmFPcJsPilluTgBaRqIlltsic3xIz6OM
7kYUHs1/b0/AU9m4TuOnt6GKkXck5VeIceG+xu6CzPgho2OweWnt35jpK6ys
Gn1lrSUxY9h0LTqH9TiVHAvt75hluoAj9Ibk/Nu7Xp1jERafEP6mPt2QtUym
W/y+4KO3/CAWk1+/ppTQKXEAecRmxsCb9nzqZquALo4FvHhxOBU5AHT0Oqj2
LYXVQ4ra9L46gakzAdBBo6fRbHdVius1Gf9kgsLFWQ+7OwjzK5PBvNfSow88
U4kuwrXCjTThAeephREzED1FJayQHkcNJ3CGccYCo/WZ3Afj9Ooy+MP9oGHc
DXqcdPJPpc0v40qcOVHKwcNyN1wUEaKQe/LUzMTuT/zKkU39RZOEOJVxTCVW
bHkUNDu25Y6Xcf8wLfQTE2qhtRITJD3lEuk/lQgP03sKL5T1883kd4cEF9CZ
aX/gE9eUFdw6epJopbiQtB+JGAh6wsjaay6gsoCBxddL99gRXf+ZOu9CARbV
Qu6lEt2JYTEw6a1G2LhqhcEe7Jzaiso8NhvBTsGxayCig6abIGdonIRlWzhi
gjr1z6GtiTeKqGdNrcpg6yAPuLd/VWXltOn1tGAlFIqj5uKhzZT+wBrU9Pxt
wSt+RJjjWvY8eTa5y2/dXo02XHt0OiEE6L4UbZmRl08hqtOu7mXgS+PcBKBc
QNUsTA9WIBE0sdAj99bKQYe1aNVZtnHb2IQnJYes0Y5ygDEnC8jQFqyNhaOd
lerQWcJktXmgC4uI07vQXYZhfRkZNv11z7OTi4MflKKsk4Rlk7CLvKyISgZp
3qauZFItXkc9/Sw12PnpfcH8RZGKhFv24ZGCniORX+0OLORcrPS0s9m9/aBj
KyLmZaEaxnhr7tACt0wugk1t/kmgVsGwDELZ9hWVjpYMI5XqtWlF/HYT/okw
c68Ba/29GwY/JXsbToFFTfMicaijQWKIjDZv1wJxScp0aw8y0ZPUc3ik7T2Q
QVjplsu5k8DvUKpDnFrD6yXiKDOYpfdRJoNqRN0BrpHJUA/G8y4qhClyJztz
PZ62ccehxPb3DTWsoE1VKcFOjIFEWwXSA+GNn9HAaoVRMyy0k/zYStnS6lC1
AMj0oCgBUEiqti0xeEh14cvWRGMKbO9sSvASJkoW63sVoTsSvXbcHyYgm89y
3BvCx48zUwDvVpyq6CW6sbHykvpzRNBB+s+UjXfsHn6Q/Fi86FljprSB3F5u
Yiic7FV0br3qgVQZio1Jc6AfczYQFhNEaDpqOu8R0ObaqK6/Q0RUue13n8GS
yehD2ekrMbhFOCYpYNsKWIsIBQZndVA+QGXjQ/xhNEqyiSmZU7tF6Py0mCFq
AKJfLgnDyZdczwstJkxa7Qq8M8dBFvXALmp1NfsOo+P4BJqvNUOEM7BNWpbY
UGpJa66CDVV/+bl0Yk+qhb5FQi8Io6lE2xmRw+NPPqlDUlahmmx3mTz374Ff
OFCxyMvoP6Q7vsO86Et4nzcWddttGVwFfEcU8pHUqsvqrhSlVpx1QjDL01Jt
rCFlT+lhtv1ZOstAQRJId3RcwesjLSHlB3SyUs31fROjjaguN0f/bn6dTfDX
1Lciop5UpPcnmG3+VokR7fwnhrRFlUM3slnwEfflB6ooa7o4SN4Fr+SQC3el
hJ3D4p4ZDMYCvxxfXdAGxd36T0fG3a1lUyR/Gqm2oYP9FjLnesSpXrdiK4aL
xzAG9B1h85SDHjIC+fcMNEGMhEje5OxWKUa+HIzoy3IvqIK3QUCqnYW6L1dA
5+rymDBxAZ6ZViEov1TdOeGAZzWcgynBbiqG7+iN170dWWvlSbcsNCleZkYJ
ddDUxPYt4mBXOSKyAmo9XRfj4/of+/f3OnKq60kL3WBtW06vQNf7WueK70sr
sx0g2lxycqK+u6P8geaWkT0cfp9bKIyboPL/hmc9eSwhTKha7bnE/VsmT7MT
wA+4WZ7Mv71v/+ylwPasyXFPfEGzo2NmdfTCfqWjoLYBAI7i7dHaFzgTeW5f
iAHNvssBdf8E1jk7SaYsYL6OVch2Ec9WnWL3WhGvKqVovyVkiiQDZMLrhBsn
VxiKnTa72VpoWrQlhkUQH6R+jB/H4DAQINe4BuH9fR0ZpBlCeIYrIbljy0M8
Sb6vO7JLeSQqIV+Tn9oGDvHVGiM4QAEuutgstpyPQa5tD1TvTLP8uxhkUxK8
BaCQ/xm4zYWDXV1IN+Mme8AlOrwDfadM4bOrFqF2zuHFmeemaxySFd1Uk4jR
Rj4VtELIc0M0b9CxxV04i1CrErE6S/wxtNA15ywFNkzxc9qULZHaSKGy3TU7
DHkBhjDjjsKS8l9xqYUmwpK8kYfdD0znu3zSBpyhIni8Qn1ApMvHcYgy4q/2
oihG1sUzFRYuRbmO6qO0MlS5ZUl3D07N/xxUfp+gWxSfMNzhXar1NQxpoYtO
hlFX2YuXYSrXTPg4sT3mbN9jtmh7KAs4LtwzedgEQy7on+WVZF0i5mhRb7Xf
mLfoAu8+Ys8XGz9idcfLSZzvJwoJevAoNH2FYGIf9pOFeJyFej1NtsBaqyct
7RW4dAK/iPIuJ1///xyclAKBt9cumEfzG4QxAG0JgWqcwoByTmnQXFLFfD5G
eAkIZ7gLy5pTpZI2/mfJOi5lS07OmFLKGAN3Eouxv1Zhmqx2E/ROh9/0AoJ+
trK/wH6T97vazKl4Hc7hKLPLCD3mQsMUhFzIpPfwtTCxzovARJdwLB7uWKey
jf8hvncNu65JfNBf8XBkZfVBeBa/OxucFJDoMZX6mhV8Io0B0EVHM4RHRl/G
RMMUpU5iD+Q9u54aWG1bJEg7u8ifpfI3kU61QhQY9mBF7m3Zy+ge5eVDAzq4
X8f5RYAMtL5+UC39+vk8j9fFG7HswFlep+MSSkUt4zbfbabCXwBtMV7hNe6r
B3a2lnh+jGuguo49VKda9V+NP87I5RxSBUUaJeJwFkL5xQuDhxBeUI4fcZPD
GXqx+GvU3D2a6laC8fx74MsyGhkXxH9g1WhonYqRcfPAMWrecqRaIgAFU63Q
NPLouZ32K54c5qGBSh+XchMcVO/J95lYjggz2jCKOsLL8Go4JS2BIsFBEJSh
hiW5uHHys7FvX6yQ42XmfzA2K/wfPhzE4XoHuhl3U+1V5j7huXqdC8ok5Lyj
FTMlIaq3fA8vu51MRWbx5FDeKxKsb+laXqFHf4qvOCYsM8CGYuet6gMsCdzH
ZO7O/NkHkhZvjDbYt1On9xPFcHsC/c60R5Faoru3BFv+pHJJPrGee2Nurrdz
P3ca2Wb0kVKqs+W+dZz93as5CZw1jSxvQNRS9L/Ks2erMdDHUKoC/VtFN0zK
m7tMR0ArDTL7LttBrCPqV6W0c1Ws8qMvDwjyLxT5zwKsTxJdusgACTQAUrzY
kx3vJMFha/m/YSDX2yUrCsmchRAmaxEPtp7VeApegYC96XjsUobKFzP6pD0D
LpXZEbq5paIOMkPNmDxGSbFyUudJ9zdHgeawNM+YUd7+TivNjva0yeGIP3If
+OruAH2xy/9vpakENJJFAovQuZy5HrbcWyCwqJ/vOCFU5iOfsTwrZ8JzpHzK
pm7DWHzrBp0sUbFWbOSS11VIzuHQH+h2yCLbp7Gpu8RqLcB16xzBRzqO9Avm
Q/crZLc8C6yew9dIhWk0FudKbXfKI/groLG9CHhepWuWi9+QQ1JVA+UmN763
wWtTMlsKYyz6akQVS8oGnYXN3ireShrFqTFQNg5fY1NgE3deChiJl3mQddPC
zlIFaUP3+8AZGvRZEqMdo6ih5Mc6bR8eYk4wBMyTQ3X7t2B0eVkp35WS3iZW
6k9uGDoTT9te8Dt92XcVp136RNJYXhOd7T2hGWAWi71eCYpzafMnZM3ugfkP
hzJByvX6JDKBRyAig3U0lpVyrwqLjMPcWsJKpUIKypzcOr1sd29UXGXK+xHe
RwSkXUtb5BqOBaB/Cjl/LyBoX/7fnmYFgV3dtfE/mJQks1BgrJiEp9xT4/BW
GAYA5YelhPXBTuC2MwCK47zburbxYs4VBo5Px/y7+Iz+tUmOAmKbPNQaPnEk
ZJPdE1z/LsURsgvxegNGZGJJvolUXGWaNQlmGgBCHBWJUSyCdPjLIQw4JzOV
j71UP3akUb++xOQ3l+bqtj3UDI30SsWm6wLleuaTHRJl1EhYVUpgUB5Up2S1
s7GmNj3JUXgMgtVPKrInkHlSB0ual7ldiKpq5K6l9NBHlXni+pdDis6RrpU9
BrjxXOvtkpJ6fZ9HggMnbOALIWrdXePWmVs4bVFs6zyeYZQpQasmOwQuPif3
aPYdwo3+J0bYJWSRq58mGUMpkySE4af+ln4WJ51IH6KYfcnxxwGzwACMAqN2
x+2dg0uOizoJKEJdPAAI9Gp7JxK3pvJvcLIqbXuvhWGLWyd2X2KC0D2839Wr
tFKcil16tejsB/DDiz2NqaeD0Zd1RdAaBRQMUMOmKb3+HNpkPHH8TGy8wGUa
Fa4dOBye/5OHi3WKCzJ2Fb7pzbfdgRZmmgSrhNAvRbSw2h82n+V01SApzGzV
xTzVSSeHEOb4absb4QYPzWzdOXWEJ3B7wcCxgPdmwTF3hpU7DqNNxpy1dCgx
K3xgBKtTYvjJe3cMjdjm1ZO+XlZ4CCUhfRWjvv98AV5C9kkG4AJepXoXw60U
bhPsQZVeYD7yKG9W+5deCKPS295djDsoDr/ZFAiLRwo5EYiY6OrYnqSKWmtA
9+XlgRvDz5x96mjsY8pOjK/sAOa7aHQb23tEeeQDw+rscwj85vIHhcVnP9v/
bJKbYSM3nPHAEy1BLf+w+nvM4rWZz0I72Kdfruw0WxLqumUDL4StaFJQpLGc
m4iuJ9ul5CtXJpntBDdLslcXp/d668JKuCJ0mtYrKt6bXxSSKiLziOVSR5ga
DesLfTb+dX+fsPtBBcXPk0L0f5LPCrp7d/p8C42k9LZ6fHQlTJ+u34HuRH9Q
46D/Ovy8kCFa3gcEcMdA1UmTfQ01wsZX4IMhZtOXKS699Dg1VNNWUdxulCvI
vWONjEU0RnH4++lkdPudEfPrPnnAv0M7+/CY1SSWSOtL1XjLVzGyunABfM/s
9/VH76QzPHlGav9SFib3KpAmzwQZV7/+k8X6XWct0+ppivrq7rVbNxTFsQJy
DpnI1bvvtGZRRBZiVm4vkDhODygVmECaHNh3ya7H06Z9WeB2UJ3U38wLkYKs
UhQcUmmsuJxen6KfIUAqsi5SF6yf6fCNP2H/mwPx5sw9H4UTM2+Vh/N1xj4B
ep84olP9GbcKV8o/Y6XPUBwdfeeQ9BwjSki4ts2Z3EhA+Zd8/xfwEbjBGUlf
voE57AI8avPFMTuoPwKTsNavHYwkUYCOOpLw3gc/GUH6IHuNuISkBo/HDN0g
/Qh5W/9zZVx9kPRXXIc2VtDbhdMopma8d7h3BaGOo+C+YeSsl1vjlkBI7/s6
9AaK+sDT9sAAbVhz2lLjnzaNmW3bMv4Pc3dbhddMPIGupVU9OrxkUi/aWPME
ZWoVkXU0FQ42SW+fMPhJku2oKyawknKgro3NHrp4FIaMKE4yaNGLydR4PLkG
nRcMg3Zy9a9VLZrMg+VZdLoRMPnZV1Qv8ENYjH77mIODcn6OovNFq7WSUp8L
a8AFSEEtAsb8tLvDoIIED6aZwjlpKur/QnRPTULO36x6pWM61BjiogZI5WEL
FPIkMFP5XMNocYiAhpIS042cSd7qF2LefqdxkX/DHv/acwefQ2lTBzmU+qqe
BMHlNyujEsxcbb8HI2KVC+hDlRG/m3MIVx1Cgfff711wgVkuj/JH9HZW2HoW
OF/rjlOXdZn8fSp5SJitTFFozzjmW0FrXY+n+Bk8b/RiTBI5sPhaDhDaC2/S
UQ642mxZAms4GTFAJPPU/OdoqFG+5VBN39rqvZ0CdS19fm/B7ff9w9P2GSCy
24cDBfDKJe5T+DC91/34Sa79JZ00YNtqr21+IEmlk3xa5km3b55mM+0Jy82g
Dx4/EpFy6aHxL6Zc+oaFVW+0K6c3vDClphn9GUcH1T4iR6WoKxQeDGKnLMQG
JzZMMfOd6Z+yQPkC64QKvRu53oA7vvQFGN6RVRl26PBg87Blgx52qjNuu17I
o0JEetWza8JkFml7exAxy7OVND34RDFdH07XhFEYaWk8Hkzatw3HAlUNJti8
EvH0FQWjdpC2kkTk+3qexfiJGRX0G9avr8bV37nnKsJS77/YHTGA4mDAEJE7
H2TJVHJYF8xad+hAp5oMJALDo0m+joMGUIhLmU0cf5wIgKwnuziWZ7bDjFcC
bSxxp1rQp+Lvq7/JndjLN+477ExIUQktdELdhb558ze4UD++M3TYl6kMAsnd
h1NDFCQ9Lr5uEOYaOsNFe8uxTXY7y5ZbMu6rHGnRAQq6t4meH6gcCl/DNR7v
y/Tqh3h0N2aK7aeTGSuHAFd7H5r/nlWPxuhbFGjJ0k/LX9xZuq2MZPCfg0HZ
YnkchQkpmLQ9eoV+R6ljXiR5OwkOgU4pC45jWiB2ZWKEu1MqTBw7luy9ZgNk
ZbZvBADR8wiMHO0pFrfkwQmc5He82tAZS4FDSXDER43OjpsEYrFeiQao1L8Q
UN831yEI7f060y8FhAv1WuJ1uj2XU3ago6OfZFlIeeEVNRk8JEwIXCWggqSK
N6puxLoReMlis7CJewYjt/7jcQCQJQiB0KD4vI0kE6H9xAa0KHcblLHceWB4
qi3Yj/tUt6yJ5x90uj6nEssekAEcGL66ZThQ37eXXpDd6jYWRqvmXfTuH5T1
CYor+FSTFpz9kNPZ6rAmAopM0cmhMB0Fe92plyDYqYa6QnFgvguKE5Wdp9mM
CERB5+K/VU1o/NVeciy+E1Meaan10bP8WaWTnTsYNN5Ad6SwAu+s3kRsvUcL
JexEGPLz4OgOqFZzFq7OUsKxUgmXRd5fUxhUHGIRzEHHupA8kCu8uPviVun/
TaiXrtTH+taiqIAU0o31ykg6XH3hdYYiTC6+ROwPFJGAXtQZdGmnc9dB7K4X
HLdYQ0h1rfBLWX3Av4Kf+wom2NZf9VTFikvfzPnpKOAfaSysu8aVbgoprt7x
4K6Ax8kBum9i6dy2AGjoNWUvSU8PSlYECRA+3FRcMOESp3rj76r/ldEY6W0s
HAU7Df43GNfZHEpD6slFFpGSXiPgcyhdeEpA3I+F20L6Y+oS/osww7X3bKHq
nZtdILzhpq0ISOB/qj4+EnFlvoD3iidCuqaQr4GhDf5u7n5d7gB4gyouRznw
mYjYZjjqLgR3ljkvMcd3he40t1gm3ECBYvTNMk2ekPBhNE0M05yseL+iFE+y
95JUUFzeTWQEmlmIHZGG+p6/jfM+CyD3nTVqH8Yv8RuKyW2qn2dANtGYrIC3
SHTX8bMmqHOV6EcJ/EclUIQad3AsFJHA8ljE3YzPKrLSPAonUXe21j+UlpB2
2iOOB39ya3V0dheY0cevGfNOrjmQuajTBP9lI8i10ebqBQYTNSkqJzHzlRgJ
r5OO5dGoc8+t/a1vtFxjuJQkSFXtc5o2kyt0UpikPGQiN6WCMGW2LkjiQi+p
cc0RlPj+7qM8zyRzq8oZX209j/97EAlMqLwYfq+sIYkXO9wJISxnQ5FeHhh6
/bqcbkGpjgRpN1uN35gtfHt730UHScE8uMatkWhHpmmaAtRLDw4bsYWib4LU
x9ZmC7TFVdQXNIuIeJcoZ7cfanWcrbFk6vkkXkVtZAEh07co2NYoQLpGu8r8
/DC9BtDGCVZK18gsMTjtez73fvdbLZSUjFJ5p4DiHhdiacmiVnnaqaUyh6WX
9MfbCdVQ//CCNepL2bInpfP1ICXL/wiptuSaxh8CFIod+THxXCPFlBqC5C+x
+/oANThQnIgEYKgWL0l2nEgxsuu6Lb2swe4pQEvPxh8zV3K3Aesn7z5AJT73
JRVvbEK0JzT9eu/E7I6RB1pj+fPSZ3mw4caNIvV+9DedilbLX5mr59nfGImV
aZEtYIfe6hdQFfqsc6L+n0xiRqPSn3RSXz7S3oKIjE774vagWY8z8k55DE9Q
croIguUU0hVoFoQDGkvcGGGJD3/YQzG0sOHd/yxUVOFXnKROjp3yhLeXWiXC
QBDA0HnezV//PJ7QJ2Gxa5PRm6J9bEBzx/5P4SLXLOkLpBxQSsP58cuSVapF
1dn9QxODImo5lur0U+nIp/m0vst8RlT1S57y9PCUMh955obXiHJCzokhUg2l
WlJO5+IGqGZLXx3Slrpzo1YogIB2tz/9aH/+T4SSp9aYYPhOz+1hvAhCj2rd
ur9/Y6e4KPoin7yuguiTUzzgGeNNWckyTrZE8HAU/D0H+cRJq0W3faUwC+sy
xvmgYFVjmb81Hn2sFPmEoTSXAb4WLjrodVvStRCz/eatUxGsTRW8nJvwEEAn
z6TIEsJIIR4BlNkyMYoMciKtFr9dZKy4fZujvd/pCCdAkiy4yGMJqNx86dyw
1bsYuYLFhZHqmYQSyAcuMAWvFDQAQ08vjEzSgbqk9b7ym93MeNNINJWC3f9u
5maSTZT2cMBvDRKMMqXRoQGAiWaI/PJ6kdoiVedOHxoCw5X4+TZ1ZP9xtG0P
/xAuteTuqBnZDGjWyy0eC5TE1Cpr6j2Wbi757unNOGABZoWYvqBhXVdsL+Aa
LL821OJAtrfdKrHU6SCwrTcs1s/V5WzyG1yst6dex7xEObSROUSRxvzfLmtk
DdlSvNCxU8KKistXD/7NcODrzitcZdpMnjezEC30XXRWch/QHO0v8AVOCTSd
3/LI8D/k5gLi6K1I/2K/M7QElGqyN2xMIyIQjyv5aJ1zrWDih6YER0/x5oae
ED3zQTgZz+cxpz0kYT1YIagybaGFw9n1y9YqKEefstk6QmuvZ/eWNKEoYu2y
4qFVkhiqr0ovl0/mj+bEXmF93Vh8L4dsJn/r9mfUbzGhDV8YhdimRVluuPRl
T7quC1+3oylpksf4apod+x4p6kaDnVaHgKM6VF6ZH5SJQBDi+brOK8xXKc9m
hJDGKqPrzvaCnOHSiYFHatZKlHmWgKbTBZgSoA8ntDDpN34g8GwgUq/EG1D5
Kug45G0uOtxgOWHg0/pul9/HVa41xRVRyu9RVCsQKabuYajwBiLP1F/KFpW7
WCxA8WUqnC8y6WjHKBXv2CcPzbOsxZCHrl2JF2yGox2WKXrfxyKZKKIz3lbd
HPXRmlk9b2nBtfhF+bcSvIJvfdIO1LfnDG+699vtHiMrcCMK2Z1VPZxCMQkq
aN1xMG1tByVVm0oYBtShoFLX+GTCUkO3TkgdfCreEzRxQAPGsmXaT2Tb6C7d
YnDatHjX/FINuEASotVJwc02aejzN1AR6MfnrsnmGRmMnl/HqMx+ybP7AzWa
9Gk41iMmWvfmudXJ3C7YJdkQ6XiK/mFkVksaDypw1WvRZoA/V1zSZKVF4Bb1
66aHUsmUkq/PPmUiOa90AEljyOZdz48C+2MkoJITVd0QRgchtpt/Wvi0z00s
xPYUZ96xL+uhK3X5J3BmUCBJAp7Ax6r3JM7n9akFHPuzm6EPjwA7tw4rZw3J
vT6yGFfe1ad6RIcDGp9Lt5Caek1LtHT1+S+MWSzVRyZqf3Y4kMNDJY1zoVcD
Sekl+aY+OavjioNK6oVr4O4+82UqyaMcZfpeX4rCTQOIgli+dTo9dKQWXf+o
LseqmPTLAGcJa399vSSO6DK1/HYZXbAyg796Hoj9imhJAF8IqY72G+TKJ7PV
S9OWugV6EaK+VSggbcTWAaPm07SLfb/w+g+mWKpnkyj7y7cj66WuiUo1wJYz
bNyIByMU/Cam8XsACgVmeoUcHLd1qhdgI6bpsTV3cGXDeQ1ozVS777rJ90lP
h1NVo9Ffpn8vK/Oa+I6AVbQ1qnaPUSP+V7MeoemyerTODgknz617cY6DCw9J
dr0Z8CTLFFEGXJcrDhwUClBLLaKbmASueDM8xziNuSY1UJUMF5/6xNBgubpa
CnzqostobmaYi6jGbbvnQgxf0MOvfNi2tJfRuE2gMtPfoeKJd/FqYrDEDuh4
1MqC0Chf8e4xBpLoQs7CXObmm8R/+zRsd+AZCC66J8DymeZvRy82na2IkLAl
WAE3r2D1B6NUrsE2cbb/EPip8sRX+rx0UAuFnuBeZXv1GT+aUgogCE0xQCjc
/IZWZDscUFkPsOjw6heIpw9gXNvLD05Amedq2R3W1TOxMHaQmLZ17rwXlX6Z
lQjVPdOCQMRBNIvkRH+woJIK6OjX30RoDz0jbmuc/B44ts5wA49kK927sxTR
T0A/BsUwoye2j2K+F478owN8k3aN51MhsyYQQiWMDF92s2ewg8JJYBkHMfpX
tyG1gymI0z5If7z05dv3ijlVe/Y49xylag38Lo6zmUsKl1YHSStAa7aAh7/m
T0Ckc9dUgvo69OTMqlKRrwFkWcwHM2+E0BSZCMYE9RlnG/RuGLV8vNRoT1b1
kULuxEWMxLiGnuIGW3urL10VLgwmjZIohVxWC3/wo1/0FfmO9qGelP39l2cI
Y38A8odp+utPA/oHDbjM0zbEPaZT4xnQShtt0EHRkqNbbVfkVM9QbEaYGWsw
Z5ne9UJ2ii2tdLUadvZ/LCMspNVx3dpaeYKPYcXbCaltRnOpibT0YwLS3bmo
V0Zk95McrD3fp9xbxV6ywBQZ941DEVT6R0UmSnwaBwl2BvzlOlmmZs1fgJlR
9q4sQ0lU/XDx1VyTqs+1f2y+1n3uPzECCfzGpFikSK483QC9vnAYqzcTDcw0
b6R0YcC5ICADP+pmYXlkvXSK7VJRTpgaGsmLwtzhJA3kn6Ljb76cOZGWGtQr
dy1f7UBiGxDhuJ8LowzMIgjsPLCwJYjblS8Ki8+CzG5FaXH2S1bHLNAL4zvQ
nmWVUZUiVBFFTyWSzwPFF3UiiGVNoaZeecCVg0q+mt5bpGJ1hry2hqefPB87
m5X3XvoZ5ATY5z8Yxq0C6chZGEgAnESFS5kghovxiYbPjTdtNZfb225duA7p
TNeb3pbVgOIXLEE60fiHgaoLsxhYflNa0gJqUGXF7xCgky89+2JHRwzIhHEk
K4HlcH6PIG5ux7HVCZmsqZ1AdxnFQ6KNJc5zx8ADbztXc9p+OdDFFoI/HO6x
+ukT8ZbLdO2ldiXhUX6x7zX1kYuogverngIC2NLT7JKPaYzc40k5DwWq2B7W
EAxeL0gNN75LBBLGHBgNJN/765rAFOfn4LAfIxwyJ0V57r6LVu+1uswG2I23
QQTsWN0FkT3xAkAiLg/3LqcF+U4Gy8Gba//wsmOOXT1B5y2d+oSZl1BM+eUF
504dvCtm3RDRl8+75K6vfdLL5StFQf8letZfzQBSMPRH36lIUoOyAj1xW6q9
JjQyGJjceUdkPjWaONHYAs+jhNWZ/5C7sU94y6FhrmnvCV5nQaQ8y8amUxW7
DI4+RN8EEcYE0zt5IjzQ0zySyeeo0qmfgoxN18WIfwVPugOEXygVI0Fyg+s8
hvuQcY+9UBI01d01DKymsuWOGonkpT2R42nuJ+6pckqkgwjKoUJF5fgpCQbf
pMFPy1Y5aFB3Jqro2ydgD+XqkP5vR2bhSVzQadC+U/Y0dsHBzs2KW1Y3AYet
beX5W2IhJGtfPT8BpYia4+4Oxu0umakKN10wmjSHJ1USgd6nqVtqZTozBIkQ
D1e7+DYW7245KMjsOfmwKOon61LSYbIyxUPyCHOU3u6sfEk/pTPncAiWmqXu
5Dq/ZHOOZ0fPZv5ZUCrV6cEM+M+0KtmksLbYVW8JzmwQLcbt8zn4kE73Nr5t
aFeh0r34rNaIhWskmsMwNpS8sLbc2WrFmL3i7+FeTBz7zbm7B86bfGFXOnjW
B8HL3x7k8kju9l533eI93orRZBfGYY+2mWE3sZL273VBbhcRJqHo754U5FLk
xHPfEVvCM8eukYyqkobdYmbR2CbMAHUf43CR36ED7EZJCBxRBiU0HGLw9iq0
wT7oFL8LaxpjdqQvUYC/gb1ioNIGWWaXs2z8OapVQLYs+4LCgw6OzqmtKDpc
/LNaoBdiMdCNtpiVPfSX+4zAJciF4ePc9Jd0j7wtOPp7p+/VAYVZutMLu5ex
ZPqE/VyqXcI05Owvxgs4jZI9lrjvNXU4uXnfSakCP0q5dMQ3gErYCWJkm3fD
+WFC7WyoTBKtwsmQOYc8JWqdnN5+ATci9CR+vE6holKQU4b7AHFd7nFymyQA
Uh1/p4qT2NxHSqkyDzmqKcliCv47+WEwQYJEm4YonHDgS0ITzoyOGobuUjF/
KaKY59pYyrjFGGGnlwN51+OUNK42Fbhx7mKNZELrcuOmdF45hXC2MUt3rAq/
UrIc5AbXeNS9BLiVRngGAPvZFqJ2OhaS4CrWwThCjhKDcKQU0xK2UB9HaWxA
WGScEXLzZO7fjWItcExeroWv14v41GPS/64rLrUkwQv9MAwllm4W/mzR3GZ4
+C4ckwHM9VdUU/GehejJz/SenbiyeCGJLzphCAAV5SiGOnubI8GneLjTCD3F
NZw493h0m9ScEw8lIcCORdRqtGjKe84VDuOPE4nfWXyqaTlroW41zQXcXodH
ANCKjb1OAdI56n/cOpfE7RdRU/KW/bX1ONY7hY9JR+KfC2WHnC8XBRQTBBIj
7llbtZ0r6GpCGYOcvCEfcTcTe+Pn4DBWTV1swSzvmPPjR/7tT1kBjsx3TxBK
nsbsMn90Q3r/Dz3U4/URMr+qvbyz8IgYpBRqyhi2uhlB6YPGoxLFDHxKYWcR
9CunwWQwtwo8jh+/tnO0GLcU2uzr42ZyOAnMl/YUSWaEdgddCEnCpOerszum
BLuOIy04/JXJ8ZzeSPNEigD2eCViK+HroYSlipglTYRRWBJVCDVna/xarsnz
yFamw6Zx7ndi63btpHKcJCU7AMigJ4UC4cUOZZvv9FsoVQjmfC5JCozJ+fNk
dUXsCYxHaYL+/dTaF5nMwFEnxW581RtbmfqJwF3nfVdX3Iui3ceEX4iDyg3v
fuqbbVmRgDZrXT4/3sijDrYsclaXvCpRZxNVGdApOMSb1i9e5P0aTT27Y3ED
aRt4NmH5v0H1ojKwaAR0Cn/VapiWPivKhLbvUKDpNjvbgsSgbgLU0BK/qhm+
ku0SMrCe2iz6pzKKXrl9V2dBS0lsrlAkwk+gxZiw2ztkvycIMql72TKZAopQ
dQK4FuN2DvaxuF27rEKDE1f1K1ANE/PwO39BFmsWegxrQ8Q5vZhpmeeq5KoV
DOFpugAAy67CHFARpc2kQE6cgtox20jRvrn/K7gn+I73CxNS/CYYOhMBotec
WNj5EvS8ZqElTNCSYkWyeaYIE5ip3W+Mbp97xtmJg8Om4C9ga3GxWb36Xxj8
fx/7NLP5OsRy/m/TE+7IKhEn0oCSdD4W/kf+b1WK/cUmWkwpbYNnz0sTT2L5
s7v9N8LOxPaciITxY46Bmw9U+IAOM0fcpH1WO8aSZIIJEIEfKFK5UKwAQYqu
4j4UzAWFSS6qVb2lz2CDjKoJEFhY7d1v3NAU63PHFDchcgtKgpHFWruxIdqN
m6Of4ZR1s0CduKgNRSj3C8cG027Q8Sn5p+JpNIbiGXA1/Y/9fz+5RTIF9LhI
zRMmojWbNRsstER/pt5aR/vwdauf3j5Onyg0BnU0NvMemM9b+DyJyQRMLuXw
3h5j67HAzd/Wyq2twvG+0CrMPWhzTxLYb5PE4Vaz9pw5BGk4KTT63EhfSidI
AFNbKRrjpK3Uxrj1hOvDsEiKRveFTBOFBMGFIgqOFicGMOYCH5fWKT6gxSRF
O6HClKHJ3cumgw+UHvqfTzZZ84mZlvdkr6KQIk8c5NwevMCSqyJfwPpejYYG
6oa/OOJNGMWOEJH6ZR6EYQc+jqXzzJy88tBKA8MlSrrGeh9KJc9j4Uo24uWa
fi9o/jDHaEF81Yep+6eIxoPe0NuOd3efv81SHMhdDPN+HVD+M2bNPxqMmYJx
fRzjGQfGyt4QmgA73mnwB8k6Xn0rTE2Q7eEPv001mdjVkQDvHEIocOFZV/sh
6z4mRz7YBM4iYrFb2bjBg3FNBZqIoaOeeL9c080pOobWvKJQC6ZLZrHY3Wal
9/82D9HGZKPxTJO34sNz+cmiBcNjxAOPxNS4umbrZVjHzFPC66Paj9mub6ih
uLIfF+eygMJkd81qSeNY2NxJ5zrMuKbEfaBvglZtX/f6GA822Qz+xxTOIN5r
D0dRF8QHVvhTyDUhl4A1Bw3V+uPrHOT8Iw4WCpoEwoFhnXodILKQOgl1b5n6
dc6m5ikpnpat0jEgwtxElh9Fn0f7UyWa9F2rWMgdUOKQ/UcOB3liemYYT5U8
ZkMHeeuB1tKFoBm/gfvMJfeHfL3eFuxv6VUTqKufmZMuPA5+cc131FvyMfmj
OZSP1Juh1t0tPDNPJOtaLlhChbfLtUJhwYyAQaoNNnBlAe7Rs/ldAnDGbtdr
WaLl3yfeCWce7PF6/bvxsfecUlbjKUn1B8DzR5dlKvxu62Qb9Yti5eMbXEJz
piRuUkS6JPtaKMopTS40SS68IxDmv6BicqrYhpuf72jzpYf746mdd/36IggE
tSBDcNC5L4xUEUmsM9llRcbChknBmMaHFU8reGaDvQEZOsLX0dwA//4Lxe0x
DN91i2bSO7T5qgpdx4LzJgDSCoSsF+136lmm5YeUUFVu5A/wjW0OzTnAYItP
IuZGSGHofsO+vpIVf41B3IWwMnn7wdF51fKwzhRgnUU9J+doZsOWtCmoVzZy
B4+QFo7jPHSV5SiLYYbuzNit8sKRrR0bGJfPBS2PQVsvG+aNtnuj7aldM2wF
SodUp6ylbzu6eDI2ok40rgSoY/JlqOpaUEvi0orK1U+D7X/xtB8itENxwtqu
xZF1RFKhrEk2ylc+f/3aRGQevUfxlFc89LHR1ciZwdNeAKYY9pZCO6+RXhll
pvec6T5R/5H2sBblRKDocSCFCOEFoOXXH2ke5mLYVVpBT5e9ZnG9eB/BPjMW
7DJ6NYmkIs0c8kX5O7qYPUabLbLY72bjDznKoTw+2RK/scsnfi/WcbkzJYuo
BpYI/xLtkUf5gM4GYd92udQA/NnuZMaax2bNokODDJtNpLvMY2hZ6oc9TapE
Wdmsn/dZ+9FApLWSm7UeCGV2X4ryaQER+Iq0fL/KgdRuybe7MGMVxmA0WqjD
1E7ne/+CzHM7kRp7nizz1m8PdNhUHQybFZtQ7+dAGhTRtpKnd+Qn/eUZbJkS
qpga4WLuWf5PuZeraMWJ1+ITGplwBiV1QjUU+hzY6AqdJDYW2NG3Ka3RSCDU
w5jEN3tI/MOJEENyJDR6Zd+dYz+DsPHtooop0q9eB1+rAw4BlzrJE+m4o972
tsk/5Qr8mOC0wm1zlq/9pFUDez45rm8HyydOedR1xRp7MOKePRpRMST7p65O
LcpuNKM/+pc66v07qITFrdEZiuEo7kIzV45BfgjnPbPKeCKIPqdviLgoztdE
+9jlaKluNorpL2tLbFWZRAnw8xfR/BiUHXbAX9wT8caMJJc2xxUkvKQtjfOH
8N91pSpDxmM09YH+Dt/9qDFK+EaLqLrD+SzC1Pb29B+j+WjDKNwhXluUDuRL
ysm7KwKMxY/l3+qNkb56GaHX6lJjTWFfKiyjxKSf77voJwVeiewt6W5BU7tE
Jd27odDGNasdmfTkY5YYauqGbQ05OxIWyB40+3y+4k2fesQF/F4V5P5eb0Kz
C4LyRZ2WwrON6er3SeWEF8E4hYxN4dK9Rwwa+AXok77IgrzxFKdav1nevlT4
SkBLA09szJrhm9xetKI/ivssV4WJTOkwxVu9XqKBHoLw4IMMOskdmJNgj4DG
XRORXH6Q4Jv+h8JI2567OJ1yfeum1ZTvRdpBdntUjBtwnR/Dg5ft6AdTUrQt
fYgUgeYnZX+UOPFFmkRWCiY69ml+7brIdk2OUMIbhQzn0UVnrTANv+gsXEYs
rZPaSrpxm671/x1k1aHu7PfqpMEmJm11gwv//Elr+Id161GqniZYbkyfT9RM
FjZubyBrZPSc0u8hwbmIUy7OzCPOP1G1hfUo7Fkmt4brbhlJGCvkwy8KhcRl
Qb6i/vVh8mRAEQn17VKf46CZuQLs+9UecNCkLlD+9KPGZmnvjbpPQj0CXvhe
YBJClN0xUkF3EjE8mg/SDnWc4LIUdf8yqNYacgRhWvQzRlRV3zn4DKHTGTQJ
WQHJyrq4Vfy75lETQXnMaPMP4MJJvgszPXdjbkZIyGHF7v2GgdC6e7QmpFYy
84wj5GKWrLj2/fgXtJNGvGrk9I7NEtD+/S8tSrTtGwKJrKq6QU0eAmU2gZ63
9JqfkCUZhYtESDI2CF7O/mZmihI8FOJor9FRXU63KDYWrOb/6pblF4OpPGBa
01VbreD2LyX98OX0Mi7FYTwq/sAkmFxRAD/W1J4/oBbXUA5ef63KIzbWZlnn
iqJXjsC7SezB+5jR3kDqaLjnZWH/AWOIqjjnx/N2tWB6abjDuQvIlVfuNIeh
Rh75/LNrYS6zRMcY+kj3F1DVDt2YiGK/QU9EJJE19H0gfS+ZQ0rFXgxYHfhh
apxr3PFGs5gHiVjt+yxLhSdFFs6bGjcBe4FvEN2mdl//nRddTDeapfMc0yi0
syraV1+uc9l/55Sq/PXZHx0InoudQdN91gln7THD49qzmFYhwjYSetOYIYgC
MBV5/c64qQHjLAdtmRa9XC5wUHtmTphYGHypsBm1w3PC/Ze52W0WOBw6Ky7w
ln0LyiS82Rf3m1omC5OJmfsRFJAMphyQyNeOFSaXXFS8NbafHGCZxeg1d6Yo
xbTMqCxpm9oJQk7oFUX1KWDdhT203N+IoVHgLd3fpudduxzCfvvINVKoXFzA
Oev/+ZgEVTdsKk9pm7WFD5CmlSH2YNykKrEo5C3HNgusyEbanmSnA/ih1RFF
2unIy3AqmKBCodEGPXQEKFygtqTHOme+8i7TQT65gORu3b7by7j9pbM29Ixa
q/yGG84O9SsWa7f/yJk0fPCAdjb6j0Uh2XCiIuqZbSsE0WiHsjHGz3Ov/WVu
XBcNBchNraXSKqDQzqoOY7AoS1yFMsQCDu/d6+ilQq87rR927jncnZTfuffY
uMx0bgnm4/e+AZ2z0QlmZTIw7wz20dfDxf/yMtr05l1EV+1uaiREcgayCvnc
abWYn1IWgwd7jGoX1xKaZupwSFdas8Kw0j31yR8jeLp/hmquayTyI3plQFXA
bdgIE+SkuDzrPiwqquLaquJKb6e711+uYdRZdm7wzcwKBwgvR69145E0yvpF
SNbbMGMpB1F0dfWBAdTOnL21fvEo4Z58Tx4P9TbmuEUrK+zzfFjy8471flqb
LJxbiYS1yf+NZnIRqBlLrKK9Rujavpyu0bSSfJWx92baFy8rcASSwGz9+svJ
xjeBwbUsw4IqbYdEj08zkvmRZOwbmwciQIX1NHf3l2lMODp/276wxb0jUQgY
Sajr4LOD3xr4j4k9/nEGhMLVrvoDSLF8qN8vLJAh0KDr93hCVZ9RIP1RgDO8
07bv0+02Uao9GXmf/VMX3eC1+LjlpXDteOxbitI+luwLg2fkzy8MR/iJGjvB
sJselrlu+1QqM037BzfMbrpJASnSRCtHdWmcSLxvHc9oftD2+TOfeRmNt6fh
+T69f5vMXvNCGRADi/eoO42AKU+dpQR51SK3JNyS/W5m9x9CzFrBU3PtDA+3
oh3uut81SPrAM3UaRml5DYynvEbpzMQr36ZHGUD6+JBb1R+ShRfLBm0Tw8bG
tx1acswKOFs1gWVim3IFohJUZUNcArFAp+YsQEUEWTiRxQgclj3prpov6obX
SZKrNcYQDMLJ9mf92nPLYRTPJN+Bc3CiJ3rnU54W591DesdLBKtgrTURwuuA
NhGqopZTxor1lxgnrLnOV6UI+vUQHgND6iBwz4WYcKHbtH0PE4e/BzPvlfg9
iYebSdev4mToHEt4MtAjyPeZwd3K/8An92xjSM6+x3qCu13PUcbcCTJCFyiZ
epL2KF2Eurab1ohKFYoQ7cqW1iP29XqCqv/DHRRF/wwaO4jGHmLIAFZWX5ov
JqBq8KYPXqhLCxQhXxfsEagmVh+hsPHu4hmOgXiNcBNUiIHm9HfvwDiLVZtO
Xhi1XMNFuAfUURgtu43ITTIxwSJLwf0eksKHze49+C34oxFzVcOHPQcATwEn
RKRM6Up9ZUFajkxqWgpyMCK5Th64/H74Mfpcoc01u+Kcm7fRemGnu3uLB7Jc
OzHmy47Oi/tk6UvtO6vdz5B4XZGLoF6uNbPZTjEnMRNLZqSf/w/KyDrZWQIb
/Zm0F31xo880qImXYNzOUNYiVh2hYE5orQv5rEfMyk6pn+jNYDmejHljh0Wh
erMkoxL6ghrls3ysYfDJlmJ802K5NV2XUdLIF7L+SlzABtWc65f9yQ4quM8j
Kmxp1Kgky0AYk8RsdvD0mMXTxPGVnHj2mXCqaUCfXI4e7cQLtsfxVg/Tn418
1kGeXudzANv7e4Ij54g18qFhEY4/ECwJ0f365t+iXw6Mc1fXtd3ZbD+gH6ev
BNhRPek9dUTPWnjr1ghul/CkELHDcM5zOpA4BH/izIzB830EMcThUutt5PDd
4ATkGfxLo6VjPfDvMSZnX8bmVZe791MqpIngiILPN5dxRlC7ryfsLKBP8VKE
HzyCXKzMyLd9jvIz+Mc+tU8wncfXlS0wHNM2XNuWAL4jKWFK6p7ejeE/4aly
ijBcN8rZ81GihhfUop/t+a0FdxqB9xea+uWEq5nsH8prvKwO6plzuytR3riQ
YqccV/P+PpuGUf/+iAvJKI0ge7zIFYWL9O6EFoOsxqXFvwZydtjQp0HFuqVd
EtSUMfmxBqrhHySh2YqT9NSQ7avMLM0KhJ6J1MZCJiydwTqlLSAvoZtoQFf7
vDW7q1rYxwnXzyXY0cxCDx+PvrEKcUW2Vh5FwvytI9oewu7jAa0zLHTU2IN5
DYhCoNFCuHOJN9aqTduxN/yQg71PDFaTq6cH+V/8pLsCrlEy9ikuj3nJVP/9
Nvpp4ZM3Y4r9igpGeCCDvxiWOIRqIFuLY1e/+GVnrqbSJ+5shK9mMurNSokB
zySZ2ktzLQc0hc/ZzRVnQsNye2owOM5Mal0o6Oz72yuuV/R6CF7P6N1pqqeV
X6G9b/EXZWHlbltRF7xiD/lMd5lUCZBkusd9CRqh3unXdXyD/kD+XrLgnwkx
IfEgUEA6gKJzmizXeZ4k7PXw7HvPhye+q5nplrFByWHH0BnnuGr2kE1RQRTr
3Vc/1wc0bmpD66G82c3A0dl489w0EoSpEwIc/twDr4zZPi7fWmj7KzpS6H5n
8UwrUqzgBTDzzc2iVj4uKdOXGxtz5oe7W97TDyT/Ivyn0PNG9yMhhzHTe7E8
RHebWfwLKUFP1ThcvMQCtYBywYurG74pM48fpXXY3qwdff2Fys+nncoFF9M1
MuaVBhiOwyPXqiIvgVDmo0en9aXb/ge5MjdmcQ4c79ezCwayBAEfprnqu6gz
1oqHU8Y1n4sYv0vVAVDkaBc1xrldQ3fP3Szbn2NPTMpKWOSGcFGBFY0vKU9L
tMLamCXNxuvdTjrx6Ufrituk2wTYZXVtF7NEvY0txoGrzglYQVzA3ewNHdIP
bB/I19jpxS/2yp9rwUd8yuckoTELXzxe10klx7fqGHRfrQt3tceYffsrJW2X
GpSi66r24kAVApiIJ5YGEwGpr9cuVDMFaM4NXBa1s7kqu6xt45C4aaqIX4KW
mVmrxs/rG0cwamFBldXJGRjRq+eIIUeB2qlMxgEkORVh8NrlomW2BPXy2P6A
oAzV+WnMlQKo1Uvj3stUzoX5T9fU8rBDcXuvHOk4cNn2se7LO2aD5tQ5kuJ+
HzaUX+TMEJiNBlR8eF5MIMXTRu2QFJOJNfkykA8a0GHpyxvjyD2mRUbbkYjM
zhfGbIvcRGO9eZjSLuOpAgJMWfMaeG3Cp4ySSe79xYrkS4AGkugUZbaCsHQm
JbuLTtDS7m94zAi/5OrMa+LW3PInmv4NnsHnO+7oEJKj+j2bPAwkX+znm7Wd
XMvBxIuIrKiB3/voCcjVFzcLa64PFm+FmP+BU3DIN05JBE37Jfr/8zUGa2RH
qHmwR9fC6L5xkxAiUpOzg7uUrTR1dbsmOKWsGQsI35a85nOudfu9QsotAyy1
QYLvEvB7CfJA/LjwHJ71Cvc1SyaZkoiY4w0vy7Uce7EEt1XNpn8PYZ5Vfqi7
lOor0jwlFfLDTT5pZzveWt28Gcr4IE03Ev7it4BmJRtwI/rBKRhdjgWI8juh
9vvi/ZVy0JsE3377MuyPARoOBGG8yPbmR9lAyKGWtqjfDs96DX6ErT7kC8Zq
0W9ZIBs9qTTTs2uPKHatUxbZilY3+SIYlf7XbIs/yOieF/TKZcChiJ4/rZB8
+C4zdMJEWYFvcmqBsvsz/v3/no1hxIqcDZOE1EQwr0CMKt8tU2rscWlyQnFY
G1wN5w0o96ej67NBNqRn0pQoRrVuE+5jwJPma4HNO5W0qHrBdDwuGUXQZTVv
31qqO9wREzhufev2Pur+i9XmH6euLYxHI8vmino8K8L9dKQaBSVEoCZEa2pk
4ZlIs2mWU+ZcywVcS4KszfwP8W5hDhRMdKN/vrS5p/YEBIaxWZNV6ZfRlsyu
x6e92hR28xn+kQ8dhK0pdGJhFj5Rp4MbH/mQT/5VpuHqcKjjRXCzdl87JPlC
IDrYIBSSMevF5WlMMkxsSzTJ2GSIernHm6evxiW3oc3EKBdhleqEiih2B+71
xO5EDOqLIOXp4yMhzKqHVwT7ruVPd8UmWOLBAq8XI9gR6rW6g9JivUhssDq0
oRIjc9L/vJBl3eiPu+PoQtLnaETWgzV2eoZmGLKs4zzclFQUP0d+N6dSywOM
yh+l/s5vLpiVGlnlshUOBI4ruyD/UQWDKRC6F7BXD0rcVu0GYYClMNvqbtLp
X5Esg7AUXxDtiYJzvNWvOhn0AMJ6qNjKz2FSVnkgUQzz8LEtC8CKCrsYXHdf
FfNzF3ZHW+Nr2rC4iBsReT/0qu0/oQiffV5ifwyOjIK44uZlCDZyBE85g75N
p38Xi3R+NcKzz7nR02C3UcouAuclPQeqJOeUokOjG/U0cAb1+VSwRR9fcYpA
Fq4QH2PYcQlYAvuNcv53HwTDEL9JQ5jSNyeqM6YaLSmnNDPiidYqzXnRBtsB
pQQJskUfRUyq5DTX//k10aaqeHU3KT6VAMllJtYtPCrZRfPjZXkI9CSyysKN
wiP36m2DnsuoWLBJ5QG9dd7LLEho/enYIVNN+4VQr/7H/XCWjKz7A8zjMSjP
TwtcHGRI9bFP/R5QLeKjfhutqNpKuonZ66JkPqqlPuiglqtvaB76KgMikQ3t
bx8uhDzv12Slg56ydtl/UD5gU0kFfuAdu440+QjHxC4noG0ml3K/rZNtzmGi
oiUhdJ170s/nK65kkWRWdIE31S4DruNEgWIqG20MObcIYAFLeP4qMzP0fayW
RMM68shim2uGZ3uu/FfoglBp1W7lsPl4KKWf0mqSFXe3TicR7i3KzY4/Onzu
HMKa3m9Exxx28KvypjMafQmSVneD2GVRwQnkjzIorLRe7yDMtsZ1RNpec5nu
JVc4MQVDDPVa7inQ06zUu+wfYY792DilmQXtEw3XU0dRqlL3AjIV+6KVLfzw
/0N33LWuj5qtgCgKn1GjqAilRdughFFWhRfoHULAPZCRLY8L4BjWtVmEfUno
Epba2YZmWZ+JAYFH/ecmZcutj2IbdQkJtDpC2vFJzVLvtXyYbPyxPQcfyfAX
3BiISFm7AFvLqIEXcjbzBcQJbjEt3UqqOJJf0DwsDi1A6KBwZOacmMUNGf+T
YU5+y96G8CUJpB0FJO61vS0tT88552iemTFR+PWKoM21oabrWJCYPfXkpFNf
YWtC5SbgJUi/JqOSmDNLGz47XDVRxmpr+GSedXyr4LCilL1Mbb3N4IRqCAAp
+u/A3k/6n2VqlfgfQoNTmENoJIiLhTsLWxakRmq7H8Y4hCj1nbqA8+GoiNw1
fASZO7hj6mDuYsN1kbrKQLn4fjH1PP9t3P8Mw0JYl4lTxPxgFGRCP4W2+CLe
vbcf8T0fx9rmPL4JwXnwlqgr1pR4oTFCJGu9pEq2l47sq7+12zDAs9+uNZ0T
PsaExjF0qQj2UhS9fcJEULM9zy6kimdmWSPJADu5WkJz8UkauNusoYN/BGkP
VJKkgrWEK1WwWKh15EXzMHHFYNoTHvl/S2x7Fk7pNwI+e5Mp1rvSNK2vxByZ
slC5jFmMuZ29r/erKPIMwjPqBY7hVSy4U9GHvH7ud5mgmhhYmzmz56A7igWX
77X7X/rrXNnrWQFXe9W7/rIRQuB2WVqpE1Scwqi/GtDN01QuZnQxSPLLOLcE
VvrPkSu92wNA5hd0TDM+QqyI8i2OggAysHzNghWQ3vsWGpQ1XzS8owTnyCOv
0HDc2ROjQXJsTCGJVAymjqELF9tOTML6wXKeZ/sgmS9gXRO1bUkGZIBNQh5c
FllcAbemGlRk1Ia6rgMuQSDjHXRozCm7eNjg8Hz1wcsys6+kx6HqwPaBN7/M
FmI5fJsa2T47MYpSY0zePty4aJXAhsgCpAr01sSXCGuLOLqENiriGO3CFCeV
jup+staA3qSIL83lfgbHL/5cUtNCsOTiq1GAYA6PNDbdUilKJ5XHfXk4Qe/Q
uYQlOXpKN5NHegOzX+Or0QH8WjBxsuMxKK6uXTJ6e0Dk+nTC1dsPHYJoL85g
EnTAAwP9u4dqRMRXouf6ACYIkPOFmmhj0mrlMr07FpiTUQbD5WOZGMSFdaNG
u+DomgZjjHBENhfLHfJ+67Svmgt8PpFxSEXpPwZGZrec49u/suS+mfp1Wdgm
0Suyiu9fSeYMGfie0JfHUWDyDEMLeFNAnR9bvcAZRDD8kktgksdLSIccAT0Q
/RoZzqhxnyD+E4mjqXCBZ8iJMQzwMknPRWDuDIV5crg8nwH2NgV5ES3GNfjY
Fa375fMh0bC740qrIxoaNsUQDvM73Q/xUqw/U5IKqMgxU3+xbJG/Zln0+wvb
8ANIdqyRpWWwhnFwbNNDGAn73/oQtwa0dVB4NpfrBai8aPsr8Jz82OX3Smhb
f8H+4VNisp8dgMZind/P+RFJgEe9YBjCFIcGlqq/zMTYQP/H4WNdJYFXTqAs
+lzB04aXxiAm82235Z9v+XLTyVtVTvPUexrmDaGGhxDDd5eWeY7mNAG8rzkR
oG8A4eZZ4eX95vorbOPzP4u49qqTzesIJ4MqHVVpxE5eyJSUFHcuKb0EVMWB
qKXNRcnqbUjvUwcZi+rJCK5zb396iL1NcuWO5kDdehoAVTZIGLawMcgICh9r
URpOzL2xSgdrCROslFulMQIOfMM0IlrGMiah+b3XAwNStRmeLi5MfzNH1tql
YTSCyoPTZ28utPhD8SLr5ukpQmzzG1KcmQHm7RiAUtz9XnUfL8t+ZPtHk2IR
6QkvDPa4uB14jLf/Hzy6OgJsVIeJuQmFEinGQ5rJpQQKyt7EigTY4/bSFgZi
PnGfFBJc9OW5bYjVcDoJ9LcGYcdMzDKhwJpq1/g+8zCBKeO05anvGXarLAHr
l576k/shokx8iKItPRyw2zxhaSlLgCMn1EZ/hZD/jv1vtNOI8fwWpJwfj6bR
NDDaY+86tfrmkVMblKoaLLi7c1XqntfZ0ZTyokv2m5cYM1sfP5ZcSR9Ea8Wg
tFjL89FmLXaoIzGXFRLC3HbzcSnP51Mg+PMadz8QB6JjLUTJrxaSgRYWL67A
IWmLHqoRyVmSMNXy2GXa0Ou2/tMcDZ+5X8klWSDcqKuvUa39U2DoNAUGrkRV
YoniLhr1I96SD1N8IYOnFBLwE5mVlB3e61Ku00TgbCjed0FOKf7BTwrEvsuW
K5nIXGB3KcCX7BI9mw4FREFR6YdZBmVSow54Jplz0JrXQVDxOZXcBxaItgRr
f7v/WErfT5vYX/ndnLrdwZAzF0vNhBSILPuE9FWWaGJubvOzl033+AjN+oZw
NjJJSufrPt6iWy69tv2FufOKzLYJW4WdemYdgagfxVM6c+6kGeApI81fXPR4
syOU6p6NmS0R0trYU5VA0PIcIWSokGnEp6Zh1QHygX8wPOcKByKL6Swqvqqd
kRDKspQlwBYryyyazbyJnXyZFG7gi9HyD64B4qEbZ3OR2ODonrl4YJ5y7xSw
XgTQhckkdmBJelTVNVcD5vdgJTxhodxeXvYrCipENrPmyXTNPeWnduxRWjHq
2o+e+1Dkb9j6cfmbZVTds1GjPbPcHmigWBzg+4TnuN8cJF4xQPndAWemlBu5
+MGV5BUSsourQeYDBIZvfqrotEqg6TrwvqfNSlDOxuAN08BH8OTAAHjPTLfA
Wh0t8pvu3KXEKvmN3CMElUEiguAtlrca0CIeA/KqwbeURY79k7uDWeb8iPsr
mdn6iZGioADgC33/wA6AefGaQSafkfb5hpRn5gf/QeE8EZBFlpwHb+h1Ylu9
GPggADRTWiWbW8ZdnL+s7YLEmiNgV6+N0sBamDE5ldyyQHYuO52GVYRgAEW6
+r6Ci5bZKwLlbR4Ip4Uo0VuGRvtk9kLTjVh4tiIzlrhLXZgudkb5CXNFLdGr
58UvtsnBd/39f7aryEbTs/n3bG+Y0EiaLmABxK4wznwPaF69g2YNpkvjbhGb
sqd/pkW/KKkn68ZnJPWsS751HfMD2Yu7dh09lN7k9xCN7+8AzcdqoZekHWIS
XLyAtO37ETf3PvBkbm7jfY+J7JoU/1rVqDIl99CLagHfMipwQyqsL1+p2mBf
DwA2ZhUtr4KR95Y0wy4OJg7r3gYef2WMNqr76CYjWiW5IAf4B2rpFlyoQtdp
ZzJcBaoF3KXn+wHU7beGWBS3VJKnydxzLIVpBSFSewZHkdLl3vSSTMZ9ELLD
rTP67/eWrsgJskVUzbIG4ONUk20BWhS9vFA/nnh9rdhepoefpN1wkuO8n2G9
mMEHVEc8v6gnNgfoapBn7JdUE2OqkY5uQNMGWlLjnwm+6NIZoOc5amK4s95K
VLEEwDYCKRhqcSoWZaTso7Lm7vJq2f0DcnUvOFLJA10ygZQoqHEfwyaHk6Jv
obCeveClpo2vw1iZTeV6IpIZI/+FV0rPeA+JMKFJ/Grv0Y8Pkcyukj8Mgtrb
D5/uiEURReumEcAL391NbSXXc/YM/wRGjNBbzaOIol/N7eAVAlc3e+RTfHlP
7xIVnlnblBsZxEzf5Q5GseNq0Y9bQPkHG3nu6DeqyqcorrFZFMRT+HX38djh
4MBPyQsYABRoBwDyaXupwM3Jw9ifVcC33BVQzdurEbdbLPUiiGZ4IQmLXpGd
deNHsT8B/Zc6mlgg8GBvnztOCU+IbPqAE0FGOXNG4HnKMe5h1rHeUe+jwD35
I1XXyBjcPyH8v384Vn+tWQ9bG1KyT5HpFTMXe9IcTUNfe6POmC8jJd5Z1zIx
3tPaewg9LAkTfGy3rr4RQk/51Hm509zcZrOUv+FN/O571CV2MdBU9p6+DKCG
bBpPq8fzbWk+pfcGSrqKSsJBUf0ftNAWeL54Tqu+Q80MSCy16w/uS7Kti9hr
6kT+KXi7JxphWKWK2XkXnNTsGTp7vkbEOsWTVlL3DIYyrVc+k4TjaBfXrIqm
DBVwq4GaN0QSsxOZB1hqpBHKA42BB2VzqZTDPV+GZioqtyeo0en5ZaxmJWBw
Rt6vor4NjX8a3Og+CHlzjf8Di4/BbkkvU79YBMB2LJPmf/SKlgOYTHZnpAv7
LxcRuu2rnoGFw0+QlOKtBEWzt8GdwYNrn/Cj3n8k9oxqJBPJ87DoFHgqdpN8
zSYmXhSoVmjX0pndksXWdhKEOmDbwOXv6o7BaiEjoiiaNoykM4wO3K8Zng/U
Yxb+EwfsfHbIed0LdxZBkRiqzPcQORkqFXnkNC+bVU1rfVYmiJObwczsmC6/
dpXy0Rha1LoHocb3smJx2mJcjnUEMNt52XbxfWQykNztdJ4sw0Yw5/wtZoki
8o/Z8vQoiE6vN6Vi02L8MGBNykKt6jWb7Iw3qKoPe1E8YJa/bQrIGcEQ0x43
efCuyxqWkUO06pZmyE46zbkHUaa/7tPWcK2HUPP783VQV7JKD/6AOfwtmq2z
85X91S5NNOeGFd+7x1r3Yeuw7drckRRGanlbFTyB1kJGmsu5eSv3gl5RkXAk
pjVVWOhPVYM2HN44UiyRDmO6mjVU5Ivicxg5FNR7llV0Iwsdcl0ZXF8A9rLi
5guBr+U83IEQV2+ZuZfoRzuSmInE6cSVyBuUTZVhb7m5Y/IgeIg0vP8a9TF8
49pPK1WeoKZuw48H2Nc6tE+KdTvECpV9oOo/MkobRQH6Fp617Pf1pcYFQeiD
I56jfaaagd6jpZb6VjYL04/bYCaP/DrhSoUgOaM7ux6UiBLxKEYSbwukaAIW
zIvQ2uBzGiqX6fuhGL1DHQs9tyZFou1TSwKvI7cV7FgPoApFBgWvnparWch/
vZYnWEeSN54FmXcVwrIzgIFGWsi/zcODDzx2HiflZ9r/+qDDcselLV1Hv4IJ
MCqU5bBtjMElAQbh1MM+edUO7G+/vovOZlJYELBW0lqdcRngmXNIN+tIfJTr
DsWPXAx0N/vymJ3Edw/azAwl+nykF4SOiYI08WEnao3jZWpW8wQzEXRo7IkB
Lgp7fW8qPBwWofrLtyEWrfruqMSiXKeiAvOPXUIqTClv7WzUnFnf2G14W1vw
0WfoKYvF3LdfjINmvz1FI4wi7ij/+15FUiwzlY/mURzhhk5///RQJ9qRYDSP
1wS1bcm0H/HoMt32Y5HBp80pflmjE2nwkWi8EbjsbWJoCV52DV9bZpzgYkLP
oTLRGG1wxKe0AjX4Gmq8za7id6Vbfh+kEVHrLNzGXZ0ezYiBZNpRpFU7FZIU
bfVU5z4dWgOr1d76eqMJxKkcWwMLNtkGQrC1vNXEwqv316BSWJkOnlq064gM
14d3oIBGRoEZwQuC+90jDKvJfFabeOe9GO/3PT9ITqgvlU0jOXgbztzFZ9kh
efg4JWQoOfnFY2hUPIxGLn4KL8Jy273KFsmfU0m8K8FZCjC52FLcGDxXn3ui
NUtoWoj3mIdHjh7bjnb/l3POKpwPHgKadocfyDqSJZFoe3pY+v5e3NavVUyZ
knGRRvbQGkGcsAsr1hvFNl/sJPUE1HRdRNBavRyZlGR/VyXHfugoytegPYwp
VVrbdCf+sk5mNkA5yqLsOEvqwkszNFDjzNg9VykoYYw5Ec32hrM/nhk/hWwt
CoGKw3VvC+RpgUF1qD0cMYaT7318d+0Nw9IgHGSe6NCGpxqq4lGGicLMq4f0
0Uk8SS8f1kfRIQFx+roWQKTYbwzB8gYL5BHQUknLBnNYSZOIMZ5Vo2uw5QWp
Fe174m3wf6+IBbtGfbPvgDOy8iVK8fsO96pB2mM3TH5vjCX/1EKNk/p1m9GN
kA3+l6YJA0sHbPOJ27DkGHgQaxYFW0o1YjV0nM5fsuKgr5DeF7sGjIeHGv3L
hk0+pymMIcU3tmm5/A8na623aCueJniK+QQeObsQi2lzACz+YtWaEIMTSugD
sdqNsO/rXHBJRDncZeyb5GKQmyECyHeFS8lNs5zGeRKYGn37ElirOr70jBvQ
JWRD/jH+tl06vIrwq2o2jhivxTkNzrIaqm+wH2zU9y63e+Qb5RJJ8o/ikRsh
6Sgn+aYXUO8FxncIDUdyEPEEfEqKmX6qQf242ZvQzvZaWdHU86pG8cJfxO5S
qzn1a/Ppn7QCj4FASoAyPqF91lO0mf0IbKvLjdY9T50H8XO96LvkEShg9g4M
eU8IUFc7KmhJuyx/mVO1mvk1txMaMktnFaYE87v3l0e1Se+eGCKPVVwVX42q
V5axKpjDzppeyZPJOgg8R5AJACW0lgT5ehYB/PnRYYB8ertglwkACqHZ1ICc
IIubB/lO63B/GTYVO7mVTTLzUDuHXFyb5iSK7dEUaHgI49XQIX8Q2hXu5JzT
y6MMMoCQG0rPFKbo7WVHrXenxgcW4NrBn29lrichwxBtlds+AGG7Tep4NStK
LOQqCgh9T/2ywc+2lk24G3H8QSTVJ95VA4DWC4z0xi5tlHLUzoIbxRd5AXDB
oBragHLeRtxJPE9GzSIqeH6OFPNhKdcdxd/702U2nIVimS9E4N7EKDF8Kwa1
VopXxuFSKzo7llyUChkpCghfwHC9S98sdogkbnQ2jrE0J7YnKGNylgY2+G8p
PM6HLyaoZNFYIWioL8TEjo7RtM8+Q14MwQ490/dd6wuJzDQqS3nX+z7rXVKY
9EU3dR947htc8edWj0LtYggOAEY55j9eF+iMfdliWsbasCKArImsJwr/NHrq
0hCrN6aGdzmQCbRCBnjmTp97EdW6hJMbLRFEjKcfh5tBapc/ZzGw8DobJO0V
D0m8Kd7YpYxi56RlDmdEmCnBmpkMHJZdSLd35be/8OrIU7cx+rSwO9OsDX0f
31yino9GeUk8prggA0u5ZL4oZGB7p8neuWJ2yaNC3RCGACRoUZaWPKsWJiF6
q/Iu23x0ilTde7jTV/Zbtmu+/R5GL6Y+fNIPhd87U2yfVt8W0kM+n+Rt6Y+X
7AeAvTwh250NH9aVahJG6Fgf52oL+Xrz1hlHoRU0OZhQd9o9aJnAcp298YNl
ZJJBlVElLuFw/UyopJJZcns5zrCmNyyn5ADDNGhoC726WGYBQBR+pRO/bpLt
nXt32HGv8yrGwkwW93EvwXvwk+jYNGBssi+a8wKREBUd+FDuog3/4NkQcxsi
DJjEIeS297fQW2xOTzdhu1bVaG9gFPcaiPME2RkAwaXfbVIx5rzf+t8GGepr
1q1q01XLd/AQ+lseVYE5fuEhkaOr+kxT295qSu2PEDWlIY9PvQ2ezd1k+dn+
rGEapGcmfMAM37S4PXk0+b+phI2kw1ZAa0smydkJBVJiKISVgUOg6L/iTX3w
FSXHMbWXV0RCmLFV74ssdFHPyXYEsVOUh53RinQuZ3DN2KL82gMxEJND12xk
FW2M9nJhqAR1A/doQvNhr9J+PXoZzECE3R6+fOMvxkG1BaGxgBFl6hTs6cmr
kcjrlv4xBBUuwMdBaygEn89+hi34u/DF+hWAEl+HLbveLhJKXsJrO8AzFLzn
Wws8NTSfXgFOdbWVYv22Rc2m0522KL3kHeDzSZfqgVjQ7x/CVp6GHQbgsGfq
zez4meCk1WsAL/u/i5iuxTnCxrFdScNoUzVT2SvWchmmJakEIyHrQAm8lZYw
JifOf887ldkRVKvZWbY6LxFCDX+SejXgdS1lP27EFP1PTizAKwkCJ+l2vj2S
Fbo96f7F9SYWTiut3MzVe81BH3OwV1gubUcFmW+JWY3fO8ML42X2E8x+2Qvc
VOR/Xdz4GVamAxUTjVmY1VgQRF3T360VztpyV79qB12iWxNdgGd2MBvIB39V
keUsaulKzMbxztNbj42QJrhR7k9f8qP/c5b65RCIdzux+uzVkq9EPu48ng4l
hjtbyGzmoosYBofVma2wKCeeu1nihq75XZrtkofseY0kAwOw9vzI6DJ9tJc1
sgmjOHa3OnT1d/hA43K4ss5KBwzAHFcIAoQb1XKQ0AAkonh+nnmWPE40ZMjT
EWjucl4c+2ApdgNDVXikIRrBAfhWSBPcsRqjwfCJML2ZOcv1+nnJSjQzpCvo
R9IrYWOGmAnlnKnI6TMDHeAqgk/GFmdPgCj/04j9cPpq//q33zxpGK1EXhu/
3tI5KEmmHOdH4N+4ZNDcGZjEM2dlXLEvrv4TI7sg+VRdGgEGHy7TkOTuJL+c
fJO0JsDUMA5vDIcjoxzy6b01+XAWaQ30CgrsMLSXa9ZTy8gqtShPzga529k1
hO8dOVgLCG1nFqrOhISjuMl5nmIAojJSS4Kz/Y7zWLTw914YW319yTlH34F6
VX1ypr36Wm2E4jqtidBQs2FNVE5CKH4qemF45UPPh3Rkh8JW8gP28mMHdxFY
VzWQYI2dM7CiMbS2jqeS0n0nCR6RMIResFxQKolVZEzDO5tp8pNkZWBHPlRA
BGWWA53057co61TJzuJUoBj+MazD60dOZWb004ebm2TbETtlLCWy4soDgLDY
LMVezRN43B88XmL9sEVbtQZdanNzdMkqyvtyCF5bRRYtzzFRe0/0Ykp3e9/z
ELHTQOD/TjC+e1trGBwGGNhuNTVOuEBnIXK4bxuIumxNmyvBybUgg+Pz2kvX
QUh8LRTrNsPoaRQTgCQA57+ieUXvtZKBvNXSsUgnGYe7a9XjTGH4r5suoeMN
07+DZEESu31jZSn9blM6VqNbUEjWSNcQzSF+DVqOauhr1E4coyNDa9MbiDY2
+zovc2qK+XhPCthDeGjx7lc4yffTQo1aqvjmOkVoEdAJzzlv5LnB3FaEBMwZ
+HbMpeEBTAkcpgHQFwuNYxsg4nQbcrsVHOeaKcPinkkna3mLX/gjUoyYdaLj
rWpF28Iw7QuXC1KS+j9T5OylqVuTs6YoOJ9pFgmjyCiFXgoYsZWRUUdfSlrZ
GH2MYjv/oWEiofoKvXJhQh08h11iDulOyV8lZ/KUpQf/zquN0Dtxna1y4IeU
796qJ5VW7cN0JVLCsDmMjwskydhVNmmAotAP78bXsIwB/OjgHmEiSeeT6AD1
cQEfyg42mJ0Ba965kU0aU0BprD+oDH3fmmrtazZxML2/ppRdPCQIUf26+B14
0jblqd3N0HBwg/SJB6Z4GRydIx3EYTJY+qcpmJOGGtrlvtg48TV+jdEwzBBb
I31n15yQ+qngFKWBibWwjykBmYNvRD5exWcdefDscEP+Q+EZt4jEu+2e4/Up
QHuMDR3Y130fO6lkYR9ge+Qp2rqfuTKgiptSFC2jrgmz29i2gso5yp+de7/d
jZgpF3JmDxOp+PAZZjEKZfYhrYxtvqKZef0cE5r4Jq4/7LIIBEKtiFekrflx
F1o3GKwb6mw1drHz/Z0TJs4d2Cs4wp3zkfvDnBimpSKJeZMcuLSfJ8CncPj6
84H2kDxCfB0noUoO9c5nnZILSPkIR7/3RthxZ1NKdY84JD4BDi44nELw79eA
3PBOkl7vlQkTI9QeMa9PhwnADqA+X1FzSL16n6qM2FoKpTKL6zCJRYfyqLK4
+Mkdyclh6euLwwatDAazhPVoeF3NL84Csx5N0gcoC33WqH6nroAcbuR1T/A9
MRU1U/PwYvPDLw1X3MgbMLQKQojIiprRiUrZrttr3lmcxdmxdg43Jy92aB97
kMw7U6PVuiMI90bANLt+nYQNqGYDTohcTztQCmvcqWaYAUg/VtR4X97nJbn7
neuwP6a/DooP/AHCKwaM6GkIQJHkcGJw+gQ72VsAlo1OtNbVA76aEo5CWMR4
x6lS59U52VhyUzbptV6g5nLZtPV64WsNvKF80aLaMfXai38qKuG1l98fyOM6
eyxZtSEi747FPHh82r6P7kjJiY2p6UcYsDxFEzfg0Dd/D5HgH2DDDW7PSv4n
ZCcmbAJ5um46ySl30KGRkP1kdZOXrNVFbn8ppvtS+Iy0VgykikBbujMZV7dZ
VGXc1Ul19LjRrda8GXO8kNeGfiJGGuEcV03OBhvSukf9cfNxaTwfp/jKYj3/
ga5qdBI92mH/gDn0wut8zMz1qWje/s4SvooWbRAqrXqXJcBkS8EQoIrcou9e
kDxbljr1rVJzArWPv6oHvGJVRLqKV7eVBHfVdLjD0Dkh0iBT/zkqH4sU0SO5
O8hOQMpICDnb0HGHkNJiQQAho0UcwO76DJTNLTTPTaihOlJW7Hj5YRl4/WLw
B6cb2S1obdybFzZCgpm50jc19QvRiiSQUXBbwhlMrqfdS36yLjHjfIJvRNmu
IYAOwhdWTiM1VPloGEawxU/80kz7o1mKRrlrZ8GBtLqmf+chmFyMKAlTV37E
bxc3FxJxR4dO/fZs9rIRCbS+GOomvibZFEHsC3l2q0N5y9zLDdGBU1I2DCiN
63hF1cqkjX7x4lgBIBXqJLwQmvvylwGH0g1E7dCN76rMXWZ9/qVf6q99wz0B
sHdHGBJzGiLNQ/+0Jl8xFv6QKlKLHe5MvkUvX3+Yp8P3iiQE4BUG6WEqdheI
gYAAM1X1j8EtQ1P5t1Gpp9Cjr4YUrVhiJjc9Ip/okEtGqVVDlmeG1xF42fAc
qjMsUxChPQ9hf8QoUDnc2mIMxNmvIIualf+z3Yby7vYBtt1/yJp/cFbETOdD
AeQnObYKQYvKE6K9SJPLpsb4scnnhoAuf6kBD3kjBeylMXbVgeoEPzK8Fnjy
+Hn7fqe9AryUbd28WTHROqwwQgN7acLUsQzQmT8QsBlEfmAhcQhcgY091l5x
y6my6MFAnzhLm0WzwPVcFiGfzZxuaorcuW2jqBssNao4YHKg+GGBdlYtOY5D
ZKabwNS2FAAPoWWCMN7t1FYLtEW8bF6z/nGtYiWiQNTe1HUfw74KJu30T3or
72SCJKMvw/yiChTDl9MRbLQv+3dvmxhtkV8aTEDTl0EpdF5vKZjysynVd5l5
PafSB4id6YmWmM2H1uH5T4KV7fnI2YtFwyy+XNKfXPaDWQ7S8EYGmHSsypf4
JQloNP44CLyAK+pvqzX+aiFtBWsuAAGXIqleX2FD6V5vda+KAQCQn2X9hXar
uOaN2ATyE6zkXLvzt171xgvZJGw+5kgquxWUz1093ccrwsqtiBsnY2PP6vvs
e2Dbov+7vN5Yh4aK+ZqVf3gGgzQRpKcN2ErIGsDiaYgthxHauv1BwmvdicSe
cD4W11hth0baGGosj9Nvo5hZqB6UmkFFmWHRTJi/WHz+t2T92dPz0NWb4L4P
HFRZAe8c8KIDvi+BpW1MbXIkRkhAEtlpTViBIsBLdMBvPxZKYp5h6kLvTduX
LDqw16RlcMAnl7ah9VLsd+NjCet/ecgpDSanmK55OlbWzpWsEcQ3MmGoJ/9z
5FYubgWMqGBxaOjIb6Go7KF1xq41WcW0bBY1iiDQRlmd+QgQtbJEGLoGhC6W
xfgnZ/5ZtlBU7Pimw/E0RFe3nY7S7r9MNZpwGDgurPTAtzFsWbGTKhWk6gc7
zBHNmqLQh4MC7nIzY4yC6S8RupEPwLYZqNnBMNEJOR2qJSzz+aZOuwL8nERZ
FXO+FC1Uk+xHvZIiD2VsV9uOfLANPRV3liCF/4qXgxqvZGTOG+K6gfC18XLF
NXkhcLAtMaTvsuK6NzpV9xwT52VCtw3UkD5AH9yh5YwiQz/zFpHJlYk/UQy0
U0lvosQXR8/BoQtFWzixAGUCETnnLZdoWnl6L0PRHGSPYjUzTvzqUuLqW4su
bLV91msq9ppWUKOgBVicA2vtDHP+z93DHTzUs9J0octIoZZUDq+hvgrqFmYU
5mAVFUqV0aWWjXFtjaAYNtiYLlQTlwICfCswnvvSwDpU+FtSeMYNnN74tqaw
S1nb+z5YfqdxYfMfK4QJOlOGD3pb+hLDwvmr20HXXXmoXFeRQ/9elDfK0GFE
epXCa9lzMB+p4eijKZjWmrU/GcctS6uIFGVyQb7R/xFg9elvi2HKn61wysCX
zsJnbQKtmEZ7+CFdGL9gILituJiw25b98n/apYox0vueFATNva0adLwqq562
i8QBOY5iSW335x9B+4so2DGVs/NiIpe/cCc3BB1zbl2AqQXm1NPxwL+ofGCx
Z1dHYHJUrbTTXSUOU87P/As3ioi0B154FcePktX3OUG3xMHgbZ1FjIwJlsSW
uQzAUDidy2sTurpei1yvMSCorWHiADTxSdGR1nmVdcA4l5XZdqoyQfmts624
atFwi0kGE9f6B+qVTT0da7GJD4DCqNEuIa6DMjsKzGpky05cmjzK98yQxKhP
EqTmPSwe2ezwM2IILg7vsMcj0fMmnzulJqCFgNaFbedZ4wa4K+jye0T7PaBW
szmjluVlNVwuvnSJ25jrVycNIhjY4zJsNwFKfBikXEkMtodbYZ7gHSl5+JV9
cdjDzLHIdzqD7VfpwrCjDmkMQQfGHLgE5dCjmtE0JZjkvYPHtaGuxlE5kN4r
J6sSMMS7FCTAqPbQ9H27Li7X1d150S12aLfWI+79wubBSDgt6dU5Oh6Gnq5h
mchHb2HGXSfsmN+Pn5/tZeIQX9zl2k04GoN9TRnZgweudTObxX2b42VDmPe7
FrPFJbJYwqljwNQTvE6o6px2tZbGdGbac2qXr+yG+rLWH6Pg72WYUoKMKouS
BfE0WxH4iwyZUUJDwPpoY8K57ywHnoITSrCGszqVk9ndGFwxM7ntCJnqqCm9
cnqICZjtHaQGzGFQMEX1Cd33L3E7SZEzUgk6mFzhomJlXYq8HR6/MJXBeX2D
13UNvHOL2ebaImIoxBh004yOjjU4JnGgBeSn8WEQc+W2Fs+wXP/AEgHgYGHc
nFvm8go639elj6OnxDqkYwO4V9DTIXrhY7+FNHJU9fzban4cD0LeR5ubb/Uy
km7/BJudjD67+jMIG8md+k/V+gVmB3WYDn6xfM++9ObzkUqpShbOxhUsc7Zt
a/tkZTtrShgDajSuJNEBX3HoA0tgERzKqTjtRKXurfAsTq7hr5IJGuFrk058
xE9mEddtz1lk1v4Ts6dmU3Yl7fPdYG0MrhL8I/w+NCYbNDBlnH7pMGsf00hk
0wk7P+Mr1c6PwGHsZ5usYYfGQyiSZB6HDEjmlqPtUZ5wIJLw+waJ1RkYeK61
Dlcry3DkOlhDa1gHM38QO0q02+bN+L+GNgvXY5ELK+cgDnekhPjayKNsPJ0y
KXc/lL2JDUDS8uXv/6dmVgWcZ5Bz2N631TSzjfoRvGGB3LvmF9yXWN6bv6rs
41CbMtpLjWn9E8Vj89eoNl7Sj8VRoRePcJV3dve6IH7S4x7MR4RLJ9TlmFDt
ExTf1wYNz8m00ORV6++OzIG2nq5xfOXrZpw79+HSkzfL2yOa3wJSnVtaO00q
6sXr6DXVoVKcVwy2Lsm8WagbcHigfNRM1h4EKG8DqqpUF5zui0yZVzYDZbj9
RWt+g2TTORHI9LgvCalWv93UfZlhzzLgVpJedOoRdGdLmbw591K80QQl+gJf
9oO5Z5qJDxPfCNZzDhPGgxvLYIRTyBmkNHyBysJrymgHsZzRrMYFlKvfJBml
zTHaVI9HySobcep8fjvXCBj+jF2Z53YR6Pd1lRuIan0oJ5HjvPiSZ+uOlw7w
V0fn1zMDaqlFUAnYNmrQ7x89msXBn88wUiCyU1AIRUmDKXCZy2b3LDPdHXUS
66MZPICCr+WBYYztrp91BmNCXg8NLPH+iltrd1yScYc6bDcQAEk1tSayXJgG
0n/27HzsxMOian769wlniBwSSnfI0F6llmiNlavf4h6l9N/0osvh+lR5KdEY
Xm7Dv7/lgN7M0t6WwdKNeofMhNnQS9GkuBsVz6685zG0z/vIT40uhQzuizmC
ZHYftkHuIGJYwoPVD5HdTF+e5hpuvZ+kpJWpbBgYXgLM7ryMdzAfessSHzLk
5QVhmX/VAAZ1a8lRz5lsrpTLRnmNImn3wYQQJlp2zUF5j0lphw8F/SLk5AXy
HyP4ev2Tvr5kG61LRCgStMvrUvuBt+53RBFPPQdb/YBRrm1IoNtSqQjdlDwv
mfQOG/Juo6CA3rN1KAs9RMQKcMX6YDjmyfOIGkkRAm9r2ZNQDfpW8AUItcE6
1YhV+l2s6mKhklZSbw3MS0LqtT/gxtE+0mXDsEvXAb2L4Wxx+Ub89p9iuxT3
ZI9jMBAnQOXRnnqmBjEclQcagK1ukl1IX60+NxXSbDgMMxCswaa/5Z6Ocv1g
rRe0jdf4a5X+c9zjwyhtWr9h4IBB/avMoV186QeCn7oz6lEziLznXJuf5sxP
btv4oFU5cxWGEfw5DAgh679AxlrftDphBE0xx9zEkjKVAEBPy/gTBw24r8vD
juavT/PJLWD1kIsZfchRJAJr7ea9JXEj3/ukALbu7Ifpiu+NcMZytIuWYfSF
1lkvDEYzC/enp2ugHi3KeDztCADiiJb7Vxa8hOJJ7gosdluZXPmW8X1cyBat
/c5RF/PQRv/9l1inVAfsfuN/jelRHVCdHCeE5ATEGzP9mcRLLqZMgeb4X0nM
FIi9636yK/fyOK11PooBCANMzZ/SQ7nkPic6hHtawwme5Zx878ZO71zi8gcv
HoU2pFknI3R4E2EJc992utegbe+yfRlHtV0xyXNXKSmGreYMOlZj/k4o9S1z
LMeGt8dhxVCflF9/PNQAqUx8srcYhUthhp3aihjZYZQet90iqBY6Xk3gMPpU
ZhMinSecH8BXrNQQ45Kw3KkXVrsxoUuiWnUBSp8NryopivPK/L+OAIowQncc
6sMSDa1yfZTsH8X9JiDImgELufNu2jUReE/kS1DeJ0UQlqs3D3hTlKhowRz6
s8NFkBCA0c0BmGP7PlBfcDf1VYjukZ36ZxtsXvJQ4U4GbDHNXkQoVWhFAOem
Wuo/axnprsnEY0DE6UR4m/2v5TfZIOSL1gSUvGnjBKPvqnIpaWWRmPEyQAQL
X/zdkjDCTmufyk3K+tGg9knvanSVY6qGPa7tJHzybYmtaNlKXqRwVAqy/VG2
/0C3iI2VFT6bNvI1NMXoG9btE9Hw5OrAZp7fGMgWj8UsLSAoTqervbfSqoir
sxsoOSHdy3bffqqGkmeuzq16CsLtkJ0cjYRxGA6Nur80vyc4h9RrMgmCmXLT
+DC1F1QAS4foHHWtoehj+8nUYy+lTvpY4CtgoMGYjJm0oBEuh44ua8TnjTqi
7u/+uvqPPdQ+EHGZtxJH5mNkYwhXDJQgsa5Gb1d99bvgnksw57cB/H+hPfFj
A8kL3EawPIhyAJpE1LweFnWKTTsC26Cprs0OtM4PuDKbXk8yiQaF7yVnAPaZ
YcFnrh8Rcq5OPK2ZrvnhNN68f+Uwhqrea/NEOMh76NWcQFURv4Jsjw3NYnnK
z3i95tjiqGa25biHPTKVqUXvlOj46GuSw7TC9wW4/GLqsdNSDgn/lPxX6O5Y
rf2hruXkdf0DlcDR5jIfS7Pz58VuxWOFbcEaaZyi+Lo8GHkLdMTdrDFqfrEo
UHw5s1kwKtK/Sv5nJfiTn/k+YNh0CBYxR4JTbZf/oZRZ7G9UQX8Rvug4Uugo
BbOrL+vdq915bKeneLbNtEcY7GICyOlf15Xxzx88YwYqQ9M808/ZvoFBIFke
CzeOqsg3WOP8OVNS3LMMcII9ftWGNgJiLC9NhZSUrNLbyb8Hmk4YotsviBfg
1PhjyhFB7+X2bESLhfaFnA+R6GZiE83ldMfH5HtpulOIAAubaiez2+rsNX+9
Br/NEjrMHhwmhuGGePNFH5vLuPC6QBswpmU5m1hmiIRwoYhYy4xCEFVXIR3b
ulr61v6MHdBfLiPHDlVYkqF8enfvBq/QGYBxYS2vsq/D1c+I+nkP60lLCkdR
SdDaxrNEUMyODgTs3K8QsBTflguLllmz4l0W8oxnhDX8CYe3vqprEJIHFiXF
U5S2bXVR2M8Vx14HZi8LKMNG7OIEExHjYugu5UeVevL7LcN1sj8hFhRTyLL1
O4pKHuN9fT5pss5KhHKHI5IHDwdmts8yTQmiePs6C8KXh6VAs+8EdsNce/gW
gGZfPQfFza7r4yoXZ9Qvyqwh5E8fchYut5Y9UnzEGf08sChAvgjKei0460ah
Z8EInZziOcE7hIshB3OjSi8rQHRSuvInBQY5lSuo39G5vrEoRsAfxj+fBVbR
LQFXB15BgqSGunw4UvDjWmwhaRiK3h4Y+HdNJ0fRPNNE0nmxWU/w8w/pWTtS
kqF2lcy3D4r+d6NzOpEMfwqGTtwdGmShiQeWA3H/zx5ZPj8qmx6zVJHHeoTk
UwNShfJHajR+zUX22b9SR7WJXsZHrEI4YloM1I8Cs1FGMGuD+EMBQeRN+G+b
TMumNOptKHplak/KHV4A4H0pIrzzth7XPYW1FYTXOfNP3+t3Myeduu8rnNBV
fLPQwEQptFtnCKPZFzOTOwts4lhetubM6yB9UH5z1svGwzm0A+O3ZtSs2ocn
eW/+/ejHhg//3RVUybKZkc2TmdhwEIjbIMCEKByU9NGVPhQNRju3nkH9+Kkh
rH2J6aXknYGHoRqEg7omOrmjB2un9yfnx4qwQPYaOOZxPySgz5R58pF9XZHU
3o3Qm5ZiZfAuxhRzsQY/AjOFTZQfnWNIveypWO/r1QCyLiTN0Vqn/qiT9YJS
KSVGB0h+qmLqn8priq12m4FWn8B4oNCjC11g2ZBzmssC+AIBp+WDoSlvegi6
ukaaOMpgOrgK81XIYt/hkwaoRQJBdzUgCPM+N/Ykd3UlU+0ZWbdZfQ1NqhED
qT8wnGObJJ01Jy0pptCWFfIT05mlSonRryiUEHWNff6CQlQSlzZix3tDoA3E
6UBFRNfMmgS3KJu1EeGbW4XUVtoa5W8xy+pzvMNwy4ERhlu9RhaRP7obT7fg
IhWsIPsHtb3KR0wUeh3PjzC96cmH3ErL7b7OITCNwP3tu6mXyd+Yj5PTrMUB
1bf54pTLDtSyJ/C0xsllxbuWYarDJ105QLRnaz0LSjBEPqFHGsZfK1mc2NnQ
V9uJzKdQUj83/ZXuYD5zKAWxGWM9I9/bkG357h6aTCuPW0RngYZ2do1/PDos
p4OeWljsv2blX4IW4DiNZtbpSjBV5hQ0odc6XrSBXP/8dRRWDPv+/WWUOcoR
hKzl4xESqXVFaALGy0XMp7m128tTmwkjmyFY7uOHzQblyRuPXT4DYJUtutPp
dmkqYTmvijOxgFj/i8IaHQiyWH+GNf6EChO8ec8hhQwTUe72I7FBjKqljuDU
AgFugBSXGA32AWmRMR12g75A8cO+a/a3K6Pf5kan6ORfVS6okhYVlN0fdy49
4ZgKce6njKZ9mjB+NDUvO9ryThmZGFWoZe1AD3uafatRkNbIuLQ1ZqpJY1AW
TwpLXgbbKK0+ovrR9/ezvBfDqQC3dsntLrwc3QadIUURY1tBYdFP7SxxKaJP
3mrfPzkEXGVnmmU5tCBGXtfrheTTBKDe0fSOFbCIUY42B74whxvoOk8H8E3v
Kf6rs8+7p3O+vwPylrPoHUy2QI8GTCfFexPhvCVdS/P5keMQzjqhkZ7LOYJA
snL/9PVWEJ756iTrq1dk+ogtznIRGU4mE8cmUFlQJnatlONuiG0eBHSKAup9
kafqHZUeE5SkW9VLexSqtHuhT8z1S0Xfpanl3ewqhrw2w/5ixP0LowsFZ4Mq
3ly+Q6ra28cZXciUw0cMoUuHRHft+1kikqI0AW6UDK8DII2mEVhHlVgzSdwG
0y2YjB2IighKtXOAqTS0nCXiVA9VNEkjuagV8j4/a2NHLzCtOqv0M7LnEERs
A4FSlZ0jtadGEfVUfIzajzqClVR4lwUe8vnGsKRdlSGKU4BTkgl9LbfXtVbv
yUeAxTPasVoQsTm8Abuxi16qf3fYo7MI1mmltlmKqjVBQZtJyOdYhZSd0jfR
iIDz5u22gW05QJ+dbp8LyPNkaRODjbShX3+zcFVEQs5U7yASy6pLAwFWepTz
huCeBkNsUYLLdoGjtMJ6W+QPCgHORAk/izfNoxbB9C0ulxAfqv+KX/e8M6wG
h2GFy3LHC7wR16Rm0PcWUgyIJc4jpM4F3C9O2IuT7apfmob7HceRQSCHVYZt
ukjhy+a2xjLHRSFJyYdqFnyvA3OVtvQRTseozmTcbp56SlZKcTSfsPbBxmsd
BgfPVbZf58wZP8LeHm32gsOWhuI/eLoPsdMIL6+z/10u3184X0nEMHyOaKLl
wxSHBhTXn0g/ma7XuD9r+iV5YZHd4jog63U36eV1lpr4J5a9MtXbr2gnvJB9
oSYGkrt4+g6UczIT6mIroMvU69glB8eo8RU7uy7yYREsxwP9m5JrLIrklpGB
m7TZMmAp3QYEHuVc4/KFxvzOy4M6szwA27iSguvl4eSazDlNzQNGGZPnmObU
GJ4wgxhRgsYfGj1nC1Y7mBGKdHIqmrYza301oDV9MX57+2FHAU8CEhBkAsUE
7msVPtg9SG71Yv/+2PrfZzog//XX1CLELIOTMqpaVoKKm7noG92KhVvHVnI5
fjmgcjMvSafeJUDVe+kH5ZRVbjKULaPdMAOwVz+iYNlZM8I5vFPTFEf7qDNt
uS0qCwq8jxoG4y9lK4JI0luY2dDR7m1nJnlj72fNLH2DfuZWL6ZjUNST/wW0
K3mANeWVIZCPYsuPauqgPMoA/rcjRXYUNv0XpO7NHvTS5zkkaYnuiqluZybK
Pk/UCprP3Z+K7Nyw824wfK+fttQ3vRjrRTAhI3p/VBI2FDgUNI8/7hHtb2ZU
EQCS/AVW2JZtHKVjaHL3dNdZfOhNk6Ty28JnF5CxjlNisdtQl/LvRnIVvmbE
HaWUuU2EES0DJw/V5dMXGGwtLAGCwPvk8uqbN6ORjZBtEVx6DWQ6jG4WgQ2m
6ivgsmRNCSrvD9uejKCpG5CG0hZinvSos+kHGOeADNdiUBy/Z+IDQCvSevtq
nrzVSAERGIMwq38M6GCUyPYgkF+NPuZC7WtdkWMSCAINVXc0KADmFWs2d9KF
5IriRFxsXo49hxYqwI2463ccfKp2JJoDY79EyyPAlQykOKKgQ22ij2rBNf1d
Q1zdQiepJDxrwtIMGUvq1wLqUztIrIpNkAAfSDZd8K91SLTxXzRIs6v8jSsY
xF1w7C2C8FnN5X6K9xgVwQAkijViHLvaJYw+kZDamuuPJiHx/Pb05X4t66ib
GFSGf8Yh4iHxkcCVJWIH8ubOZ4pcM8WsykOS8zRKN8/7J+bb8mb8v/eX8VPW
lNgzUf/etG3zD6K9xW4CyFiugBphjNVDr1S9OTl4WUqPm5iBXQdKMQ4s7cE2
fmaWu+/NCka/FRSh/PxQhJj0abaA7yAqFoUCYI8k/ARjB3gGQUDd6T+f1rcF
H5/zvm6GWP8HcJMz1ERPByftab9tOZRvEHYmqfQmm+rYX+vIKVtWCl1DXysh
Vqa4JFX2uXCZxsiE2YS6OpClTr1RqMddKWgTmGlszddVQilCWsmHdtWF3bS9
psUgOjObbYW2Yn0wwTfT0YaAQlxOYolzq2Bu2ctp7jBye4G7cE8vG/oOfbpm
bbPUDf9W2lT2vwcr3xdh0b4uBMHBNCoN7xxigvK2IvUkdgZQxuT4DL0JBRed
IYiqZjMCtsjarofKghdgOEEciQ1/5uaMraH8LPkYW5fOoQ+DmyQ9IGJDZXAy
ncW7eJzye1ULYmJWOwRe1LchqjhcfP4ByiFrAVv6QWz4KNMoWx99GOWRdKEc
Uoxc/YrbWNY1UChCweIGqJ+rubTt95peR3vUDHmdkZus3sS2pJbRajntqXc6
tmeXEa5190Hx2Y40WveI/nEEGIDUqovnb75p+YohZEr7CnOYrpx1FochbO90
bG1Zx22KduFyWUBVQiBPXvp119do+Y9quzl24yEQPH/k1MCPtxcWZ6INPsEn
4k5VcRF0N48ZJ0PfWvkWXeMeZnx9rdc5GO8X9q+xHEP021WyfGsChfIDZ+Nq
MNlUF7heqa5O8QH2vHe3TEow8wmR/7R0Y1fWVlG6W96l8pEYssXzT3hWFo4Z
Dc0D3D67ZzYrLT5agkCRX5YnIt2sP4WohIwO/NZb9V+gn8od9KIFYVQVVZeA
e5g+WCvpK2un96MRu5Ay2raC1iqsM5ZnpizT3a2JdzTyLDGq2USapWGCigeC
DJO0oBOFQsoX4unI9ef38di97PQ08OuqRjoJZXz19vlWEkAuG8K1XSMWjstx
Ol9D8yslgkKVlsAeL9MA5Y8YXQfs2GjEx4ZpjuPpWuLgqetloNNoX1ZKcgYd
XGnbGiv97ei3uHHQaakTU7q3QKgVq3nHT0zYIecfI4D9jUalkWndP10OF5kR
m2SFA1PY+jzSer5V0FUbJcZ+mprZ2F0ZfXhxL68ZcKlBpUZ8UCbqvgGgEQGC
JsFNlVCP5aVrj5avP3L9RU9YaQ3DsjicRPiQ8AdkBFuH4keUMurEh7ecjkDO
5la4CyInwn9jdLuS2juIBYyrqrzHWqd8BsUZ8KLcC3MNqAUVtmfaiN+NASXw
IgcdMDvtjklEIu+gnOSCDkOa11daXZp8/WNFlKfmpJ5826319682Mm3w1kWm
kq5fxb3E3Qek9FhzJYVKQLvQaxw0jUgNZGeNkTVZJguSxcJiufnN/e8XEc+i
ZPyHpkEGkOEp1iKum1ZxsjMWVSrozeKTdQjnEXLHqqnm+Ve05N7Dgpb9zZL+
DDRvHGnrEmWMaJxCQlSp/Gnz/IOiH2ION4UfjVosKEo7F5MorS1BS1UkL7eu
aRBIVZw7V2V3wzMnW2y7CNVmOBNOTbpxfCEOWjYY8OCj1jDT2JGAtAC+adpK
Z9II+6nU5ryT3d1bJa4C4Nj+0M2Ucpvf8rF+hAYFCpCCjdJpIALwflA2I1sJ
8YvXM14GAsMssVhM/eTJXhEZ0HXf0i+z5Xv7nS6kGi+Tt+8+S4yC+PtS7Srd
gW7ijq5R5rJNUSuvKt/7kiTV7sxymupryKVa6/jwQoiW138SKZn1sEwho+rc
U+oNH5c23af33xGCzj8wW2MD3VEtiVlYS/kQfuHZqKiYea1/OJFDh8UGlYTN
4xdh6E0g3M1bu//4q/DCOZsx9nmJpKXI1902bnY4uCdbxGkZ1Nl/GtW7k34T
ejBP8yOK9sFGNV3d5gZJQgzav0h8O4yaNJLaWvf7LrIKu7ozsl9XVv/Cooq/
rlg8vdIqVShrV9Klkf46YKM6B8t0EHCkq7AcTD5g+65AlHvfCgEG/LBOUB9W
A0AiolN9qmST9GJ0jquhz60a3ik4EaMhXefym8qdiU0bFeUXssaweFmXwkR1
ZfiFZdgFjeVd1JOEsDK7kyETGZGRcABzJxOoDnvgqQ7s9XU19lX/WEweTCym
hagEB2U/MMEpApag8weQijD7on57f3u/j8cGEQOIYWMIYvqbuMIeJshm6wDb
U1CqRO52obB1ZjR0uRy/F0i59VHnEyGbZW51cnoF9gElYIbV5zKm60TiwAx9
fFg+/L06bbnVvnid6bAdsqbswW5ko9ZZtdmpFCxwMBd5VKAp9n4sLD9osqdU
sDE622vKITCfIaKXtd7ic4jlxJN7/5Y8Wfibs1DzZyQ+kl1ECzPhRXvyDDaU
bRM6+6ZBtQ9C0NRa5T6aXRxmHCLm4dwWb2pWcmCB7NslsAxWpzbpvzVpoHWZ
d7m26QwNmCUi22CxdLjedKut3xVSa/nvEBpGsCEK8Qjl6KL00q++2AHyqZEi
J5DDQV9+aiyF51w2oU7SHiiDsjW3OCtX+dIme3D96Jdppd+LbvGZl7g5pmnC
5zSDffj1W3xt5a3Rz3bd2VXLATwFxYicu5MyE5VrXelelp84vEAj5Zj3Zx7E
/UtST69vsJF8bcyZzIUT/+creJomcvFWT4frN75CRjBXU7hLIrqVZOmEc70d
xrEGqBRVnURg46TtfoliA7w5AVBMaP2OSNiCwYW6J56HsK7LRtgBoN5zOAT9
+u5YiWUWBTv3/wBiJgRD+edRGjcGzTi7hnn8Xy/LeP6oW8PS0Y6KOgl+yho5
nhU3VVmeBEnHI9ffYFRgUY7qHiXmcHsqND5bDfwBrf834aBG7Lk5F59fYQ0s
ZSWcvyP7omDAVJkQJX8q2SECgdx5w61HUrXlemKuHfMUbARBpBAl3neRnmVa
QMBJgUNcJaSE3yzgLmuofLcrkawM1NAMjpcWHqc6/MxZAlbx3f5dn+/QJ2Zh
YCZ+5lkpNxOKuAeT0a7bVLNg0xLyE9GEYLa4phDrGo4ZTsaaaDOkyYL8VlHe
ZzUtvJpgH4EcjhjNjiT5l5WqMvHlWNdYhs14HdQII/rsGswshZoGbAMpWPEb
9ZnbhTLvP5fFoXy+b+lKOLU3uVlvWuVUlLRGDhSCwE5bi7KDH59rrpM7lB0l
JlVpmtAPQ11qcV/tEosSgcmAzZqeWYhmktQAQ87/5w4ibdZjPcUzlI32RLK+
sk7uS5wlOnDkHwomrMRm2z14kK4wUPNdUY7NZxorfYVH22crfeiuj2hhgM0X
ovqerOaxczfXcghUrGDDxxaRUqXp5NYYtGaRJ7m6O+5VchONgqRM5I1om2Bn
ZOYLO/qasNcN2p7SUNGGn4xnN/WPNmOJ7JZO4ZmeDkRuLOlifp9EXNhNlmiM
zZN9FiwHEPZI47yaaKkaIJG2sXgfNGfgsNuN/dtMO66Cf03gu03Lkrq5hiGO
2lVRwFO5lFHLSthlqQxNkR8qaInNNd3ifd7kKZs4SqQGkPDKx/MSnDFlb2Fp
DdU5rE6TrfHRJbZeS9ZVYFacav/Eo5AcPgvYqX7uNa5LWbRA9CM9bh505Ugg
ewy29vQZuFT3zOxkGi4AFjZts0iYXf4Ge/ce/hkrMQcNfFI8To7LR6ymw/nu
kKMDxxjn3dvEpzX/sT9CoxxIpUxLLhpEKeaO1pJ+uRnALt3am0GGGv65GDil
9OqnmcDaCejopAB1IoedyG9QPEKyFGACO3fwU5EOyq6y2Z95FUXKBtxlzU+z
90yFjAl7Qn9EmNiN16OMOolNNOc99IxIOnlGST69R3OGMMTHs6DWyKbGsJkg
EK5pqwV9k7muBzDgpcSCticT4iKlazY1t0xiFeWcvqG4n/5GqeNzAo2iU//v
SXWFON1r6+i/iQHYZpyPP5Tlc6RoaSGRb9H8VaqIZ7G58jDjIgFcedK7uQ5h
gg7jo/Sefy3Qm8kYtFwj8jqKkfib1l9Nl0Jx2+qdwEkAnL4Xlshdfk9RFXg7
RURUZb/844BkoLvt8l1VhvyEzwi73yZBTRZuAKMk8gY7kyyFUizb5N8al5Q6
jMTz1QS8k89SDGWZsvvOdST1nzogpw3CWRl0kDjAKlfrFuDWhcBXxr8/5ru+
uDVZ48cm5zfScs703mIokClD/BaxmteMhoPkqO1QRwpIYB0FYI2YBU5xrXOq
LMVj/Aj5vTPe72aqHlyEIX1EntWMN+7gBqXyWN86WXMOIoEZHS1Zpz0EgdJH
qGvDMMBF+BkIBIzBLcG8ptxn62lVOFyioF5SyIgUtXx83poNMZQT3yaExlvp
84aR8cbYjV4Sg2xgolaSaoOLP7aMf2SYqXngMpQ5GWe09CrOX0DkqRsP0CsB
JOMDXQAHKX7gVvs5gy7OdeMLuOPFiZr1bXlGmgxM0dD8GOr1mhIUQ4Y+jdle
eojQqMZUnsyJedCbskeoVtdfK4qYM90wF3668bwDV8wj3UzdyZIhYbm/spUi
PEIoS5rsMH9wn8jLkRFX+/pQOF8e3G1GXtdSGf6QL9pVOaesVFnjPEFc6q7G
HEkCfHnJt+Jdp50GuU/EQxxZhlZEn2A0WuP46vH1hiA6GaV72qRp4rsil0oY
gIV8ctIJtlzaA5ixFCSCbfC0CJlwUnqaW217bOcpvL3wGqNcDPqLuOIH+fsg
Mt+Gc6uLmBtJKymEtJ7x703HYg6NuR8pmXtmzdfHEg0+bnADFYvWgOmTibQu
Fe6eraCpMm7biSn+RdwkNn9Ji4AaV4O/vRbl/IRUTnnWg7fGtYxIeUQ8GnYN
+oQzJWH/ldlkRyXnHX9t7l7yj5xVjlspLYvBPKtXnXusjua7aEbdfbUp/N4t
xKWQZ2o3GOOcXijWGZPj+HIPI3EBOrdaHaFJCgzp0Nm9rFIXIqUGjLeLm6FD
k4w9AcCL33cKD4BDBjwCqlM3Ps+UYr2Oz05NJHARarXeyA6ob+n7F+U3J1Xj
/MivMYuMbl09p4yTpfbt6F0zTpZ0KpBQxK9642RUBREstb8BYMjcDtDX5M78
pcH+f6+Yre6tlOXGiaT2FPxpQf4tfhxXOZKuhSNedqUMo+akMthI0685eGtZ
GMOke+JGIaUvFfOAHnpM5k2T54ll0naQ+srTpZp/fxRDsWOiUioSxLXESY0G
RVOb4+ujcwWMxv+PCpMKRvN4Ad70CowsOfdS+Fc2WWKH1zenNTJ1k6DdNgOZ
xm/MNNmiToh+JlYOJWejsggFNc+GL/2gXn0krPaJrwFv8CyhU/dZqo+Au1hv
xdDbWt0HkcH7vPXqKM6safEJ7UwGH/1i/k1kJglNxw13KtOHRKdM7ErMuVJn
OtFEWgIAsJFhP65tMdl2Tphqo3TjsbY7okv48gE3IDsfPKrMEDb4hXyk5pxX
EsaLAClMYNY8sO8R6vmmfBEm8EABiIxWScUitPTzc9ahAbS13axqz0gKAmsE
/y9jYnDH5ejZpFIAUv03E9O5InnZwCorcz+y3stSrthmYj05tbYvAg0awA7e
KYuxg2NXmGXn5Thro1FekD3N1oxudJrwmH0qm/ihx5cmYnUfZ1IjpaXZnvh6
l7NZooAcCplTgrfGPlD3Zt0abR7TZmZw939MECTUgIwsaJPdDsgqFiqAuQPj
1vnOEast7Oy/fMBplDHb9566nFuBpyAEsR1P53C6MZYSkI7D6ebRNylLvBD/
5af7bjye0aylavy5pa/Kp0cbSH5iXV5y7xdAo/imBGEfz2bkYaPR/JJLklql
iDyCwuMLkduGeMhHvSix0DZiEvx/8LOpHz+uiBffMu5ISck3/ZdQ1bXlj88j
5bXj+UjpLgKNYHXOg1gjeFHEHtYuPDdH4Q2UetIaNtK921pYtr2ImWTXfbe8
Yoeh3jOtpugMTy8IiBYglIuDaiFiZccBdVwsVGpZEcaDql8qDTqhG5FuJKxg
YClMh/zDIJEYhUdPul9zui1ADFfTmyTR/vwPgaosuY6FuhAgesllBAjil96a
RhVe3m5pIlqp3DKhkAFe1Vt6LVFh92xCRTLzJN/iHtg2QF2wyyOj9z7GHSPd
4L/uA/vV3HbxEsgD+kG8dxv3TbTxKsMsvYjMg0ybreAd14O/ZORXBUfY91NS
CN/Q8U/DuXxeGk0F+RhRSst6a8r9WLnDcL4a8mpv4YAFMMt2Rtio9GRUU5X1
rF3nI9mc7CsQLvg1FujS3awRZi0hIivRBPXosvj+ygOIR8q/jh/wywOEZthg
kwmOLcaAv/GFusPvlhSaA9uwEy00G/IH3JEe12HlJP/zf/bTk9FN8PHpQh1z
IqdQe4mast7XxjVii7+1+hKZG3TxPNr+j/E2t+RIxXiCQG7w+E8ddLwCEVje
9lEfd3hMaSo+nO/6GYmA3jiQoCJ3Unz55g+dSxNcmnz4653NUnMmxYvCxY5h
0D4/+rXCSTGMxixgK7ndzHrYY5jzQDNzD5rR+sTsP+37WdZx1+uD9gaqPoGu
SHOB7ZUYslNIYuFECbilCZeoytwv2vSSneJmLR6KsirGRzBVOjXreUmv1ZR3
m46UTOlpmw4Kl4u28VUkbmhpg0LJfpKi7kDgSorlosuxwmQRhxjsgP+JxKfY
Brir2BCdE9VzH3yo2TFgzgxR7RGQhprdfkjl5DjEu/7olx23s2cmLvOQqrfP
VZ32xSBo43B0rQi6ql9SxXhXqVSU358JaycesW1XIjUs5Epf3JYsTP0BKYd4
mgO7lE33WXEFOQNvx/ouk4cwkAue4YNo/k6vzGKJjVdhX+6esGnrbME648No
+Odhnaeqk1ADroGd1wPTE1OZhKubj+rWtSBKjYRIbP4Rb4Lr+x/B0n/m9UWl
tgUTDeZ9WUgTRkKFi0QA35C1ZOwVAEfxPbbBURKl2tpICJiADS/mCAGFB93S
ySOFsqJuOxFTZ2S10hMZ4DLcndzxV0a5DdDDCaYkaQJ02ZeTW1+V45GMd5mI
36sy2Hd7XVyRBYOy7I0ttIEhVT6cvi7R1qW8fhAj7eAshbwTKPamINgN8ygx
NkFNyPmTefZR4TU5KbtloHTAFESCSv/9qM8pRRtuRJlcarTKGP3Eseea5AkE
gs8f/8eQEUDOY5K3ztr7WQMypH9f4lj1sJ25/rjPXokzc+PCesRyPR1e1PNQ
/c6fKrwxggSXhCem8mrENy0t58TeYOK1LqD0y4mXLqhSbgTasFc5L5pXMF25
uzQbs1qyFhUu60++aFoIaayb2OKsgu+NsEhY3jmmVdKWsh7SH3UUg2xQk0eB
dumuMgtvepJj8GDym1tezELJh4aMJqtGvr764w8CEzIuO9xJyr6XPIqcyvRy
LMeXBdT1PRxbwCKkQYq6Huu3S/y8mjfvpj9tNnWmArTbiI86bgiMFaprZmta
5K0d/8Dl4U0CpL9SH0PdFbe+l5Zb6i8sK7wr9JVTVqe1xDSTo4ZDZ+wUpuCQ
JjjSaQgvADgiEDNQsR03yK9btUIDyarmux/qh0LAhHlcPs6sbhChC81P3ldw
JuykmnsSMddaM1E69w8PLoV14kHHAPxHUe1S8DolwBf00yZeNCNVGON4GJM+
8yaHkZc/53KzjrEVdusJx1u1PUUpQiOWpX1W1bIcVi/i7fW3eA1os3jHZQTH
PWnW2HlnB7tH/Ms3ZeNZ9DgtdFWlmnv5I9E4JV6CslcJVYc0e3Jz3Zu10NZe
kXR7YA+WBHPwwbo7xWHE7U9IENJcmNihaSJfJ91jQWPWfm6n4JZeLUt4vVMx
xqwcBEV5SgdlRsFVzuT3d6hJ2TZdtEPhfv2zSLexLPtpwZHXDkzxmV02lxrd
cwJq0BIJIMSxuecJsugXNoB4F526om9sjo8kKDnSUb22ScwKwckWqzEc3Jt7
CxlqNqN6ywrBwFTHxrlyVapF2wM9juaYMJA0Gt5CTrlS8mR9kfD7AHpjFHXo
8foVxWC1OxJoqQaUL6hErR7+gSb12/P9ZXDx6tG3GYcR41/OE0vVae6x/yJp
c5bu+vKB+jIAhaicdPPuYjSagtBUr+qvjP3Hc06sDMbDAqFUdFTDKCUM1+eG
NnAxCUquj5IPCAb5Pm+StrcmazdiWCD4mU7zua6fzQaS7oMq20lmQa4CO/mS
omVeSPkByANwoyBui1JezPaS2RZ3vkYOZSS0QZWJAHuHQ7PlerOn6WDGi0OR
gxDb3KBdOF6OAPEK5JSHAaLHGgiQ3eA8rzzyaOibuk+AH4WEQeEKQu/JmN5U
Y1u1QTkcsLYGrsm/n7Of2hMszWG1dcYu61v3v6QcY+vl7ZCp9DTgJW6nDCbl
zBH1N6mC9rJUfpRm7frGSLCw/Lki1IxbrUAHYkzTn6SbAkh0M8LVgGuljreK
J/50LL7g0VgSmudK/YonJ7OL0j3t8oYNa1hdlM7CZEDKZcCL51B91n6XiL0f
Xs/vdKOnAfVq4nxCwbkN3ST7e5HdXUqkUuxivdqMOpNlxL3QjFLd3UcbfqUx
HeN06yr3FY9MSYtkGxc95gUbGmPVsktS4/giKcTB2iQz2aHfHXzBqkPs5/Cl
eDWdGDbgzWS0U8yS7dlaeXmtuwKNXwMe0t5DirqSBfOFiLl9ud2dyBki/X58
N6D4RXW57LJcWYw6qO4YVUcqev5AQacaz+DXfHUMoHS1cK/TuRPjYT4Px2lX
8BcjA9FWZeLxKdAPjpRP47Jcry2YlvbVxKSzSGenvNNIq20m3oXUV3soDRAx
josrvBAvWafcbFrFUaLi1qSQTq8YEXaXO6Eud/q7gf4V36xUR6kHnc59BKLH
K1FCnvfiN2SvWo27OnLlguW4131vOEOmhRvwWz/SEUZaUT+j/rVIOWHH41lH
ACXBlR28Sy5a2Ye1nbqpkjfPBF6sNAfOaFVz0R/ROjm8gXJp6XxVndi5BPJ9
54v4LDe5ahgq6k76lQQ7dnJE0US41yIlqOPW9b/ahBvElv2Pu/1sw1K7CeB6
iTK109Q7BCkAwU+o/KPxRVI00Z532Vxq0NMIuyAheuqHhBynNI9b5NZWPw5c
/FGSzyrQdc+97qAGXi8LHQjcahOPYUYLptw9wGZfDrMUpT+MdolRVQa3agUE
MUZuwjG+IprMS8JOwHZD4baDaKhgydEYrate+Wkg8nBCWfGeG3tOLypm0rUA
idWnreta4/Toxj+O/egKSiWrLdJyZ6J9IZVedigOOjkMyY+o4DGX+OYznZb0
se0hi4bxSmfPTMcLs30rcxEiI1hgUBnReOCsMHRO5PbKTnTLJpyqagEWhsAK
Ksss5S3RHhSqTbL8fFseeQUZqYrTHK7eyyYwsRa2whH0xqhxzPYq/brPAIEa
j1X5M6piUaTMNhe+7vxKU262tPaFschNDauwBgcLXP1CpfKX150UHW6dVCbS
lFyfu9MYOc1e0zktZqjlB56F9d4eRLa8ZteIrZMjRPEtaeo7PuxV68vitRiw
UfXVYGHdSEca3O6vB+UJgG/uf+mnwXc3i4NpFgn3fMQWIuOsKExW3E7B2Ptd
l+frw4NPTZ6PkEY8Rf4XEJ8R30ljXuxtwczdF6KZLg5E0nwD0XxzjUD8G3bu
HkBO62Nrs19AF8fqyHesAljUgrG397dZMq8BfufH9xzTYtyBOehL1FOGvS11
mmWeb1D9b/QC1Y+PRypN43rtfCBs8YoJQhtyLkmb+kPTcUhXmhxHNvgwDbLn
iay9P6j23OKXEBf6nsf7+MssUx7gu/OnAcQBL7bfXbvG6NBSKtpydRmMfKtI
jj0/4vbnABIK1GvHWvEpgPGIlLcjVoGObuwAhXyvZmxI/GyY7q5X8rL4Ee9j
QUTAFaOREPYrxEs4r55xaMWLkHPCcNHknsneC4Z5ZMfH5l+CwDHqtYGev80D
vUTFuitUI6lEl//OAAO6p9wzmnOleeU21P0HaFvQjUqFlSFqW5hLz9g4MA/T
MOfBsGpz0DzwcZ3FC8PMqfvR2N8fDrkwy7X5qAH6Gjc7H5+yKUNs9BYkJxxj
nTJldYSZSsgsVdyECkMLf2V9wgMrp0wZj3mw3GsB2wJuvl48pWVu2rNvNwQp
C0QYDUSvnlQEJ3czT4PuHemN81fJIRToPNGhwReprG8LnZ+Sd6PHI4pGlT9O
NoToxWTgyAjsWKLDSomDUpqffzcheJ5J+o5jV0WWtHzkZ3wAB2v2sDL+zSrC
9gDOK/LfYpfW3MaU1WFrh/0HplxA2lCQypsxDfvtz3ChjRQT5gAzlQNiU2Ly
+2VYzM8zp2lb2e5KCKZbogd/RTCBv7QNWuJcSGUEZoNIhCmq3iNmdaATl2dX
yA1B3bdXi0UzbNne+nXEB5kYs2l4Eags7PQFACqoo9/2whZ0GeICM3AbysAg
A9FQaKOAr0G/m2d6xwN39FlZw0HSdyIyAaMy2zGzZvLWq0ikx+o+QAe4VUxl
2w932sQOZCpOxW2peycWQ/uUmGcD1bpwv9Za0GZxtMV3sktpoMtLpxsRIKYH
260aT8b507dMT7llHuTeCuWlMN1CWoLQFGCYOjpNc2zWFoJVKRIvtP9IFNkb
EqR7ki/sIiT9d+xmQexTqr72m6n072CFB9uM6LKxtU58IxZSG/mczFrdqUEK
CQUsB0AJYwXAJIJjG4aOTSXxCoc4n7HkYVphoh2Xw6ul4FcHHcV0nChm/dgL
POxidIYYfRMhWr4ioRLg1a33TOkUViN6OF9hX/jHI6MAhCNfwqvlyQaXRzmm
BbA43/ZUivi68J5rPfWu/YlK5CllUZHTqyEwwHhcPTGy2TZQMAoVQMg8UO2y
t+/DEpc+IAecttsEz2cuwX83BokqTHx2IzqcPlblaFMKpMfhfdCtuoIDUC3V
a7uR9tQvUhjJUrn3Jj1BmpZ6V6+cmuQ3uil2FNYH11lGHcRgSbe9dYmKBK/D
e/hQ2kk1ukzfuOl2AFR4Qtd/xWPeUFIKeyIr9CsfU8DJPi8NiBtb9P/ayQ/s
e42lCLZksXdArU2+H3IXj6GTO+M8U27UHn0d4C3BuW0L2lzp/7n/4U23QUG8
LM/lXzrs0xdJl+zSv0ofP/AeYo300VDCT7JGOT2YnGPJ2dd3rxVEKncrU03X
vrrPhJ9jcxSn+gLhXQtq9vfh81R05icACLaFH0/j01lmLZ8P/rCTnjVSYxRw
ukuKHbqAZ4yBxxNju+TB429PYPUMy3EJiTqdJXaf2UPbU3fYjwOk+3fCqN3Y
k2SojR/XJ66wFXu5bGOC0d/1SYsqjzrNPe5OYdXdPC2o57i/zDdjsspkoLF/
H4V+09eygFroRa1F/UJntV5gZwF0/05LXmqLJGwLq05LwGjxnveT6x/0nhLz
8+Wl7cGekS8A5beySQxG1mUUItMlE5KaYJa54OvXGNxPi11qx696v1lQ2qzL
5dEWTtnyTFpOgOBfuYuEaEq+04RI3U76bKfYTBPur0TG4qO9oFtXCVnDlQ66
BfE/oNzaVy4WF6r/fkQ+EAV50m1bdLGaAidvkmWT4EidbxqhE+cih2V/iWeE
XuztJZa7Ku5JDK77iNZnVhxK1RluC7d7/wJrb4j82QspZ3G1Kny3lYYZdaSR
me26cDY2O5YCWsP1fy+o2UgKQe6K7WjJU4E9hXKleTAj9z3C59s8kG5F4rAz
vZ1BVes87JK2AqiAevh/+qaw85gYf0mEVWiNV6uxjGp+CypmBzZ0prIPGs2j
Wqu9ScEy2a9CCsdYipi2qedlw0b1rPq3OQWh/y31NLN6DzSVXfnDduaTJKAm
f+p9ANqE71wRGOjEhHaZRYFn3iq4x+M7mM6TaiK5GPelqUfc/4z/GmFmI6la
aJrN43bh1r4FJkPp6bDuIY+WnH8+NAWi+cwCTun4H4HjJpyCn6CErDPImWXD
Dg/h1EW5mf0b9AvAzRvWjjQjqFskP9purtxp1Cz19kpgmcAEWYy5GTuct7QH
UCwbM+OFmB6aV49vgVAS/M1i0N04KV0NR+BNgt9AjbQr58e90C7QylLNcKI+
CvT30L3dGbGt9zCz0zWU6niO2yleGv82i4svj90s4sJK4w/uBn6OIMVR0nLQ
L5SKWPe5xJe03hxxdIVS7QhYXp1mLfo843IbS82bbS/WcoKSbYjWWpp+Ysoq
Vnv67x9nV4z70rYgNQ2u6vmzXL5+MMhkBWYoNU1/6e9gUfBUOn3T0iUCxh9a
04fd7AfwR96ISNJmsWCVxWZ2SpsEkleE9AdEN7egH5gnhQSCk7SMyijJuJFs
+vdSGuDbcV3UbkF6I06byVbvP5USh9RGhiwDcPommRgf2BFWPcsZiUJK5NkA
UYDqKWIpLQh+xe1/A+5pz1iEOpXaLDkazDU1VwhdFIyHy/870ZJ4sxx5IaWi
Eati+3Nd8XYDHLGjMyzjo2Yc2eZYrgvPiWya5k7fn6woDLb3YthqUX4+LnDx
TqY/72lzFmK+T6tdamEXJ6hPN7FxOFJLSjN4dniMOfjlKR4aiSpHdcDTQhfJ
z4YhDzg4NPP4dX0Wak6VTe2N4MnUuYv1ajpATMYBacCtQzITXr9t9NWGhrl0
K+6u0nbKl/2/8TKKoCA/Ao/Y11L95hzJJV7anSZRN542cJb6PbPGNNJEaVlj
yxhSegeMpowlG07+smU2EVDi+uZW3OejeDV5w+KDYgQXlnZsHfsfc6Me+TY4
xnY4QfsRMuRubA1ba8TLqQXIGdx2CeOlPfoHzZTSitvpSOQJgts48mKSvnw4
AQiDM255FBY7dj+e/4auFVMJBQcMA9tGsPiANA/xJ0D4hYUcYZr7NcYuzQ85
DAL9+bES+8R3cu1Zap1gDU7d9aTocp8w8AXDmYU5hgS7iuo/nlCmicyfJzYC
UiXpMRJsmD2PE/OyaoqWi8z+7bf/jt3J5RguW4T3z6ONvJ8VLLBe/GO9ZkXl
6l24V0nzm7+477J5oKq1KYBltl1t4bE7gAgxOgkoapv4RslC9j2epGuB4Zz3
cODWY7UQ3+6H7NlkNBO5wbO0jOIxAOSGC2f1fnogvr4W6QN7+UojipiGHcbx
Mb2yjm8iEiMp82xVE8BQQONr8lUGgdd7y4FiOFYaThGQCdaQf5WvFodzv7F3
RAw7jEUKltpPmyruRiHWxjO68x+GTGbfMO5ZgtAtfLEKoFLrZ+0Lq0lBKUgL
wBVhCxazVnZQdrrvh9HXh4EaDBXxn4yHx/rEcJMFpZCLZmto6BrVDpA5/p38
OHLTGgjcgxb/yrNJN1veNSouJ20MTh97p1EZU88ssTtM7kEvruqaNQ1WxpDb
X6PnTpH4njJqqBsoPkKjRTQu7KWEilHzFX1O1ToMUmQ+7qxBoQYG5gbeqcUL
sOgH2kvG9vsuC0TG6SIh2ZrGhbejcZU9LOyDuo4YREfaDJHr5XY5v1eUYhPY
KHvgRNlzw+xXKvUM7WYSlZZ5CUDgh+5+IixL9cK9wtxOJHN1K4BzWmJxBwKY
bU6BRESF49F8eo9I0Sb71XDI1Km9di8RVONALR5QxfdnTHx5dgCfXmG/XY5L
sofh/PT98z0dH523oOooVIHejM+dQ1KPf+oJPx+JTWFCXcNq07mRkkORrLy7
SxaZrz+laJ0ProC5A8gCpP/yMAIKPE9WXVUJS/EXDhH5BKk4eil/1zGFo/uW
jBmfx184CCIi5LnMKLZZ75Tba3sdowyraKgImoa+7ggVkSiLLvui2u7hcXSY
nxiWDkEqm87uZjLlm9QZLQu4ylYjapaE1mq/iJaoFRiVJ5NJRhn1hcWnsJTN
Uzk04s492bLf2cGCxHHkhwX5YXTlq/N7Ksj3NijvL7dHLPUNJ9vKzwUACJhG
0SonqyKHOcb4X7M6r9xfwIXGGzwVMb90pd+s/MPAPXeC5tAx68mDLAt+u7nu
4yWbeUB0sPPDjbOd17W2olVjB+UpzeJZYWDNTepRhAKTmQ2DxB2IT4gthGsr
ZjbWJ/+ChGWrXxa7AEK8MaQIUGRQLAuqX5+f3Zzw1WR7MWeRAYdZiiD/HlwZ
QEM/A6DM7udFSFV3AqmLfq7O2bNGHFxfnBThvg1jnYa+NPadbi1mAw1B7zZe
SABQSCYks8IJQ38jycRXhFH6E6osAySdokb1mQd+15B0RVQqNNjoW9I/n6v0
5MBrMIW/OkWo5oVMc1xrk1B0hmHxyhB4rokc+80ViWuvRLxXyyOR4njpNomn
TUVKGTZk3GIeWxP952BEZpXWqZHap92BOYLMIkR2sCgfEef26S9nQJOqaHxw
UdnLOFYpGF07DbwIZSgs1uSMIT7z2og92LVU4w5tHaqx4yNhi64LDfUsQ5yd
necl/E3EE6nVgqc+1H3/W8AE9aSblJmb+MZ+OkxxJkuXAxv0M7czS4YLg71o
XUnsHg8N0IwoiOgBWHhXjog4Q7QWhAm4paGUbw/sSnrYeVV6Hvy0gMwDV+bP
ewWcCnPlZhv+BB4PLD4zPLFV57hlrCFj6MetTlNlp10Cv0sf5wIT0pXjxo65
FHA/iCnlBtgg1VaOR7Szt0R48d/ofurznIVw2+obqKIiXLa+QVq9X93Kvkhi
Dz3t3P5NDZ7HD/HqnHdfvWR5zLmOus+3DbH3F+KW0lw1MD+dishvLloxFvoF
tJ6hX+GOqdClixATeLhVIuF0+qgG6vtTKg5Ww6FXNTaApSPKwkbamQF+Fezf
Iu6uBAZRs0uRQxq8vCXmBUbbIikq619ZsDMRJw5+CkNjA1INeFVACWMH3yGU
Awb1lrazgIs0WzT1dc69qBaUTS0gaDN0sbVN630O1U1frFE/Xv3H/VgRf20w
2q/P4L3kwEn7X/PgWHIJVcL0WaxnSNTMnEqVvbG/X8Jjif+Mws4QnJlxPxDN
UT6m2vYXQMG9k6LWwLBv4s6wvInEJSmfqQspPaLK7sY2PxlPETn4nGyoko4n
irHDjShQH8Z5GTb+dCtUnpvG/t+ApzkUhWVbKKH4RXERVmWnvOuV8z3SA5ON
LXglfp98MTo4fuAPQgU6awR+Jy0Jki4Sko1n5D18Aw2LJwA1laQIQR1uqAuG
gbcYqK5UgPOOda4dCD1TEE6iMPg2opRgd3RiRFF9zXfqYbpBY3z7SFTSyzFo
HlBw5rd81lk7s/8AF3xnNEf4LM/3vlCvTjCIe4ktEKZ/wGjtJlKeZ7sz8Ah6
Jt5jl44Bqsp6x7HaazFhsz5ZO3xlBIzcBJnu7rw4ICkxEtjTVHv82RlVRBaK
YRz2WIeurdeaXesXUghA90yaz0OJOrxbL26QaCiedo1Fo/Z5AI8yMJZj+l3X
YtfoEbtB/OmhZqUz933DHCUnXeLS8SOwg6g+2UHTaWOYL8dOWOAaPFjMueWj
7BA3yIeTbI76UeYuwMkfHn5M/Z5UkYdE5fovXz68KIHR5RiyJo65xe3p8v1W
l4HaHUIuXJKvcZO2HZP2/GNVCoU8nsRwBN7DMZTYimWZTTb9BmFOBdiysL21
exzAsIHCrh1r0e5NtyuHgxsCi6VDPC//qBEh8aarnRJn7hDYxLIfd4sqhuXR
XG8Dnp6aicowKub4YahXJIx7GDOYTp4mkICK/n9ObcaN0MWP9ymHFjgjUaaP
fM7zSw6yCEXoqJXSVjY235kpaPHcmVQTBLznYOc3y3EFpYJzrEWLLSlc4I4A
pmibiRdYqrPzOu81KIayR+qXX8ELjWmjGGsnh89Q1vj8U3SGQmUQ7R5afPzB
eJ7oNtXiM9sPlvFrCfDQj4/sQ80yT1P/5x8TeRKDtNgDc2v6j/wmuhChQDId
U2RAzhKPHYm6IS8K6o2j1WN5oGfQD2F3Ls5yXitKKBqIfMFaddiY2cLNkPin
unptXh7SvzlX+HJJDpNQ7ddCoIKm0LwuFISvpg4F+Jlk3Ktvy0VQ28hOgKwQ
sypbGXNUN92F5m+90slIzsCqOSSkqDEuBvlRPW91E7kxuUQ/D796M/NPQCv9
gt0b30UMO3Q5OyHSY2XWAam5eC2xaavYpuiElMVzuZB3hyvrTDux6AGsYYqv
J4JyvSVmLqJkBtqwsQzfWegPylQmeRXRp5WJiRRSUCFLo4Lzz9rGPgsFRNZy
URoht1BNDks95rF+wWnjcCZoyE6YEvRQfVl3aV8IxPakRjaytUFKaoersQvY
/5pGoXk/sEv/Zy66mmhH7qZzBVlgfAPWhIQw/U01m1UENZaoy8PGBKwd0oeh
w5YrL6kbxfVW6O4BHdzBh1jfku2rzvAIBasi40U/oCgfY2PiDP+xBfWyJ0Op
WSIRmatqKLTSKFiSQ8nBULw7A8OOlmHaOvxshd1a8X1jl+o1IwIZKIta+qgp
L3maC1BUKYHiPgVjL6q0E95T8pYukk1HwPlZnJOf7DdWBxKPcMJpcQNUqQvr
yrgOzuNZHsAbnuM+hpYHH/tcxS7OzNT/lxtMlilJzmpGFuQYuyUPMNaEVPrV
ZN4Gl2sOplX0aMwBA68yb8k2NZrt3iC5WJga5noIE03zXrC/0MZE70PLgyMW
FgJy2ujkpYoH3eU8v6szVp271wAp9mE2XotdTL+ksmkxyqBjVak6u3lqpvXz
NWVQX56Qf9IiCnpiYnFny9oMjFrfZCt4yJ4NxrgPE5+stDlajI9gjW5ie2e/
wap55rKrguY16IDZfs7k29EvZzze2atMJjufAdi3fqmF31vq3itAdeuQxbdM
3naXOByYtb8hf2eipReUTE/YiglI9KENC9LK8zsxqAZU0amWzIIDLvZ9tofJ
8MrRtG3cEiOzEIOikp1hiEdw6QsqV/lx0IEjxwnH0LPSZb13XYuWdTstMBa7
d/n8v+yjVL5Pxyyi76UnGqoUQVWT5lpTl8dfnq00PEzswOBByMKYafcPJChN
5dbGAM+7aql8cViWDVuJFBpjiPJr7HF4ZsQvg3u4T3OPS/uuZ6LLCzfNeHro
qg0hNk0szsEBD/pOnnT3hkeBB/X1QA8ktA3O8XQ7LnW/gePo7oUzRm8P8RjK
LufOcSN405VQr/+VK6WResbcBcZCU14NBGtkxQ9eCwxdD7+eOgsaJ0TenRmF
dgJuYNa333bc1RQ2L+lmMVMXXcM3jdkZa/Dc0K+K8pmFmGkbVTW/VwAUBoi6
++x067B8Ea2jilNmM85Vmd1dis3X6Zgon74O04x53Nz3PJ0LWZZK8nZSZFJF
WGgV+2xv8lJ1dakJRb3/5eQ1qfsekHP/JNAiR2NwNIyX2Rv5D1qLWkpYEiQd
odOtb9SVPNHZkbsh4cDXcFjLQBzqDrQQWHUxj+5wUSURLp+3CvL26eWFHg6O
OCHQbEundntNhO9CR24GFf2LJJ+EjY9vTo7jD/1h+dR3dV91T904/Yxt7YpS
3UW1azHQ7GTleLKKkB4VnJkSN5Pf9a/Fv6KZi9n1URSB3cB5YQB3TpuSNLz0
ScdW2l5N6hGwMzT/J1c3ydO1HUPpxt2mrJql8khTEr/bk22J3FJlsSB1aq6B
70SXb2TOyZlZaZQaBS8XMsqSoFYRT6lhetrBpo+jqIILNtvPZUIlNbkC+hqn
aWJ1NY7P5HMqesGJFXiD+eWoy4aDBo8uZ9A4IE62rj7nfcqQTY4sDCxz+MZm
qiUgly2Bw/5vkhAIROn10aFZ6zHlBu0CuWjrrC0eXZ2O7kazQmkZiojW1tj4
McsvQRr8cejZmLsTlSOJMK9STgJ7zPOd9gx8TufZQEPIWzWKyfTbT+0G5VTh
JbSHghRzMCKTJpi3eA9J75FOuF+Ow6rXtfbJeVB8mNAV1h76O6lQ9l6YTcQt
OlXw4A5Yd540rKU2TYA+8wXhMlVqSD3ty7htAnRw3pyQQMQrTP0vnaIrYWP5
xOkIp9MUreR/rRBKYwSKsn6CsnPSKKnJrkEAV2HDQrmut8ts1A0e+nDuq0zK
95u7XO2sB6xovi2SRRrEN2KJOn8fH1QiDLHvwHvHxhoQp9L+0M65h6yJodbu
q/tJScjx1sl8MMWxipT714ZzjLFhjTVPogjhHCe5ugOAbjLQB/m//oeeiofg
hCx2cxxt4VRNVz6b/r9XpdfPT8+TuaXrlXJLqTEfKKfsEGDPIwihmDbY6Xvx
RUgSRaH2MwzcMPjo3S0HOQ1kT+iVhCRZj5Fn2si1RMm3zL5KOSdIBIoOfv/G
6kD6heDDfXBX8JcfzLMeV6tvERsPWfPs5HsWGpb3RNLPr8umrbawjxs0urHR
RPvl9/8JSKiFtpFw4YZAcKD/itJQFqtfP3MPaglCshWuR3hWZk7jXbNuepT2
bTcAq/TG36udWc1a9ish+QBHjsO417Or5Frk99hs5zgMri9BMkenghZyo4AL
C6wYC2fb+mkWkysX1An60EnzFMyi93/69s+Lhh+aFbhA68xt9Mo6KF3osRjE
WDLKVPgK2ErBv6/h+v9k68bFuaFJNlw/AvFvuw3hJCAFa7duuwR83upMgtlo
hxWb/Gv0IrBOj6JYRsDBnGBPHcHnetxBW5a2pMBF+7ciLAg/9WwLpTxp0c+q
ss01l2q9lVHfeVreGdqWoNAavwVId1APSR0PG66sS7j1XlsEvwxUIB7flFvq
TAEiYc9ml0urO60k5T6/mgsikjaOK717FeZhReeZiV4cp+mPZ016CicXIebr
8jbKnBKL0j38r/H7kjTBpWgwId2fpskpeBE7/8INqkTYTKuZ106hRnppWBbm
qH8YDAb6d1V12iy2hfuoe4qsqai33CnEh9OmnzHPcedbGj9mRjU1I+Y7XIxJ
mlerIXlWB1p4TFnPkM1qMX6gm5u8nfQ4rkc4mb2/F5C10W7efHi+fp9auPjI
+DzDWT+ckOY18UokAQ1Pc5hPXjxlK6bgDBrUBDfbgjD0LBUWTjZWb1eKGXoZ
1GPiz+cDsoYY0o/xI+GpA+17mk/m39meLmAgVLwWIafroxGOSpTA+Zqfy3GE
z8RSDFS1IYU3n5HC3RPtvrbver4AaBLKmQUt77h+fpvdY1mlUW754E0AR+zO
Tjex0bL8wHM4c/wcM+c4HLH4AMyzbWHfRsspUQQxMaWl89/3DIvH/0G6IQVw
yke8i4JoC0vZZ4et327RLM1nuR5/OV9+3g21tiP2AhCh8tJi2n2k73dB8KwF
sWju7ry5rGxXdnz3SE2YkYIl1Eg4VGEpG31FIsvyESwA9B5MBPl0rB08DHeP
P25OoebAXpHIbItLlunIEDtCa51bEO+cDjrGk7JS2eDhCQ82tpgznKY3k1oG
gRFJlop3Kj3uTO12l3RRE2j2NaPRokjxPo5GiFAGNiJKqi9OgbOcNST/eRGv
Trt/bj6tflYQ0nKtkRMR2yAtCTc+DsNiHlpNb3Sk/MTCnMKvv8B8mCPhcVIb
lqBEkHa+qhC85GEQBqx4EVVlAKK8yv4bMf1+6C/cyUjDTX2jEbwV2BAYxsaw
jPnv14FBSknBxtCOLlHBafckEtdtyU7scGxI5jH2SDPnMQnKlNN1d1UFJtVw
5W8DB4jSrsNCfyu/e9pSjFY071vGxw2tPS7r1uwg5TfURbN5EaS1nfEdwRd+
8hY+ssyf6GTZBUqUXW5ZNfDntKMv0JEHeeVO9g/aewMTtbEPRdDLdvCGGiuz
SsxaCvvpRzEl0LcXNT24dK7/P1B2ZaeEJz+zFYyQXCGZfTqnODhXkdsXDoCH
YfSr1eWJjBZ1OjqS1k0tVw+G02qEIHa4xlHEBMwontsh/N6dJ8+s9jv0OQje
QfWRczU1tcwbeKg1vDcg2kg92rDyL+szLE/JSvo7FcvN0QBZi51k2THLFJ0p
UCPJsAdXKZLfQulMLZ4vdkgYVKqq6RrktMxzbM5OwhYKoCbQMsbiPj8Fd5HB
a7DdmFyP3ttTUvSg+myPUUQb6jH8nEkcpsRDViOgucapiS07vCvXQsSWe+Zb
CbCkxA6mKzX8U/r3BismEXa99HQ96aEhSPnv6ncNgGDqsqQYc+PXCspsdrMf
pmJBxRefgH38s/V1yPssahx602ABbdR4CwGnINXC1yjwiHpWB0gFxry8YYdK
b6GoJhl7qKKUnCII9Cs2kT2ZIcUVUORg8lK9poPK56MSJHg6jt9rOrpnyZ8K
nvUVIguw6E84t7nLS9mRG96xCo9RCn+UrX2zWN/5XfKsn394UT2lV5yGblB0
JkdvqFuPFO8CmFZFX3hEzQr9tJp+67/1gLQ+8YD9H6EyHyz9OHum1EEEPq4r
HzEmDucspqwNX9f2RR46aCEwK5n8MqTb4k7ZMlYzi0qKZ6cxeuOjRNtkGYvq
5myZLqhx5kWo2iZTosWE8MUA326Ayl+DSOhzLfkeLgB41gyDWfoA1+xtrlka
sA/jmnwx6epRQxC9tIAjdlISSs08FacevGTIfJrzJiW8Fsm7M4YLwMqWMdZm
k4Rd7x2mnsHsm8GetX2JLdyk5J1KEpJqbUOdipXITw6AK2wLpp3boahS8CIf
V9rmpWIA7CLeMQ/jtiDzCKUGVqYmFTk9jUYPTucid9HliO37RcxdrlvlzY61
02NpmcUJXN37zzLVKCkphUtgxEH0+K2jb8ls5b02sfEpum9i6/WRuKh1KoEd
RxPdWbuSsDKj6DXPnK881QD4rPY6kDugsjskKC/g9s46unKhK0gCqhP5LGqK
DcdFwVLWppDF/RjsKUH7wloevx0Pc91AuKRR/PpappZdrpr/rEiDz1LIgyYO
CJIUlEmW/hEcT3hhBpQAYpPERCTC4S/CbJ+xjUivyaBCAffTK5E+uqS4zf5r
/pmeyH4aI/SPAMQuw6SkSRtZDHZv5ILd270AtzFyI+xoSXLBGC9zDliMKK/j
4QW8VUvWq/x6VbLuUMLRjvb5U9WLd5p6owDMLqfZg21XrUOBUi5L5MArvAOk
6QbxpOlbOAx1ZLbHYccPG7pzGgFh9+zHli9lj0Hl0Q811vc9xht2kkGaPhpQ
URqFG6GTBBpXt3aAbglRRxS/8UO3dJ/ghiLnHWlFDs51rxGchek4Y6+yamTD
ILE26+Nw9LYyVccktJgbIiN3C6r2smecv99TDMZOCEZYzu0YH62k+rOxIbiv
hQ+Euw2sfYnlyaDPQKaV2NHYGn5RXaCYG0ssKbP3/qhVVd1B3v7ROdKGo8Lp
LH8ozDFY2GbBs/PEDXE25IjRD+uG9xCy++JRsvIfk+E781Ph8jc+b+/V841/
jFzjL+musrHsU5Wg4DRagR4HtXPBfmGkLdoE+pWtI1b756MDmbmILJLh4mPs
q/gcyXdYQcST1pxRBx2Y5lT/5W5n44kbFNyiJz6P+PgNGBOSdlW7CsQqO4fM
2kosUq8rCWqgDufnEYc7FfNmK2Y0iMqcbP07Hv0LRfwkAg8Ghik/NFBeCduw
ZWgDui6pPBnTcI8KvXhMCChOi15ZmDvPLRdR7aM4kozxVoCA9adzi93qRmiN
zndFpkNUmdGauvQx40WlIvpiX/qYCx2RTLaBdPBVt5sIkzium4qYPEhj1d+Y
huyYiHZx4JewvkzcCxusECGGieyv8Qpnhfi9vXfSlivWOnJk6auube2DegEx
WDRIluJNqArSihrjgIfyOV7OCzYvDPetziMj6dxbMaclCV8uF38Tu3beK5T4
Fdsjwaw/BrhZtG+59iODZBwGF0taTPLpSFay3V85GnJ4WLVrPUKs91pcyavX
Jiq7K/bIXgPPR5WANFFclyZKE2SF5YW/YaaE2kragScH0TO7Um5K3DJuULpI
PV/W6wJCUgAGUyzLVrGi27jrPducR/sHq5EnRYi7UTENrNWktQm7iwPoB8sq
x0YZeGtzxZ6GBYpi/1M5TH+dw2JyUytKwUa7fFTl6YbJDY38rUuzUBWijfvf
FbppUge445qBHFOCKTtJPidCI1310Z43AxjVC9DKkWxUW31UOBEuMjBXArwB
9ESOvdBWQgpPtWmIlL7wDVVKAd42unDcWLhRxRHy9qxWxvpAgMzxDfxr+YgY
uOZ7nm6W8zefeEtgS/2Olkd85BF8j0/N7DK7J/jl43EkKUZmaL2iwwZudDN/
z2ISQmsLhOnm3PrLlef34OC9lr/TAJ6MZeh05gd5FyO5sW4QWm8kbmxi02LP
QDPJvyEdKs3VfyyfdvdmSDRCQU3nsIxzjbC/bHkMR59UACUVjOvjDJbG+k+u
JVD8qK2ABXj9xQG0t9VQzOfDGtSljY2seZeyNlIKu2MsIom/ubWCfSJmd+Fn
TXwMwurYGgGRbUA7izPXutyPIkxlUriNDqjUukT6EzTlClLbqyb2LDdA+++7
3irHiC9J6XXH5Qj3qzQ52ENd4jzcm3pa5jsP10beJm7tTw0D//dttyUsFY0I
mrmqZIbDK91MLAx5wC+tUQClaq1hz8ESZCJHpr7a5C3VUiI1mQDeZInRM6Rr
RQmIH8ITwmk3keSB6tF8Hrayulp0QS/picyC1dB3//zUtzOD4eZlOs+0SAf9
dEljCTWO8s+MzqmbSb5z03vvr2E+mr2WMMUI0kAHDXZN5i16EK229W/wNhC8
lMMYhnf1Qu9DsufjnYicqo1dFtDkbXfnMKgrrCSYVQpsDwYl33LHdm4F7dd/
N+rAggLSVp/gWju/TS0dlXden3vVZO5HoOWTegcbGomYqy/nxs2iLcFIAmET
+shHMa4uiche9L7rvhI9FpQw8N8D7aUg0elqmriuLIgeIt9Lit6ic3FY6Kw0
4puedfWSkj7KvOlJ539Gr9j1VktkoWWKOhqq7sUGBBy5rqpU6CszyikbMl4F
fbCuW3Ch6M/aN0SR01kUarpJO8YdJveU4O2VinRGHxUl0fCrZPa7NqdhxZcU
70E5iUZCfpqaLm8HuwuyuNsllw9aQFL24Qsa8rCmpbdgxa5rPqyGn1q8bIxH
4ELs1gaJJdH76pGVqdK1bodrrEyla7r0ZoGzQ4cV2vSGGLWBlnBdFVUN8p7B
iDTczPOyYFxIzJH5DhB6KRQVBj6ScXmec75B5gSXDfnI+/dqe7xcOKB9qHNg
L4pL9hFdL/MWR9nhbWXoDHQVG/CGGa2NSGDY6q4gScqLW1Ecsap/Et/Hdu2b
eTEAo80KUTcEXl6GuBijHR3VdMgezjpYkjBTqcFM+Qf50W87Jht3XJjXEqNA
L/dRPrHR3G0/vIJCVe64vGF4wccrsFYBTqw4cDImJe3FTlK+jv27vA09zwiQ
svIfYpNKqpg4GjTyGb2mUCAy9TLt2Uw77VbDvPl2eZy9D9MBgSo4iORD1jM/
CowJ30g7iXY1qglb1iAD/nJsJmVuHtEzK7g7db5VgkbgpZg6fnIbd7+Mk/kz
nUEdQNONsQGHRwqh8IGJ09HTcmoewKdNewoWTXUtS5RzqAbbtE2/KEtoyiLB
XfX5fy0FUFDtm95X/XWTppABjzKlW38OngXxfhhBLrF6vxn6IIAEGqKr4VlW
8AxoI9VMrG1kMttK0U+9FhkFUZfGkdR1E/aUFPIsdU/6QjW0X9wXbBQo7H8Y
Fgkh2l4me+ZWARPFszjbFr626eeA+jNQ5mKcmi3b2YXdzuUtl4F8id+sh3P6
smTLwYIzAaAoU7YjrzSQkbQH2wBwHdt3r0Ne5SIm6iGWCsD14wc2uEFpQQwQ
kO6bMAtWVUpOwBPXx9csRgw5F58tNkrEZBuisSHeOYmTN74kyUsY7KMeyvk9
s6efE+3fy5PprOhmHgJymyx+2jfZe4weBGl5ordo8cfLFq8neEMI79eznY/t
hNKLackmEn+vXPk7A8e5/xCUQKL6sNl1iUQ4muRRZkVEDfJgwKCrr99iatEh
KxcSWglzPLc2ZDeaU0FjrnmF4nAIU9KpxUbaDo4F+BTzOreom1eALitDN636
JnpQSqalmoljcya6jV9iMUipZTBB+j+pJCPADD4dUGMi/EbwMky58RUcs+za
V9cvV7k2kaUsUOnHIX4wf9hel/qLBx1O6bgGhQ15xcaZbZYNcYBny+gY97i3
owy2KrT0sTFbi4f28rKs79EOpRK6uDDtOo4po1RJcvxSNVcUKZu8+e8l4bK6
t8ae7OylCThWG9DNpBclHC6HalrsFZFZqgP+IGvJaVQtvB0fCALq/F0blxW2
6rJ8m6D8ckMP/SF+P4Q+FJM2xzD2sXPi3Ray++SkgH7p/Jvr8F3xqXjFCZw9
isF72KKlLZZUp+VG25UZGSInnAsK3yUxNOURGtcB7F5pA0g1jp59VL5K7Hsz
v8HuA/jYl6lvvEG0Lg5bvg7hL4mJQCi0Eu7YQxSvSSWuT7plU/G7MoB+872c
CV7LLG2AJDHorutWDSkOcP1z+ulFRVMf4WKtvHSg68HDxL3E7QUWEPEev+iD
mvta+8B0TA5YLl9YjhjYlLn+HJQ8O1LYR0wZYIWcZex10L7drj9VlRD9VeE5
xBIAwvyLdRt7PADTHcMwdpDW2sIDrC9POcMr1U89vbhx/ZxluoQEaJKC0MXR
yHI5ILaM7xwwg5zG2+5pKVCwSx/BF/XrKOCH77LaHOVQO7lyyDYc1hn/AV71
gcHwaBy9kxSe3zMXvNgYXeKR3awpa8dRnUgDlBD6v4SOZcMFh5Sc3ytIn8h+
U21UPFyeYpD2gcR+K2wxsvRjP87XQxqniEYC4GBjTWaPrUQmNEdB2idi7tLl
K4vnlcn2EW5qo46FHvKgrIigLKnatV4WG7JLq/FCGvrYRtNK1Z857Hq1RNeW
K/vsZv2xhUfl+xzLQkks2sXKSaBDRbJUV/jW12mEQd+ebbI7kEk5kQY42wDG
ih2GQMOeBYVkzpwwEoCNHP5Wl1902bPvzNQ3XfRwwVgPa9uGg/PkhvKZAfE2
2hT7stOyiaRpy+ec9kZCgoL2pVfmNWtbvVjO+hqiUb4IPJZ4Z/div/LZu9V+
B7KhBUaqPwVSW34l6+d1uHn/df72lENzuBRpZi/Nji6u9KoUTWfrKxBStRJq
uYPEripeXPd3rlVLu3/WtS2xDL6tpjBF8/xJAt5iYy2lXq7Ru5X0c3cFi67z
IKC83u9+xtmsGYnjdqMBe9nXyV0ZWWo/4jyWtyBRp4I6y6B7s2Q9npVoJIhU
B0hqoJ4xDoMcS4SCsmBE8ZKs4kNhavsAcC25HElKDoYcKeLzlJd25s+Fw1sX
dkhR4DxgreEV1zld4Fh/17d5IFD/8RfoYVGeFmW3pMdnxA7/PsnlF0dLfOXB
Cj/Z+OrSLRnS5O6oM7YL5GcqAN2qAIj+6d1Y8GjNak9WxsnhfWGL6rxSHaSJ
2LJ0w0hNUEowmg1qRtWwtJ1EQFDbtRYE7L6ru5KUZ6AwFhI3+Ny04CQ3Pf0B
NN4IhfrtkcteJVN7LdMgVNpkGHQbPrc/I/nBzpBpWQiixWBQikvSsOUChzlq
Y1HUMcHgSDyaIQCiNJZjkhL5XtZJfIfM/b+5zdcuCcebJFZcopWSY3+6Fsr8
7YetSbEIcWwQTyELGqkaPeQiGq/v0lPoPrbugHGcZJbVcyaROlsZktEmd36A
P5pYREFkU4aA5Cf53lSTzKVe5ODFHy7xL1lOUWp2Miz1Xzu8zGWFi+Byopxa
mDNprb/S/C2mMz2nIH5wBkdn4sIvtcR+JiDCWD8KjDpxkS4bIw5fxvmes7E8
IdWiBZZc7VAM61WyIjl1o72Rfjsr1iIbhJX4B11gQrhB1HCOnP3tGzhjZaFr
ieoDqhqBFC/175RP0256mbzBHf74fXpxan5j2M0QOu+OapGfjAdz3qzi2Y3e
QMcGIxDNgrEYDEI2vmoObnJYAIyOAFtMzta4nPDs3tJ59fZ5vUmFz56EPkyx
0/jZ4BSurLYKWBzbpFxQSrTpHlgq2GRHuvKDlzQPX3dWyiDWRVxm3iTkyTis
/sxGxh2GEJgWxJnLuXiYPiWbjKtST7uHumdKcef3AUBQl7KJZ4d73SnkqlWE
72iBKCUE4KEXbgN8paVa8p+agpmBhLvdwGM2VMjbUmna0+7ne3349me/45nR
Erp80ClPSw8EizrUL+Dj6t9AKYv7pJ5DitNGThzBAJ265D8WIhPLMmhLncD1
CaWmDSvzd+baWic3Gi4CcHzmV2j+1tUyiL/QfH7sABcJeJxS6V7EoAC4fOmB
G3rdM1Hre4CBq071Ez29wopwZltazOHEu8hw1cGZZM9c79Ws2KY2YrzCDIkO
B2yKoKV7v+hU9QatRtw21Gg6s99GqcYRJ/1BUMn1FUkeZ7cDKzw92PiXh6mh
iKsQYDDJBeGeCbOsObFbrz3DuXg6q3CCkzjmOpUnY6UIdcSmSDfrBh/QbsU4
1UZIcrkjUd6BzXq56pOeFnvHlD5hPzTPeUZ3oV0SYXLR+2V+y0/H18ury2cG
7aQHtMp3SMV6DeuqL3FqIcUfMDcIrx5Kw3on6A6PDzwhzx+aOEklS5/9Ym9B
zFZA5wZemHNMgBh88dDZGbDTIJfbjEnFXToDYlgaVRpee21dwQv97YE6UeUI
x9S7vPTRMD+trIsiBIo3vE2TGyCvcCzlRdXAW9Y4NUdR0Rm9MOuwNoXBCj4N
szvgAj0xiDtsf5w28S+1+UqzDK2uNljo4V/8MUvH0QsHRBC8Ne/4DawREC/4
jP49FVS78Z4xOuF1PXvUN85+rA0fApEw9V0E4Lwk7wKwCRadixdBkPvAfYcd
SX/SCuHLjGBR7dVwcXa/nCijEMUvZyONFif30xmrx8pbVuW2XuN10hvjEi4G
OOutcODcRUR5X0yhMSJAyy41DFYsypTKoTT8sA5L960WzGyO8cI+LauBuRPq
7J5z8NBPblSAnQ+FSxpxzfz5tcDChnZHW+5FYMXGoDil07Zu2C20LE/HLTxq
6U6iRhITxA+vk6IPi1zd5qj+mhAZYXFRLzmGU/o7jr6l6M4YgEJLUMgpK8GS
Kd6ZU6se4/J0ST+OdacsyQVbBPtyNiX6dxLr10cTercBzGvfjSn16/YS+Ndv
maJzVIjryXEjYVmcq8eGm7i+Wv1l/6N+C0RCZntpXjyUiBNDFbIUbncsZkoV
fa3IqdUT5WM3hW925eWkWEg6AYZbyr81YASexgiQmlRWEY40r2qdMxSM0axp
kgymChzK4RHShmkIeXl7j8fVvCzKlm4DTd3PpNBxVsVPyGQDoczf2N7sPNGs
k7g+n9hZNKx+15OdscN2DtvGcWV8KJR0TyTMuKqI15VzLsPEH42ePhxXq1zQ
9Q1Y/87/E8qzcYxEYP5Gwt8a8GZAmZuu0r7xilnqRRyxAXvfZAGmE8gexio2
ULcQy6h8CghKLCsorTbdl/n1+Y4gcq40UxZEA+9QZDb/zryjjI0AYoIdMDhQ
TjkcY7dfDLfwLz5lWnWIYxymYQ3g6OJ5nm44+j0nt2dejziHIeZJRwxLdal0
rPPZu1+yfOqI2tW94PPOEln7f8/3gyvM6ssBSYhrpLKGXo+9g7oKZ5ew8Lzq
9vwyGJgDN55mZilaTaRaTd9DlLo0gqHmqgoZAXBkm1BzANjt329eptKNpSYr
dtaKJhJJAr/JfbjZ0GGLzGsm0jO1ACVluRAqCvJXWwvJx57IqiHWmQDV1eiD
+vKQkBtHMwRXUAPNYd8Nq3VgvlWwT8sWDYlI3n3Ib3C7uDxY2haAPiizIB+Y
qAHU1022MIpGUc8PYCULl67qFeJf/G7GOhBZAj9gymYg4YVL0p3ApYwCQ/9w
GsLr+1ddYD2iyngqRWsKZgMrzwFyJEZj3pVcfqtwInaX/5V67RkX4mBp9N2p
SEXahWh/lwbdBpoFvmgvq37wD5GEPSXla5q9n0EYi+HyIY9UdB+W+oYPTBO9
8wE48tCk3/1/uyDNI+Qg46ysarO3C9yTQwgr4YLoCc7J3uJDduzDC4RHjkaf
egpDCF4BULU8s+Vc1AockgN9Pi3krghwmzpO2S6Le01RmE+RzKaECWUVsz5g
BJu6Ex7qiq+KptcJZmtq5xxCLr986nqSYcx3TgcPuMcV2rWn8fydV51yQUwR
zeQjaGcYPi8qXkc0i41B1q/6qHPAgxDgKHi0m0FWCe1UqGGf2A0/uwVuEjK2
yEMwqX7MO9EO969Bl8+g+dwx8aNOOGilb5GGUxsC04gsKF33VPQIpY4GgWrX
M6nc7toQR6kfZuBC0KQ7oQ89X8vSdIl5hV33zrLTBZY6UB9TxMo+Qf7jb18h
LIKPMwoyJgjpq9uUjIpsOCivZ8qiWHw+4wJMqtT69ddfcvNhmiepyUpfKrDl
zNzh6T1IqKchtWW6BTm7p7r+hC/EKO7vDwPpB0ExoGQekxM4P3aMzpgckZEj
GLsn9FUh8eP7buOMVmaSU50UEgSD6OwwDhXMG5RNMuY2rImqWeBG/99M3y7f
Rm2AW3EsempU0Z3EI5bKNoB8uSxHHdQrjVLj+88+QHq73PRK4mCYek2b2k/H
tgXOUsqtpXfw24AIH1dHGtdB2sqkLdmMt1eQbKlp6mLZiKQ7PIjnOcgqdjxE
kd92loB6l9jh3fPXArZg93C7uyW20rpYqRhtvS8FKEvrMefzNNwX6W8LZrFa
tm09kKOWqkQfwTu7uaYO7Yd+WSwSXX/lVWkzF2Num17zR6gPJRJoqRW1K7C7
zNWKUGBl0jTQKAmBJ/mLK0SCOcDwoUxFZ6DkvHgM1W4REVML/huHMln3YmWj
3LzgO+ko0rvcVP4f7EzVsUWmpf9xE6sEqgxncX+YX7UuVJLiesb+1jU0LwdV
CR5ANFx9Im1JCgW46TQOV6nlspj0Jg2DEPlDFc7JpaNCXosggYnTh7Uz/8lu
OaW3i0vIa8dLoQD17CRq9TfBjDjg+5Q4j9ehxR79IUw7rr9zyHagp+tR26SG
VL/KimbfavLxRhkTetqARHDsTMHF97rffSaPtBB5MeNBmxMR9R6Ss6JONeHy
67E0sddmXsjnxM3d2RzTeIh3jkORt4KP6b99PfxMtXvflm/mJodxpO9z9ilm
dGOicn/5ngKZxjW7kKhKezBOcLse5HsbU/hFHUCRaRHDJtjn14IkLCcPrmuf
JWyhx+1Zqe9ODqdLeWIzjMui2tzPcZ8pkDuQMfTJQaRaQhPjl4Vidur5HiMJ
rAStWY4Hf5pO99S2VAdVl2dq1oNdtkaqE+tx73PfFG/WE6OiNjO0qxoMS8LT
BSk07ekdwTT83hk1lX8vzAHQDDUeRt9xPcPAoQ2yYtOqAtT8SD/fdWQBbV4I
S/1YVr8cPN9ObIbVsEDxMjbcCpN+EoLdKdl6QxwB5jwfWZfLWRzFh+5EYPG3
soGzaNLC7x3iAMBSF7bu1ulKxfste065NaEoXhoh/NYByh5TJdO/EGk8ef6y
m42vCHt7hfnqAbuyY2asQtE8sByqIDihZX0ZyUiI/sY+THOoYwgm7nNFSfSO
+mea1kDiKronE+Rz6gB0gmhOlDYmswmtBfmv70iEM3iW2gn2YY2DTK2NrrAU
dJDb728g30wLfq66v80ncdCkirlWLzVSIdZIBgYYEoyKEnjHNXSkhsp2aX29
yqm+F4ERFP7mbZfTfdbgq/yxUej9qKRd+PF7bXQLjEMEkh5PpmDDNqN5Z/9b
GjlzqTagAB6bpj69uXESAuKZwRiDQkexZJoneDJ5WvgUUaD64sHoR0B5NhO4
HG/O0LR0uS63zgVU8IDxmfne+8p+0gJDXxm0jHudZWVjFgCMeXRQspveFz4U
7xAa6tuk1Lg+e3YyfQHqflZL7UsNuujyeTygT6bRwFK2+m5CPVLSZ/jRBN/G
6WVztQ0nOvHoS677ja+nAawUzx3EiChgdIHra5rX9vfEHjDJFP6ZA47IXP6g
FpDczt69bkxhWR+XrMx/UOVzfI/FjxZmN3/wVRAlCHvngtqx+i/Lwy4d1IuC
KjT1WfF/PBGNh6wNzDMZ4eFM9iFhQBvKA1JjnQGU6jtXoJv4FzA7gzqZiPGz
BV2knAv9inyOy8dua2G1u5zJZa+6Dm8tORdztlo0iDvvEHNKdEt6C+0GilhR
Lz1qEwcjkFO/ZOqKhf/e7TjNDyWcQhiPp6IauOXoCuHHFYa1Daz8SaSrmQLb
VpiOwsj1Tmej/grS1VOBFt5uyz7nDjldYFFibrl9Kqha4S6yipKq8jVeX/ti
8xNN4nYzC2vQ35phVPkNDq3R7DL7SSWDqT/X5YY7EjQfRtZ8CA+e6HANiOJA
RNrbfS3bX0cge6TY99DzZjhD1cab5vqJmH/aTv2CX6zP29krtW5k+tr6bvuf
7ZWg3FzluL3+84Cv0yAHXOYdEIOvjrgu57wVoq6KrDOc8wXG6E3AZS2Yyq1P
nPKvMTU8yJqXibNOq3gEHhMSFPzYfQ57yznCwpbqG/mREWVGfjoFfrfFvOGD
+ijoYCxvNdvpT9Vcs0jUhqFwOVkmqjCqm5wstGDda6FWeBIe4vjllVsma4J8
KTzSVGRYtxPl0rR8buNnpCJFK6QMZzyUiheLX0gXPYt/cD1vJXcb8QAtCYp+
oT3hZd661kXiYUruFsRkedKKlPDZ8QEBdIP5NOHDicsim7qrhepV5UNi7m7M
ZiGCvxirN0keIaaf43qCRmDd4KTPIaJR3QwExrv0wWwnbZVOs9lmHZJDadgz
ku9n+sriwuzJDrg4bmHdzFx1kD3ry2+0EcTe930fbqgoX1XTEQKZvQjMqMHF
nrObvl81s0qRUodjqwXQ4YruiBOYEMpC48E1haSdhPjQRwlJCpbC3D/ss2A7
8YIpgLI+EOoX9E+ivTTxFsf5kWth5SdOKXmowO1kxLJSwMv5LPYsVxItSSCk
gTRTQWK/470KH/rA0njh6mSX3ccQM7HOGb8ZzAxrn1T5gaLJGkI004SQt8L4
FQMVcs7nxaQHwXpbwI9uBN7zf+K4gqWcUi99LS5pLpypzZv1zN0kgC/PczKV
e/K2Yoq/nvEXeMlOBSMelj7/Um7u6YyLCalwWYPfIWw/oivRNnLhYGpwzQBe
QVu+Xo40qZAFY9mKzgXyl9eMUTtHgX5dx24QgRoNNfvOC73FsUgslkgeDd2B
mqMyIbDIUi82Bn1Ce0kUy8NTQKnDUU3gzKe+8PLCXGt1/Gbp+mXm039nkZ0n
O0NvEKnA+h8wcFLB73IWUKaGQLaVbhtTtZ8bZtDz7ppM+YTd3hjRkX0erktw
MBW2RrLn/zOLr5OrBE3Oc/JRqrMJZmpGnZpcY7HNO3Ea7UKkDWzPgsx99b68
29uMQugY0kAl309hZx6ebA7b1CJbcJaU7ppJF5hPRyEzmrAp9opaFAvkaPum
a7suEhjdKsEeN30WYpdShKMMR0JUWbktlwsIapDTJrBqPAJkQYH117bq1ieT
/aZ5Hx8NlAX5VJw93zl+Rwdaei+cuRssSmxho4MUvk6e9Vt6qkbnQW7LC7R8
CB36lTk2cv1CbkrJRDQyhFkHtV3q9OjX7KgCd5fZoeIyFYAgwHOqNo3lewPg
OFMPa5Yn4yoK/zP8ITP04p2PdeO9mTK0s+N27H+GMgKzNQqwGkmtWpa2fAuD
9OnC7JiQ3NwqgBxOBKm3Q1c41UObnDM839eGij1Xzb6F1WcaSZiU1doTjAr5
X3GFQM6xGKJgsTIBQB3GshrufaDyHlQz7exfeFW9gpYpBoK/6+53QEa4Hgci
PnpBBJJZ6Or8YBV40H30ZJqZr3kaUgqdAISIA4LpiZzacS6ji0nhncfSPuMG
HSoANOZ5DJyhehkODuwgNGO7YMe5pEX4tRNPRurXSvifunpITnG5DZc37+pU
Ngj6to8lXUwJXViITS3K8DlnUtklewJ0zU+xfS21imHFGGbLA/Sa2etqpB26
IKYVMUDnx7aJaAKfqkcFx6rpvcPkMZjsFIrx9ezH+iWiebbUt96mQGJhrPMk
6eoXBuhe/hsnyhc/6OMj2C44Uru4UWLHDyoTlQkKudmeaw4XSR8Wu+ttR40i
1MIQsdU9kpmtHUL+9gY3RHL4hRdtuhLv4jVNkkUsMIuiJZxGa6LHEZ6daq/m
7/8mclM+YrGQXVzdFbkhS35cKVJubjyvoKPV85tyknn4Uu4ipbBm53XZLmuO
wFpAxNbFtVGF09F8Nyf6du6jRneX0ZaYsOfGdeUmpZlRHIsPwQtLQe5CKuG7
AcNPJRWjA7L3aUyPJaE3LEcGufv3pFUvOU1QxkXaIrUV/kvJf9W8I71c3u+f
KVaH/k2gkW2FkIptB+3mpulVqBxwAgwOiU7L4dwuOodg+B8YGs1HZ6M3Mffd
UjDpcHLQVL52OYJcEC5cy0oOblpnF8uX/geCwCZIscR584WAxdwL4MioiR9c
V8/o6/Don0as0QYjukb4+FMecbdNS7Pr6Y5wvM2WF/BStIXzpXk6IPj75Rs4
BBxVVVhyqEshWYEgnAPQwNQW9bFtSY8RtK8kCI/h8GuxruflrXoqaeNWDU/Q
D9TKYv+IDBCosytE/sS2Hb+UlsPZdzg0nuLzBy3RDD6oQj06aJhvmalPGcYj
6+5nTYVyMpfCINv6wkxRW/YdsYVtBDvthkGxqEfHYaTRaXqgUdx/9QlYHWu4
Wfm89C5ws13lT1nRkl2bpxnpty+GozNFPunPfJ3yotuZc3TJ8WeLFupWo+jW
dCiOiLKGKP2ZuYWuJp5D6/C7HgB0gRKxyRQmhx3LhqLXRtsEgasKJC9kIenP
Ti97PhTU+MRGJqIU6wD4sXZLM2cvywOhGSTe+XM7D1g4D8VFv4d+JoS0CCTF
pvbQNAxnAuBrWHZC7ZqaKlqvntaK0E8g1BMsaiiLQLhcg2hv8GXc0V9fvQmd
8lmga6k2dvhYHdbtj9MzHowCPCBEIYFxY/+mJqGUhdRCpKGVDdLZ0MurZl4n
I7Owx00cp7QctMzZ+Bd5O+TNZAisorcowztEFEZMxmDVZHabFhdu4qPQPiWv
xXLrNrDT2zXBhxc26yB4A4bHDf5iEN0Mkq2zKfq57P20q3sNLFJdjMEcEUG5
YUpXKdzEE0v6t9pkQZHBbEYRCgyYvAaLDgwnIiJXIhKwJfZcHut7zP1ptQsP
Tjp2sWs9XAYautLgukgv8BftkmkB9k5MTnLLRFZOVHvVSQHDqArz5I6pm4A4
KkJkyhg9MxtZ87u67qb1ISadb7J7HWhQGn5EesVLy8V++qXhkfdY8ISWA64t
HaoCelDwvg0NGN6ZI9bHu2A5IaZWCKitNeo7PLCA5kXo4WFr9NtVrsQuEIPh
jcaMe6h1yhV5VMbm/2M6Zh1xaqWsGGlLPmAjc7Jgnk8lNBRE232/bWaS5gwW
8EWWGPg8OFTkAqxTRBxd1RlJKy8M2UXWXuf5X84F0AWBPYgJ8/gyw8ccVJIH
KXjFo1ljM/bDJg2yETt2z0p21uef4htUfdGulUE5Ve7dYa1eaH9vvu2V5P5W
279Gcw+Ol/dnpCLZ6uPwIWZSgjhGYn1r+OtJKGScotkSEdlModee7dhMrq9N
qUfhnUCksHyPombcWiGEBN34WDh2R1/qqLATYYLSURig9EtzXDLJyeo0FILk
Q3kZw5ZnmDhoTPib7aOK0Ug6+JFS8Umc6nmSR0J/C8WE/KHz5pOwVqYiz6ZM
QiLldlwQOBsTbhi1PaTtm/fT5VevkHUDzyDCCQNvbgrfFylcH0NTUrCh2012
whsg3dKiMl6hOYF9INLV3CaHTi31pEBflY4Dr7SvE+3S4/PA564BHBN2Vd99
7TmdKV6Sms8FYF6UDRft5u513V3uOwrs+37I9xgXqoiDOLkPs7uN8QmiyxZF
6CxCVVZOh2FIwcyQ2OBiMdrF8p1yIjVqQxWVvcB/QLyqGbZjdrEep3oiPAM9
EtOVbYjQ4y8AH7S2ZqNajIG+rpfqcdjIuLqK+hJ56xOKbNdjmFJ217WhmcWR
Y/9Bog8VCavoWoPeb+xvma9AmtY3qiS0CryoKsPGgvtOeAjJEgnrngLPmIOr
qcuV+B6D2/MOThkRJ3TLMUyslOOQdtx4QxdHlDcuHzwdNFCbVkk25I+VkWZW
gHd3TQUhHLP+SZfDcD5I/tFeTEk+bXAp6rSPx/6j6Y1KkNlrJGtXIfZceWHJ
Z60eamoRSKLATQgrfxTLiGxZhOQSn2Z7cVJ6Qmeh7sr2SpS3zqjvdmJJbJvG
+mXCnvDftSbJk5IQ+snZSR7tQ49zYTN1qGPFVtU9GZjpfGMfzVqA7BL8Yb+2
CgJUum6SUKBmmAynzUGumkEboQBr/q9hgV+bSWJBEXY5BvXN0Y2WH2F4z3n1
VFjfQVlg0j95f6VfclJYQASrLsftEUHgRSrkh6fRrVAToNoV3i8SLVKLA4Of
MLAocQ1LeZbEmmRt9bH0ALN/Oy4FU3er9lCVFhgQtVsOs+JSYNxK0tB2ugoo
niEDjw2iVx6I/uSZwna9FpCVvmeGTbIYSmAKEzxEB0EEVE7CmQ49pIG9PQM8
hQFkKiThgsxZKavj8E7NepcCqmhBop586d86qIUn4BTqWJIWyWfCCjVYOieh
thx9DxzSDTiAHTvLpSQnyC9pEiadNVZuOrl73Rtv69F2LfVJo5N8iUz2WN9R
KqBc+prSYbwuC35o8uzg7rZvUpV126XifFubOowXv6OAKie2B88ozteG/QvA
sPPQapkJvafgxgxO+j5pFfhaqxNzsq3G68QVN+tir2WwmT0kx7ndNG0mle4g
Prtdx66FjGjKD6ImynKflvMFZji+t1CBX2OVn27SA08S/FNm2W+ixmtO+YWP
T+tTTqJbHBRjgEytAKm2kc6Kk2wz9q6nYoVB/YKl36a3hLvfEh4QgO2FXoFO
5myLlIGeEMRDLAzvvRtQIcZTOOzcQuL9VEQLalKkuEN568eBimn7tUTaoP8Q
Ce/ZkfMp5napeo6XdM5aosArk38dZp/bUkJg2HaLd7MUV7qi7Kaq5RxrkQCw
deCjWQSI2SX3l5pSDqCPFu9klV2N9JKXd8btEvM8+2YGFlrjlFLMNO9gzJc2
4OqySPgg2jDfFh2o3coGqpPAvLOywAyPXKKSLAbkq2a4u2nYN2ICq+7LTFh0
BGkDs+cDPqlLVHko3vTSZXipa+eCDdoKE4bqL08B5PCBRgzAYwqAtIsoY9ks
lZmXZApxEv5CkBwaAgowBf26CX/Du/wrdbHyMFeikmRxssuX1SNsVsqYkjnq
Vv5q0ftuC/dkCxiYKm+2PJFW4Z+3n1yOXldwl6WnJ3KxMIt6x+2A6P19Ao0e
MOe5kyUEinXYya9CfY1JPHmZ/3IvG4XmCq+UGJjE2v7r3stO9n1SReftDb2O
ak1TJbrIFXT9kaWGkTnItx97CbfT1FWKFCgFcrivQ9Ovqjt6qYBS2ICTpAIh
ZBNShcuCzb8kfhHYGHdZJEZ5N/MYnVOCDhESXrDLdYesXLpZA5DvLA6kvH2m
vlydjO46YjtAyaVQmgOsY+ocwbQjSsIt2tF+MyLHQC3c4WUc7GkEeTDbC7TV
gochV/3VoUT8VdAfR1MWh5cUVyAc6bY7MRfMiwMuk/sZmpzR6kkok8yywJ2X
AEocfooRyYVGDf594b5qDpuORsjdXfS5J9PthsP9GnnNT2X+PksSRsOr58bq
Gtk+2tistdZt1YGfuQNsOU/bJ0uxEcegzXJngHa25MscU1RH3yRTsD7nn8Pg
y1y515j8z5niYufJ//bnRtHLr+iWEiT4AAcFGibuxWWLYw523lqFO5G5Nq1p
n4wosdSqi4gFlVvgKuw8CNwPsiw8HUjTET2nnJcjzPH5nTiPlIbpC299MiBv
13cGhrIxRieva0si6a/5Qu0B6yBYaweyIflflAWPrAuHrU23c4s/LchuCc9L
lvNNeN+xPVFHFYqh6xo+0rzxGKDUBKAcWZlSwnEMqY2sC++vWHbzZfLRGBsp
+EyhEA3J9XeHL9pCEt9PnuWz/z+MN+pJP+EB5H5bpvdlU2uNrp/71LC6Sv3n
bqeNL9iaf6rzBQ0rCsK6CWmp4cnNNXVtM4KjX3VB+hCFVeIRAtz5CLaK3qNk
gvdcL31F/4VkZhsb0g541Lbl5jcve6RHrvTOsOA4qS0ipknM+hA/avEUmlUV
6LlAICXsb86kag6ngBzkNuFe8kvC9DDfczHmFyshuzxYLIzYHmDMJOr6uzDm
PlRr5fPPLyt/7W2JKBmfW8YPDbQvLP5LLLU1c8s6GCj4yRrEiCzXtYE+Q8uX
iSN3Rmd6NkuJvpOPhy2jIScweCYPxBMSAyo7f+owjS2i4lG9zLZcp2IOoW50
PupePV4J1zX81+0+B97AG0LTB02BEDXy8J5B7a/n+MTx0x6ljxLr8cf3GwYM
0EDvufptxjX8QESTmhhyVEtuevtBcixLvheJXQaGYjP0UFQElQu2tarZWW80
xPReTY9HhPq1egI5L6Uc2hT0Gspsc4GN7W9y7320TNtW85vRlkJV2bhIjS1X
Ko1qoSYZgACOckAFKFFdafrumvCWdlpt2VmP1lhRV1VquF91OFGYUJ2t2GRY
pAT9E7SAoOe40Ufv5MDFsxAHzU1He329OrqegA+CZF7yIbBi63j07uc3T4j9
nJ29qtKbeKC9EQ8OZe+BLduKELpbRmuOL24Ec7HUaudI2roOpjZKdN0k9N4d
eFoWm+3gyGf54JqMGvDwIKxKIBaPBTWc22EqQYI+vlSYAu4bnqNgMZxfPkZU
eD5gM10n9PI0IaEa7ecm4pro+FNxWcryxN8D5gfw0X7rVXc4+bunFWnj0Dam
wYzWJGn6z6DedomAc9hVYBNpbCSWOGG3QI10YfkEZHiv9rFjGamgLPTQUwAY
vZ71GCMUbfzRaEcgn5yinKT2C3BpeCPJYczidU/VbiaPVe3qHDuXopjw0fED
x0lIZdZY20MRwFXljJ1+bwyuAOzq+Vwma46FbhKkJeHnqHjMRIBBhjr+WZLH
vpBIjUONci13zZogRsbdw51woli4Vd4MA7x+Uk/OmtdKPbRGWK/NaT7n1VTQ
NUE0i/ynG6pebNyRS+61EHT0vIxwKRWtD37jgIebfbtfNYpuvtSMO5QnZc5t
r2DXvyJohYxViO8aKRc0nncQ0sIshhF6Nwia1F4hu2hjfcUEhRvwFJQqKhkU
h7pJyBb49teafVxnGCj2hdkubsZzrCdbFZE3eR63D3mizM57KqpTLE5wxt4I
L0Upw3zi3rQj6065/CbFzPqgGMoM2aE1a2fa6f6QWSPj6E9fTjxYewY/B42D
7o6pmo0aRbqyYTQp0GCQAOb5VDMacj6YRM8DslDvv9PjGewXt3bl0WzCCWeJ
6Meu/H7vhzSHS7hs05KpA2rUOQFQCIFq0FtNyGNaeuA6gAT6RVzw0TAMJTJ7
QFqqxte8ylRcwZ6nDbBmYQ2zjziCAHGyBEVf1jSAAc9beYsI7fp/VY/l19x7
EcacwLzWg3JPt80TVt806dDME2J8ESsK1iqwLwo8HkpHrAAgnzsqMZi22Bk/
qQokjIfKqaQkkjUF9Ryhkhwjac4feh87HLPhzL+4tR+O2/oEh4MgiXlyhV0R
M0gZS3+dmcJlZ5FbWmFsAs3r9PTbf4SYdOf+ExPJVemuguYR3HweH/S7ThnG
u1gZkDxYcZ0xNuCOd6sqCIbeA5TDEz9fYNaJPusTwmHK2YQtfDFaurFIyOsO
tw7m2dptXI/eGAo316nQHNo6ikbAYaPpBiC8R18h0dbhE5+UxNaJmaKLzqkU
Lft9hDWgefRjzqQ/1pBnWwYFqzoPZHvmKlobGSxZJgIq14gA8Le4X08C4cNJ
NZUsd0DXDqZDyFDuZpsNUsXQuuBghn4bScQOSk1Ig9Qllr1mEkBnFVQ/QQRr
TfuU0jvw3Jms5YMFPldjU6nNIfupcz3KOgsstnN5sCsYOcZimLufHn7Ol5fa
4IAAU7uIXKd9qTEfuzmv+otAtRIRNQqE4DcRjNChexamL+uKNHRndwNtt/4y
yB3aRz92y4wqG0sWs9O+aZlYQsiJpnEokYq/NZxsNpcBTO4gfiaKMUXxx4yS
h5yHciSR+2lao/Cm660bKNEHoN4ZsFkTqSivM+t3LNl9E9duvscocjYauUf2
Pr/sxzH9gWbKYM9kWjsYC2KDZagjY8ZAGnbsBUZtzPEB04RSHQ0lM6ZejJ+8
Grr0HMAmkv94Zo4Vsh7mrDGbMrWI0vVENKFQGla8DIsLHKfHYI68Y/bbqcYD
t6mMokbUx1rjQk/tRAhyIr/ug4rpsmuBr37ZoGlrVmf6XRLGDsHSpcSy6E5/
uLrRYYacHeLMMfylmwoGVLipJpx8PEd/ENghKh7druVU9egunaXLc3ggTFTF
h899/cinitDaZPabaajVM6u4y3lohXuGaFEOoYvp7yOzgfBZM9YpWdpBBIvI
dBn1yrBBzKt3oDBvFFnpgnZxWFDXduOhlNe2F6SxMtHwgFo4sKf03oUx+Zed
WkSAGQPQonOCcOkdrl+7LBycXUio8MlJHcYDFoiZzinpQDm6U6y7bfZZcpEN
0aoKH2OqmGBWr2ScQgYePLrExDKDxBxtcOxFyUjhW4o6FndqT3qY2dnxkFmn
sgwb/fn2WZ6kbtxnkJ0knhPWjzmijnFegqARJg3N89JF4IB6F9NPhM1rAOUb
/ADhU5aL4GznMBLuyJVP1IWm/pXAjuuMmADTG43dNTuttkeOW+EIeaGwIfNj
B0PFAuaDxTQ2D9yoggYGQ1ymUhEwmW11RG7jZ7irEmQyTdZASUWyaO2vj37b
fkc4cShukD9I3FBLm++nOtjoufYAdXtno1z6SH6mk3ya7P+qJbXo7B4DaQ2v
sNSv28GG62PRTLeDK1grrl2L+Uf7HSUhbNeRrk6rIEaIo1j+7vukHipJmYXw
TSpZhd+7r9RcvYVjmrmvWUoyrQFZRxcALonCOdMCnMX5lSANbOgNExy8GREJ
LDvEagMDaKeViIROKABsuLWa3q/l/q5Udav2GEHvSaCyhHeePyNnmY64nQye
xd43b+rAEqdouNYEhFVYx9OsiILw0ErpexJ0n/v6uX6TMhQi3FeFN1JtTc6s
UVBxwNDrDoFx4CqBOSd9EAq1PJQHXL19bpVKYitb0EeSbB8RZ9r+VxtdjPsF
RkcTxpeoB6Hjer2YkPHODNEA6ZZaqBpKc4qQ2dwPe9Wf3T/U6FuQHONqjVCT
QbIjJEjz3Skqlo+XW0fb5UbjwQ2WCXcRTeb/q+2Cpwkweu/2JiJt5vzsHruU
pO65TQq9tswTSI8Fswdrz6A7fJX2RhC11Zl/Ceu/IJ0YQjnjP2ClDVrB8TEN
mXmrdkdTC++pLBM2h5aDrw/1h5cm0KTnvXCkLYrJDW6hZcAJMCMgtghmYZUw
Fik+G0QYUVwhthOG8DR2YKaUghgbc3V54hbzz664eNy9IAYRJaxQiLrogfK4
LMjJPVk74JSkqsTKNw3ICxD7KmAnyVmRkUFCvDbd5YPfuthoIudRU0UjIiFi
8+iNo2blxq9jH5EidYu6vfM2/exxw3OlqN9t/1w8I7MCzkJ5zJhpPRA1HoDK
9fi4EWPKCfPDWloD6w3dI3yz2+FLpgu+4pda4QQnQQ3VLcLCq1DKE8I/mZJG
M/effk2EmK4pIusE/2/OMwQmUN9PSKRkRbtpz/ac0zT1+poxTuFMIICOLxYv
9F4aXmMGV3cPTc8BKEkati7r45Oz12Dj9nSCHbgGeCAwc/KytAkQPnM7U+zc
UlU0KPgMD4h4NnE9h6BlTQE8NsMpQz6JIfkvvEdDrWIfPKviAhnbjy7Y3kVI
DmkHNiOkKrcRnhQB124HX7dZJxcUc5YQyF22w6pghOnEF8jsoYTVQpaJOwjW
Js8Xa9Ye07Ic5tQKfrXBjtQo+5SFDLssDcq8SfqMn18w2xvrNldPiKkW/l4m
E7WJ3CU5+J561UVE3yKjJrPBf5Yp5wi+QbDkcHexBiNGayqpDIZPAa/ov9X4
Pu6iOMT97zgp5qkvANBv/GyHmXQT+rhhQ6HjTwa6g46HyHK/cLW+DJsu4MLk
+bM/aZgabJuTK9nxzmwNLugBsYWpmvIls+PQkX9sG9nfHUVOepcC+7gA90KP
lnRJUaEP+dnl9C8geHSzCxTtfLJkgjcBGUYPjSQLocYL9g/XAOTQ14XKaRiT
QEW5aLVOXtZDD74tvYBdC6C313H5grl/YCppZJMtHCJ/hq7Kd8JMlEc0HCVa
3aR6El4pY2RbOYjiok+ePJBgNOmYQKXv5Hxnxrnctm8+JIz7ZbydKLFt02LK
zfymdT6AvtksLT5DtSsIXgG0gUvEAUZBkv4kNnr0NGC1ICDyqQh1DBPiYt4T
nB2FITuPxmVLe6tii47d7zyGhvA22sDyXYaI+PXphOjYmVvueYXbWryLu4S5
71rONt0g95PtXV/wrWhZDf60GliQDhM5/IBNQb7fK22WSrWSE9Pu6WvJNfHs
0aGCOiXBIM8YwhNww68oEOciI7rJtt1vfUxBEP9kdZdFi6cPFSRNI7bGIN7n
HpbsW34VEth9wMqbrHCvVRPvoGGJqdR0emsj1KJGunsrkYFSsqze/da/rfWF
+dUBvKPvAuWm69nB+1sTxbhdO3N7XonmF7RjaOWEju2yRQVeVtMXrlkqrUaE
ZJikLwuh8ixsBcsQKzVVm81zRVX0ffMrcBE0cTAfwJh4wFDagvOH3peRUcF2
uKFcN/ksuNUYgu/rmnrBNU+ujJ8UwYQibKrd0KNWVhGrdVZrlnKhqc59r0SA
+qmUSodtcC5Bp4UDGNpvTIVAup+OICKD+efyQ+Ky9ZPpmox0eFc39i7Uk1zV
YlISBMB4dkjzOaKL2docCdcM7QDxKc20DRj1+mpBwUNEIqGmjxNzdd/v9Qxz
2TBVCZeQM3jpJ0H/ycFEG0a9TmKQ8JiSQ38lAKDW9QZlT4DnPyxm7gPfihpz
cdWGp2pZM5ceJT92/oQIJiixvrqgEkLHcPLwCC1KPqSVZ5E1WP9P0t6QxV9b
LVYqHfgJFU6LWsTQN20MJvzaiF0CT80aNXAzC0eAtUbLjOwRrPZrV+dpg5p2
4FL0HhBsHiwNI7eZmkx0xcPzo2l0Bnyauf0OxR8fLX+o56n5Zj7aJjJ15PaI
LhgJ/etttZr+ocGhdzvN7wuCJJjduSfhl3tpZWkwK3+8SY1G7Kfqji83XqiN
LNyThtDDYV0za2wKUlgX1DmLF3DjEkaylQWuh1VqlSKKSdxXBITO5PsCz6Lk
QXFUVZ1VT8wqtLFUZNu3DLEzwr+NHeDbBhCvBaVXHlxswc88VttrFHLsCdlN
bB/Ft50TA6JP05B8AMCAjWsAi9V3j+0iVrlugl/mnOkWEeLqqjLe/eBPhH2B
1eiWOQzPFGSIwywUCl12WAoNxaj698o8L2OnH6vLUUzT9Y8SF1vpl0GK+ys4
7XNJISVNYqUdxXV/38K+X1iCBnjIE//srKDPl+c/dZDvpDzs4RMRmMScM6Ve
YVfTUeoAuXHLgJywhDrOlcx4gy5h2UUJGQzGBEbsnxINaaIt+ACZU8yWM978
Zeuvcd0daL98KGtU5lBvktJdv5do5w9jhqQ+kstGtId3kSYmEz1UKxnCKhaQ
Lh0m58n8d8pEQVAMyq3oN+sNVH1hsgskjRjl6TqKVlGSI9QLwydj64A78DOE
PbzclKWz8o73dTg8lKefG+ETyqtF6hXZRifqQBzWunH2dRnCzUDdEmrjhInM
GfvzCejyIVEGorre21b9xQMkHyAlBk9EKayMOgwn7PWboSo+PkiZtsZHj4Pp
yA3yzRTAZ6OeOlFEivlnkcPjKtNvpH8jy+rxTB1ohK86sMoYmemcKwyL47SU
5lF9BmbHv+WhIE8XTOvb5eF7er8iwn34YOUYPK0hleXjJDLuayEAV/3LQYkv
f+O6ogLY+vwAkrxwYKd1Op9UlqPiTGM0KNxNoMIx1xsZ9kqZbqz0Rc66yz1L
jqlTIJzi1KRKrSj+i40y5gGOWb/otjO1NAgs1gTSBjIvY51zj8vX0xB0QJh5
+GabIYHsgIhQ5SwXO61xsQJCXhgipYJK0JZYXEy2HUq6cORdSH78ZoUwedQW
8HhTPaUFMoMaNfVgBPUjyrR6Ca1WYAjFH0b9gF6F1zttPxI5uFQfWDVhyfUx
K0q7SRixZubMnjr/y9c1v01PWLZZTJBUAB9ujHbFXU7MRzUYP+XfXXciZgOg
Pyx35EUnGvMLHorwBKvE8Jx8Cpic8O+nA7Hk2z24+7I8PXmEb50y8pj1J4SE
ALHp4rUVtQTOfLs3kbY5p4NxrauAXoBOY+/zwHEtjlCqQuJwUnJHiMv5KwiX
eAua3Y9tQJmEl0nQwXCu7XIMUjk1EQx+CsvyTEmpDB8joJWKa5wrl5rREjzn
/IvvBFiOADNOI1acMTLsXZde24Ngvz8lAstUPal2SpLCo/nvSf6WmJoqw2sN
AaDuUH9Gfi+jt9H+B3E2QGiABVSSRKMVDPffR1JO/KYIEWYV0uhAbQHrlL7/
KGBmTUxzE9mzMeBVCyHvPbRHbWxc2mPtC/ALpvjrRCMrjk7IL/XqIv5ExA5r
BeMtuPwpa1TKOIHgaGNRE73OFjaeQyX+jM/rPYNpz6yeoXHxZvqIDVb004cM
ohs7L6MjfFe7n2PK8eVEtvoln2GNn+K5oYi5EaxviN64SIPb/pocJmcqa0wY
JTnmijvMDVzw7VHtXqL+tkKV68MvKts632iM4ETmO3Z2grYWXlQSAph2Egen
Kh6unyQQDDIuzr0+NE2Hki5lEl0wYmMyV8CM3SuPb5n3lEkuBv5B6P2sd+mg
Fvttni/iBoqyrlBNToLSnSjXD/yM9UFs43I7ZpaQZwTJKDJwUv7pMcFLkCEW
W6TWlhg8oueKUylhe8nEpI0kMOrhFKrzv257czWWOxyeUJPMMBq8Z/BoPZ2i
RQiBRlvVq0SDAAhcl2/wgnHOJhgs1ntE1uOS7WGBC4DMjWl3fKvG1AeC9yOs
bgRElkK3tfLh3a3APaxR0+w0Q+mBvZZ5MF+x0WQzXEf5JMeCyYepIIs+OdLS
hqAPm6hxVB6lGlmUnGn0PeGNZBVvENRiQk0oHezCoKbmTgKebu+jzx2C6y8+
AX0eN/riCp65oi9S5JL7E3GA9y7O3tyIIfdXpjuptNP4EBbELmZPxGBU+k9Z
ENJIK9uBeXifdiFHa7aOSJ0o0jOWHXEAZBKNYvHRZN0vDeQGNON5QT3gSyTW
U6ZJN4vMp3mcvYDBFK/0j4gYaPAvL9iMMzXx3vWsFnOZtQhqj0zXy+Mp6W6y
GACQL6Qp7HhYG4OqbvPcHMOof0YhflX+GtubjCAkFh1NaezRv/6y5SosEycS
qyo347AftK66RpIdqzGPnQpIIkhTf88hfy3c3CvE5gnrZI4Fnhex/TJkGUPJ
6ngnWrpA3z0BdWIUeYcEom1n7UM/Mz37fgQK11xIvRKEXss+xG5EtgIoK36z
fMuXrAQr1/2UoeJbHt1O68iw66Rr+rzFCU6bQkzyDV1u7tVf6wXKs2ETQJyn
7lvYEf3MxWRSl5eaWyvW1vTSeSNlHVmPoKW4IVPbuy5Xt1emyoGhGHdhexVq
L5zPXbZYGJdB3B+9CAqP5F6jqZYRfCQusbee+e3/cuXiI+Vdmuno0zGvioGY
Ja4J5OTt78hFiDH8eLZb9HeSiH8DF2hI/Is1jfxLVpiYxQqA7vi+A96bJeaP
M3/GsRVnd0OfWd8CrLXOpgIPKKDpH97QFIHRYj4QTH9GxS/oSAgECIkUONwV
86ffv65vVX1oHdNqsbbSDu7VPHpJXL6EVpu8R9ZAEN3LXwwUEYqzNt03glip
6kkdlwNUi21fDMNpsAPPmGduN7TDG3MhpMWLS4yUJpK7is+DSmmxJig/rFvq
c9yDQLA9InQfGMdbJyiVwsl4WYHIP4qPglfiG4TgEQjJyhBtasiBdQnEJmDM
fIMOaIv2Aefm1Ao6rTOYvUqWjf5AAqeM7n5w9KDyghofvJHr9IAiGiip4wOn
docSiN1IvU7wEoJrQae/+1vZAxkM4si8ZHLEcj/6jOPWdqaNxQzKLzpHn75W
ZJ/foa9h24ML083L95bDzNhaY75g3RzXe0kRCH++pXYF/IvNBbWFwE9vbT6W
+QZ1TpRDYMfnij0JgWEbaWqttWUJEwoIu17XNlVsTDxfX7zXPZFchva6/Q5Y
7rAVtDaRMgLizdWNpMzTrUAIELPPllLstUVLZ3RMRF0B/Gw3Dvc8F1YqfvMq
Ie2evBPNqAlUVTw6gsK2pXr3O0hyfLRTeA5ELOBy3WPG3M8bjdsRNaAs167G
V3OlJsFYx7qgoW+C6vr1yYq0lFdIenD5lTvcaN4MHoj3fHQplUizYt+u5nT/
Qnv6Qyb8a+UNw8UMbFV61or5ASAQUs6z6OVzwIwdDcvxCydySygZNSDbreo6
C7XdYMXRGLH9TAjRUl3InVF+kaR6LsLsKJvwsHQXptjgbwq5e7hPmGQSoV7M
tJvIEd8sR7EBJ+znzuH1zaFfsxyQrfsvSQakpyCH+Dvm9ANKpLB85zEOeOmz
VMNPE/Kd4E7gRUHiVWxpcM7aTNRj5+Vvr7fS5W9NgF9j/q9jov/R2IFR6iTk
vMW/U+s1X+Z4S6y/OEqzd6H0dlavbMWMNFUifw9nAu3Ikd6aiQAuOf6R0XQy
420y/xxHYn1A2OfuznnJfn5quKy06GJzeWaYHxVng6e3t0DOxobD5itWTen1
OE1Q9jjFe8LLbMfjwuba2GKW0p2AETgzEoyhiu0w2Lzht/tThMzBI3YaHYz7
xYseBPUuygiiNKy2HYY+rcX+vr9eLBhcEK6269CIw0SrIURMnNFoaVNFDE+I
8SzGfEJfJtZ6EC5tCoPRMXvrXkP5ZaXdhs18KrXcPjpgp4JR/yVVmm5MJOWc
CKD667EfdUsL4JNNj4lsh890zoQPRfDRx9ywDQq7mTzZmxD2kZQDIDdEZdiu
R4ziqEF+x0IQDzDX/mVw+y7FcS3FDZJcdFCJLdL6iKrPtAl3vtwOLrC+ujtA
zDk/KvaN0GFmjzdvRGQY8EB3UH1dYlmNv+GCWNXePL1ZRVCkBrqiXek7X3bi
Mb7dkJZCB97eoIUZUWYfvR8EY4Zu6UDAU/Td4ddExQqN1EscOhbbYrG29x6l
aQiD+K8M3p97bnZDzDcs04JnFqJx6ZoXSIam1gQYjtpK4XWxSJ0Nxbim90XM
QmDSHty0BqQt3mk3gI9LjlsvfVHhZXD9GOlSlOG15SIbdxKN9hIaQiyl+Wqa
dfN+qcogoBEKZkrPiSa8fpVxOS2WJcXhA9JaOt4Q2lA+YAIfn8LEgeH4+2Ua
3lxSY6tcXTS3LauRBVTTOuexy8gwlaBJ5HGlJVxvfjg7hylGJb+ZnujUXKMB
pB4GGX9JzNZdeqhP9gwardWty+C1cHYs/oIpYvJWq2IHnqDHA00irSdHyr7B
yAe5ZltJjDR7U4xSqfn4yRuw5tEJw4wNI6uW6UD9idXz49//h/kdjbfDJkla
cLWqQPpXtr3sVEIGJMbleoLJ5xnHtu3wD27XR8n9xUbyYujuUFftdzPWNuyc
aySdrxdTor4enuko/+CqkhA5flmYAH96ZFY7fYlB5/oBnRU2ezKussdVDNBq
Cn0Tyqhb/VIV4kqTVXvQG731nPZJpikfV5CWnx7CadvfwGhA32lzVegPX+nw
UF3LWmP65dNoac7rNUuoG2xSWzXUU6+aCj/H1ZGJXplT6dWq7PKMuSNP5JgK
G4RctWm1dCoJP0Jl/MieDSXhWCOra19zXhozi6xqqJMA4qqC3iT+cKnfgzCF
oh3qeCq+Fz9WkrIIaLejgLA3jRo4lDiuZria5Vx64H7dOzdE6r64L49Ocnxs
VOpcaletka3bgQYdqz3WSjjA3jzEnU4ImROZVCH1KL8cCY/NlIx/Uw18SBNQ
Yvgnx+09TPFUpwSqtT1+o1s2+kkOtNihaBQNdldPcApw10IK0Xr7m5ZS5vsz
vN+ICuhZGzY5XrB761fMI3g+HhkymQCKDvTJs+BJrYMOcJaw4O2YzIvqwO1a
bMsDDUXu+pJyX2Et/vddIjW4KfRx2aHkoQz1ZXM33w0LU1Bk15FfuTRYFYYm
tM6db0D0qCcuWL8v3Rnt6faQIKE2yDGEnl7OtnFA044GREmEVdwYpNYfZ9wY
r+OCgnjUoyDXmTLytPLt0G+iYdsXQB6OpwgBgyULDJX5WoHMY5xw6Jq9nJWI
1T3ANNwKkNhXEJSzw7iWlJnBoZm5B/jhuvwLtuNmCV8CadkB7aXeGyQjwTnt
o5bKBf01THwlV5lFLCx9ZsbkBs8ykJMEZcXKgEtpID5Hi60Gfrpd+n3r1p4W
A42Gebt/730LyhjkLgwPcb0RUsM0MDlySNPdAXlQsXtxJR1Xj4Yf3bbtZSL7
N5wDOQTsl/8U9YMslv3H8nwbn9JYm6AgqKWMe4c7rE2aQDUV++9KLESJ2tSM
Gd396YbCSpTCDotntNQBTjP2mFkVO14ZnMMXkbMFNKW/suFRSxJX5wAHBSjS
w6zSOsD5wWwui4AitwVzqzSwHIICD4U/qF+rO2T1iBZ8hd/MaAYjL6jYzt00
W353O6Dw679VRzJ0NdsQuQjEsakiTGr+o1Kn/jSGTYz8GCYZW5M3egHGQvoJ
fTat+b5cFaw/erABDWWfadu7DS5ryBhl6znPjoSED0SlZc1G2FRTXJy3CQw/
qZLY8h6tnC5QKKsdrugr2WJMzqO+uu1WVTpSZVgxC0x0vgIucvd66Bb1pugj
TC2aQRoF3gPQS++SwG+xJP7KwtuTZ5o49Si1NUcAkzRNbI1atxUEjLe6uTAS
AHOqJi0g1X78PMQycIKm1daJFiqvP+nYLehgA6nwvKoIIcZHWYIvKDlYCTc8
CjDJ+IulmWbmo6gIYd4siMYCJ0xlNDDCZTtcgP9AOjJE69C4L2/RBxwJOjGr
oCb+JmbQGgs6uJ5g2l0hc/4+zBzO2DtcltSVviHEkqlVHcc5RJdHGEDQxrCk
/uN5Wn5kpt8KcgOKsMhJbPnu8Mz59Y+aQUThKTuM3sHbuRlClPcppYhuNcji
1AvsIuSiRjnU8Ts/lLDDAPVz3c4AAiQKEYgnX1TpQzEj6JcKm9d559GLpbGq
GVEwmBhnXVUvVFy4fFpEMCpRvVbxgKWw8mH036OlAtPIJns9rB4ZN6yxbnT5
3m9xq8+G8bxqe4EN++w4xgdizEwyqj6NwZmKAOh8MjSKNQthYhNtDZZTYvG5
wiBbPpGZV5Uk2deRKeDEBww17+KLMbmaRC5qluXaj9SVxRgqxxJaUJNYwYwY
0Z2dPbqsIY9AjFFdJA/t7EmA1pTWsIczOGFg76hFlDHdQhmoqQdofpeK7bMy
84yxZrq0lVJWx21lTWW+Y/zgjSj9OLwpR8iAoG0jK6PSzdl1+EmgvDgOSLUV
sLUifSLiYejJPj2XUeTQ3jvI20NW9TMBM3tyr0Kq07Seh0W1utCPCBxGEr84
9zJEZ8gF92iMlp5MtYzo9I4522o2GpbVmEkLzhmChUl6nUmRC58Wi6qz7csQ
4HFKj9IWXlHUmJe8jradaYDEUIYk6rHJNScsDg7giKOBb5sp3CN4a2WxXFbr
ho3f+omcIdLJf+f+V6NNxwyzbeg7NZTkd2Rut+dJbF2s+anzLACGlO7qopBR
bWokwV74b6FJLVZ7O+7Qw9n7s6nIgLGnoldQnaNMRqYe/VFisTh33n++ORPr
jg0mQjNWIScABZip0P3PZvfCylPxQT6IkGwqbTFb+KZzdTcbNEzvIhli4a59
Vg394MNB5KdcMTmTFVc/ARepkAe3QQ6nuselfdSOhZe8JZTLmktTzGZxE1P1
FH3uQnI5lAeqyPYp3YPBgc212C/1zipbd6KQ8Zsxo4S8T57P53jAC/P5Ap70
zOavA+0EfQeKfe/IGN6yqthY5LeyH2eots+gwjtP0TvNKGFkpTE1bwGIuCfR
I0K4Xi7EDGSmwOV/QacMDC+BvcZmHOflFvvrZqf2y/uVfrfuGlN0VSkwsPtD
GYP+sOYx08c16SadB/uJwUa1nOhUUPmjAuEFXcBasx5Ylp2y8ldYssa4NiQ9
2FN6jYSLCwZugJWedkz6kSi7eszD48lLJDZWFu63yQiO0Mp3ynQjWnuI+BXr
T4FwPtjQCul+sNKt7NyAKjARGUQIdrEuF2WlfVs4geWbqGldw8+4bk8GsZCA
mz7NLsOm4NprwvGZnO8/p5pE2qD6i5tbDm4wMyvqitJ1Qlj//VKZ0hada5nk
qBXmIA8BLj1YNgtAQUBW/4sHJmHhiv65gKiusqm+Vkar5t5q0RCNfh2AJd1L
OWUGeqOtj/qNCcOLoEZlb/EpeaZ5it0a0IZDoKBgGAkZG8xz5pgf3NpOZASX
1spsITE+xuiicdstayrhxCJROn6N/086RIYd2zEdD1hcmnJLAetvHWm0+yR8
5vbXk3avknZMKqGuphHf6YkoQsrKsEc+2vt1D+agnGxurTlAJggZzekEPHMM
cw5Z1noa5RBocGIGSUXa1e0TNVRgDjd0KvpK3OwL1854hyu28iZDZ4+vlpC5
XH5ZMJ10S1LrVFFzQMZVQ+Bs7o/AwEyXLqogDPTN5r+eP/U7uBXPlX5cvuS6
3ZppVDx3SS28GTocRfe2YIOJ5Hr3n5/oxluSNFuiUEfctcyOmhZ+/zV1XeGT
WOu2gkElXQ6rQFI8Iy6Mw7XokRs5QJUCFRmJ5cGsKrONnhABH7tEvskGgvF7
77D9yY2wj8SCB4VX2I5Q81MzDbQwBnW4zeH7Esd9MoBQ0BZsmcRKY7cojAvS
XSMQ6xP1gGGDR1CUwYcT3rdk3Pf8Sn7ww3ydmuYoWtla1jJ12xJun7PrhmiS
k5aePGlhQGrBhnejB0n/yT9kGLS0Pq5Luypyk8rsBiUAxmTxbZlTs+DrmHlc
NkuxKUiJ9nl7NdMmeDOuouOdyEgQDzon5s+CnOf++Gay0YZhfSJ2jGBhvmUf
nLj+f2pothFQiofRfS8P2wrfzNpbuPr3wGpQKprwlHNxPi8VvXLYpISds5jh
mr6djUaBsUloTi8C57aiV0XyxIhav2JqdD5HD8bnrragT9eC6XpEYvswTjvq
98y8v3/6AvUZVzCfE6AIQPNLvZ+b0QoIOhwYSI28oj59gTkD4tBHDNhUrL1b
zdaG+x/Tv2/K+csFB5eHNFbhhJizEneilCV4fJpi+itZZH4JJTu6OU1V/2ms
5Dyb9ZII/pFsjjpQYddOzT6YxDe4S9KQyR5bPdNmbYwpX/3TXRoJQhHL9mTG
qIjJUcvwP4GBP075l4n4IA+n07gzXO4NYSB7JVAIw9VTxGTMryZjMiM7iKoB
EY5zg/PsQKK1uiePZMKrR9Zr9W2Q8IyISKpZeOz/0Db00mZEXovGljTN+Bhd
qGMC2R9tH/OJla+ijz+Zi47QLuJAExkGg4uEz1r6K2ZUqEI219CZ1pouqj+U
p0GS/Gmt107TMgw5ULP5UwZNrgepwHdV7ijwm/+N1gysGy0W7kjosm3Tj4Lb
L887Gi/cvbHWSpNlXVyslu+a2U2FbowEM+7JJADsUVz+4fH1ZM/DsXge/8Eq
KoEhGBqPwauSEZaD+gbwPQ3APmxMnxjWPAMyGQkssfi2wAllJ8+iOQuid9jN
REKoi+avCzo/ky78OO+nbVF6SE2xCUmbBaSAQLWP6bfkUQXAGnPIq34xcDh0
UB7F3yIZjqvNmNNC7jwGFMpBlagh79ac0DYRfT0F3vFNe/Yf9w9orVUro7Hh
xapC5fCviQEJTTbOAUhM1M/uVpRjutNjUJm03QfWMWxE2FAeJvGT3J2dgMau
UDCmHkXA6mG7SQAf6m3tpI0//l/ZGz5bXuwRHl570shzR7HSFLSiFIYkF1mO
yEyOA/us369/9sZ+1dGUY959lcj6lQIjF0m1agP+96R3KEAQBwVqDIe9kSHR
OXTdzKCjmHtJPxKzmqzBJBO9wS4fuHrLldgSnO4j2TQyM27dIIMmP9i0w2UQ
MiLSTvr5M1cWVnzpa+u75ZAFxPLKm8cMLiOzGkujRi1mQeccIXxkGqI03SL9
d7uICZsc9TraOQ3GB4Zb9LdV2YCFNVb3KUT+NnDnAsOAbXZThclMDBiJf9VJ
GdHh4Fp4Z4Io5P1AheIQz49LAggES9vnQTuED1/hISonrcVu1rJYM4RrCS7o
z2igqGaFaJR7GSqYJuJAPGh+KqrqK1RBoQ7aXU/o48INb5Zh759j8n5uO3D6
plCfKeOwuN4yoqsAjhJaOLssHhyCz79rEKzaZWu/jBDeWi4ozRa6iRyzj0rJ
KlRd3ExCBCoaZbYMtgoaMmAMuYsmWmtgaCOtYpI4/2E+h60yO05tNVNMd6jX
IbIRugMs84y/QO9fPLiRn0DgblKrkPhbTGUTH6D/X+GKus2t1LdBs2iNH8/I
8ac61OVE1axgoy0flQlJOZQkxZHSjjmw4ljVRBzM0HdVBQsiULBkpxiF+pmw
W4EikeQc2dVd5pmctzaG/WqOb5y4gUBATapMIh62Gl+Y07QE02bHQdIgfKP+
Qo5hH39OHcbNQvYBRCxg2lvAgpEzXAclW5hytoaFpNDA1mn5oIe/wmfH0OSL
0vfxB8Ntx0Sv2bZXf5aqZCe1YaD0LY60N/i/JcWZrzcn1wi0Bx6iHBTFeHhp
R7pdUC+KlGLMkLNlsbsLgZ1vVkOea2HSJJ+AbtKukOxhPR91/0OJXwpbwRkQ
O7C34qFd2SUnBU6ytBopRZuo15DdV/D4ovTAAPJjnDqhPr3Bn1IjAWT4CCPN
TIZ/wWgj/wLD7OaP2FfArbD+EZ4UsvFs16JdcMrXi3dwosWahckneAMhr/U3
CiZiBGEwRbpI3YFpqFH2a91X3QjMdx7zMUNtApW9+UbllZ4QPX9sn0wjlQIA
bJDD/vOLBspYt+M4t+2kY91Se9k/J0FpbzpaOcmd5B+PTpKxCIbNrPrJYRoK
0PfLJrlP4wBsMHeWnII0JoT9OZ/juppoTD2vkp7UvLznm5lO5z8ubwp+VkQQ
WhmfrqiEH8f6qqIbS/Z7vo3qAka3jOhgnstjQztCjhE+eHzHpMchA8CVVBro
+ag3pR/eeh3MAIQVbAhPFL3ObjuYl83mNaY1exct5bGyEyeZNExEJ35Rz5pW
7f82lVURuiiQd9EvFZiDIiam7U4tHZ9Y3QHPAm6OaPHBIlVOnSUTB1ehi9Wz
FkmE42xMnThY2hVT7dNKn/YzV6mTKjCXuQkSaOhPdf6QcVJq9ar3LxSexwE6
a8S9DA8phGpTc69O42yUN3ssDeAoLdJ93EJ/9cCB2FLZa3qV3HCcN/DO+/X6
j21BWKmlRoEaDzNw60Y8LQqx6vJ9KkBj9qXp0rmF9QRE0WysOkZqec7422jh
52X5Qtr+GGDSEEAJ8e2mt22qZNOal3yGbH3KIIfQFv6lUtj+EclLzLkxPhiV
TdOaQb8zL7ywNez24Bscg3Du/jvyZEn+Kh/sQFZ8GL3H3PN85g+VuxLJ/jlN
OuWAn2h9a337iJPpsQoqRE/7tyMQjR/0CioXILRS5CIEoAp4c2wpy0mNiHG+
62aQ7JbaazTLhOSgTZzsN+e8SroGiMAEEeVVBtj8Qk4QCPW5zO1Ldp+cCMQF
HY6AxDpW+L+UV30czXdq6SYn3s41UmBU/9qMceqa5WSDz6/7bTk9R7zl3ypC
AnhtMD4SvHWLUjGnZHfNEDrj0wh8RP8vt2sMbNNXhobern01xDy94F04QVMr
fGDuZV7AcEPJSkSHSuc/waeBLg+kCYxXiuuNJfri+3RgxahGvkmYqhl5r7vR
poR8Nb9X1d4hxkyfPRjZ0bpbJt8S0Wrn6NpYLfeyqZhFdXZb+gBiiFDv6Y0/
eveTgOrbzhObuZW+7C7www2YSRrbadyu7rgm8U9T1CiCehVGlXZ6uphFxaQh
5LbdoHgP80pm6imo3FlTcVqyzwCYoN1/v7O16Yu9UX4xYFoVi7jlJpy0G0eq
RNuYT+XmUmSeD8o5ByrZyuSrauH5Ckd8EqkJOpizbslfUe/wzpvUiDm47d9z
4AT4RSDqpNZGlrf6w2monLMPVgVGvTJrGpgvyZqXWJB/d3qunAaZ46EwDtbM
vKyiLVG+4AOM992qfE4b39XLUxVfMlrCKPFkRNYgcKyPX54SkDVgVp3JvGBk
eNn9fPMpXKycfNz6ZYeOu7SYqaPSziUQirvpp5b8+pBjeiMNZqkh//BFBfx6
eJZpDlCtBlBQy2kMUoCi/k1F9PCHI/RocNB4Icr5nGN59UguhSxPlrTMpuXm
NRzoAKRHjEPmtDFkEcXK9ANCimY0HKiHaJjWCGb/I6MBN4nzIsJN9GK3maBY
SRwXHp0apdQZxRRqD4007SJEwet9hjuimnDskoqniBmK/lQMN7TNM2Qqkh2q
Xy4eip5MSRRG1f1bff/NcfkrHkaSlKpDBw8YAaZjOWY1pn0oUGbIbv+6FIMf
BKB3biE5P9QtBt5RdZQVjHf1JtiKrNiIO63in1lK9MidvJB53sxMjNx6JMCk
qACk2ADxblaABrTJJXiks2CH8lBHpiecSTtxyL52d9yGJZXIFVzM/R5pzPIj
LZrq9BSvuaUSHjdG2oDhRxshIA0NAVn/xbbnWzR5BiZyPr2NVSjpg18sSUDo
BsrGuGwyYBMjuiKDUYD86n5khZncU5EmkuelNmtexyBFbPiHtXVFzgwHu8et
cQyB2P6NlvqUj1OJYsE1HVUngiS/f6957oGUppo/ssS18Ln8+GWN5wZF/WOj
R0D6zKpBNzGiWG9s/YKNy7SH6oHkG++Ta9ZSow/QsiUbKiP6Z7ADUNieZ/C/
/Kp7Ax4rb98FWjX+wFiBo1RGlhdQLsEZQVuj9EBnkGdTePYSuDy04l1nHwRq
JR1RQPlmlPdsB0aYcgha+8XgGv8wk7GJUs0cqkCgByMSNYiuVR/jguUyAoY4
9ZDudgJf9tzx+CrjWAT8/kAthYTOUCFEecfJ8biCOt/Fe+kJXSpsYp1IAEBn
X+xZIrkXE5vB7wTAI7YYCw7+9dchTr07XxBvZv8RVC8tICxdY77OIoaivSid
OAE3GNR36zk19n4USG8paRHJTeLa02xBlyztHKbyz66/XcW9MxfSET28RxN7
DaUrLeLSrTCpNE/Ew4iuGfNw3FVAft9zMjS6uXutagk9QWBHpQSfHlkYhY01
GNM6awvOTj/XVBH7SOXQhVWF6saSkkkJ4v5BpNAPGVdR2hXTUu/B8nj3jRtz
5knurc7y89aUZyXW2nJHHQAdlwNa2bQhtjfRSSlJLGrO8nzxBrmAfp2YNxa1
rMVKI1GKiZQ4iTPfs1k3yg0xOWsKsBYS4goTaEasacafqpZa+0bHcbig6e9U
fh0wDNpKx2+UmiDfL3FVnKmJvdANVify5cZDDHYXzz6ceypk6KBFOKS7SRr9
Cs16CnUtQHv2OvfPI8MX32j73sOXjo3IptzU/8jabpE8ixz3SMCJmw6r4OFO
RXvFqrBz5tMyFXsGFFTs+jzHvZRE7AK8l28h0SZIW99PQzT760y8whTYiCIT
g2uAB9zp2S2mIN/CvI8QX4KTtcSsREJR2ZArQcWNPYVRg/k+zWEix6Jy9bD3
FOipgCw2EOgHMzG+d5lUgIaKgO77IAG20bE3b4j1TROOWEPn2AxaNPBZsyPC
PjScj8XkcIC1EA7Wco0kZvhIW3kjnUW6KiGsu/dBiL0vWqsgjt5ZHkgIFdDS
NQ0PUnehSqquq3WgXbxmSMl9LzOBvZFPlxcpNWv+zHkT0SFo45xC5UERm/5g
G+1ebfbUpR2OMBhh2iwjQHIRksuD404akqczbH8RC9JOO10xrxdFIrbepRbb
RCwQUSU6WT++Bj/U/8/ouJwyw35G19ecRu9mMxcf6zhseKoLZyOya3unCXtf
KX0v+Qs87e3uoRuvExQQhKQV6HEjnjAjP2cGxInX4bwj2o8AzQflC7pES+VA
KiChI3PEfspeUxoU1lVPixfUN87Qjh4AXdjpy4fRj/TJAFPG+on87oI0Mcc5
IELbSpgkahfWNzhDzHJwrDSBd6Eg4wbV8zlKyXzqqwBPz8M6xW9HJ3kZB9sI
zq6sQzkm4uixkkHd4I1Y/scmb2D3eFikd+lIv7zo0u26GKBt6oUfm+4vnRVk
f8Qsj8pxquSRHde54TE4jh7kyJFkwQ3WlaN4mB5O0Yu9cz2qXQiW3CnCWkF6
6Nn/iHc2vH5ZkxDQqGyksCfGE+JGFsraYshyvExKtPWfuUdpOF06agA1BBDZ
Gf37Ec+tU9RgRz33SeAP5g5pMWkriZQDo6SgO5xQi7OCG/P/ZWLGamxmOKox
g+VVVvsC1FXPbhsG6A74PMXh+zwnPiCFUyyoVTEEP8udoEVSNL3WLSNUxnFZ
ufmLEsMIOwinx7UHqfWvvakO0wxQvaU2v0evrB8xsFwM9dWKPr5jm+5aLOQ0
2m7sMOpW1uQ/F6NucjGOiCd1+xnb6h86mtNG2ARo7PaFarfrfJVkOeWfzcUd
nUVUyNqw7gsYZz8nrY5f16KuS6Y6RmwXQ3MGdvTn+AJBrvN751C5WRtKQhCU
ayjDaH0FbFkHEfdWF3875s839Y9m/uJoIX7GLwixd3RuC5ogwzUADKwAHZTL
3tJTROJ8omBTEiG6H/4PjTSvirp2U2znCNN1SJUnCJqr6q36IpMFJyYdDZoU
ocqdIA/B/+byHU4mLf37bWZkLr5tYtItT3bDS5l8EC5lIDhuRTbMLEtPqQVx
+PXbIe6SM2urj8Hb2K0/vfxmKkvM6daUaykZF6ftxk/Ebv5iP+zXGmkEVeib
+rO4jAZQvnW2dMtV12QJ/n64iaifE3gV7FSsHyYUJjw8OljVg/Tq/ctBPmvq
sb0ClDtLOHrnwKZkedJ/alXCU7/VwsKc6AaJwFWuihFX5BF1Hzsx7upKCXOp
Lr5bDHLxtO1kFtHQFGaCkM9VnQVFOxa4q+s0RESHizw076esy3rfFixBiL9D
ZJvBeK6/0hgq/K5G4uvaBXtZ9ojSiHuli0MYIVzCHrPGuRIO5nNiWR0GpXe+
+I+UBPcfttGtpaGKGxy9dE7WRZYfPxpt8pgilvD/JBIy6gI5lEfj2FHtZ7t9
zxyJEwHWd8UCCcJLVy3rIxBJ89E3CdBh0HyRRAGFLln6FsHPQT4A4t9ziIZp
6/UwoQWSIOuYSr+hxsTeNo3Yz0L5vUlWigSo+l517iDgDB5FQPBmUGIpSvJA
6XCCzyb1ZivCWdRAb4R5HYjVj+fwBuNUTu4KhF42HcgXd8xMJQxQs77JaBpt
61ReFaoY5l2wUnMTd/jhSPUd3dzINVtjKM5xOvqsS1I17M1oIrrlIIbD4Bzq
YiuMZ3MU+lAGh0/tiBAeLPvLC0gHu002YdS8EXelZt6BUJYhyhifmWp8KCDV
932Z3fnNcYSBiH+nJ+oI/zKhElaa/sqiMK5IVhhRMQcYy3NsAGeHk1VVaGfl
e1uDwcA5RGKPTDoSXrtjPkMpVQ9cVV7MZmbF0aHjMrPx1QtLiAFpnXufUf1i
zyk8Bu6EgjegJVH1whptjGds9vShIdwL3wimcgBXjGGxJs8VbY+JV0D1oqVz
8o+yBrARJdcFKiiKMXwxJzIaqgduYt6jqPNvWKIm5QxdRwFw7qVsEtfJjL5J
gSMa8eoJ86VYrpLmh39lcuZwvDaMq1Yy5UH0Pq+7wzOaM8tJL4/x5avBwXeT
mN0CEn7l+XnBVm2Pag/XWV2k94nTwi5jOjQiwEYx+ZXju4hKChtHkLy3xMjy
rLHgDgBeBYLO6lt8Dvx/HTcPS3g7XjBP0uleI78230O5nWeMVXMQ3S6h+geA
LdmOMxiiKUWhDKOp6zRZGSuyg4pqcB37PX1DTMVbnPv2Z1WHZ6TuHPnVsVLX
gMqp3VYXuhcl8PmxVc7eBcKxUMEMdSEMrODZvrG0zudHEYmh6rnYqLljS/KK
inUPeqeruYgH1/AmRVANjCF1JqO52xt9jzge0hC92ACDnnSjeNbbA6Df9Yku
n92FwvqfCruKhGY6Zfj/VGVB1sqnnz5t2dAAJn5nMeVFyY6vPuymzsujwSTs
p/zQFITOoFfx/thDjo2w0goFZ/ltMkVuqrTs1rHX/HW98+PE946UbBZkSdFk
i3I7fnD7Vg5w5ASszppG3xLYm7pAGRTcJ/H6KVN2vRrFNyvV15q4G8LIzOZe
y0GMFTY7O+UCjSy2h0UuDJTRmIBN/7jJeK9OEtHPXavYHUrVDpa0v4QIqpGC
ytMRa+Kz0Hl4OtbHMB6kRBUQQrq9RgkVjGKb32Smj5IOT4GkYvl9d6NUHQew
Vux0DYogU748h7kkSBLTmOQ+Y/JKY+zJka9HBSx/eU+UEJTSHe3VN8kZBWtA
iWjf1r7X7mB/2qP4C97QEomnuU0fNhsT1mifJQPMjuiwcFVLGWcpF1Pvxnfg
P7j1SPxpZ5ZnwkShgRnMgUeyLf9isXVaKtRN0S+dJzOGRLY5dLm5c5P6bKQs
zA/rV7HQ0KBK826EfCrYKHvbixiGdRIRURrC9Xr0LfgfqU1yNmj7UXy64OwS
a3NO/90sDKP4QBf4ormmAkdIPz6o05PYPhO2yN9LJEvJwYT6iwkaznK/PeRz
W7DYNHpR470ucXfZn6BnhtkADozoqfQIGlEEyK0DIYL6Sq29NJmfWAOZv1uw
gb2H25vv9+ToDaugwMxaLXMZsg4IBYSKOMuEbfk4qV1aFWVbwbqYpBzDTI2h
V3Y3OxJvUFTIL87B26eHblrAj+cVRVn8Fm7a+UvxlZQf+Es1W3c8Rbqsqz7D
kUHlGI0OGd9x5UrxGFCCXZTp25gd0MYnMGLnunF6CaVbG29vy2rYh5ALIvWp
0aglEBnfhRfORltuW2GMQH+c6mnwS4lQGldmgQdlo36xdA/Fm8u/E2BZHQA1
LSrW9+Dm4esWFOllqhzI8eO3QQOw17/Kg2umgMQzjhUUCc897/ammIUpGTYC
FPwgMbvP8L2caio3CqUmGmaKUE6QNO1ByDT3sXeIw7TsLaFu36A+ItWrb8WF
TK7+z3UnAZ2k37LcfUMMQvJzoB1g/U4w4va5dXc1FtrgsmySVNzzX811Wpdf
DlpBQ/BH5X59CrUscMqO8WkthNeoA6h5So6kLJpfJqjIqQ4EV+Ft69uAh9Ki
qPgibfFz8SSz85E92yzQhzDy32UtmD2BzZZkRQu1tolSbBAjd5OdQZpP9qml
IeddwDgZ5gsxqDRl43gKEw3lsNDGQwF00DJ/vD7xZtUHHuZqijAOgZFR+uKp
W4gLZ1WAg8Y0yS6G+O8Ma29pZEELZYx5EVy2RgJ851T1m90MjFgSVqsipEap
U9XnSXrJMvrnp4cc6Hts1jiQ/HKeAzW8bb7CbHYGPx7YNHiKtXOICKUcQZxI
pjBhzyzdfsKXEYmPRDp5Qxuu3RxP+WlSInEdSfN/w2k7HLzU8RZ+IempVUL8
P3RjxaGthjAI00ktLoHo6InB9/zYVhnD9P+webHSP00fuE9wbVDy2QVgCEDe
DyLMwLZ0dlvTf6qAUvQylJ3HvzsjMtPy5KezrTyyy7trWj74n0n+NMnKB0wa
3GphQMU9UJXBb+FMrjz0qjR42f68UuXgHKM7Y3UNO1ijR7CefRC9ymt7Hu/g
bCaLpuo3Ss+xWQbeN4hdxUVZti0wKC7p4SzJ7zRYktt749BzbVCWrDHysOTx
651ZPvzASwYk9bhon4A1ER08WZoAk+64H/4sTiKYjQsJMvi6lBJa2QRByJvw
0VhqSMBt6oqR5zjUrHOKEBRCvMdQL7WTnqI1QEvDiKZBW9/Vsgm4rVvy2zBZ
B0A+mSmsceEPuhFGlWayhEVQQP9XA/ZPq1nveH1eHP+rgYnhrSL16h9qvVaP
j5IIcq9lm0Ss5hnQgJj3+zPV8/6VEhH8zGnAuT7oIR1uBT6fkajMplGFynQA
99H8uIIT/Aamx4gk9UjETxPJ2OcYimSfxyjL88arKSlhPAdrXNfJKN8saIqM
B1y4/oitN9wxgs57fYW/fjffsnlyZKzzDRYItVnyqlgtACQHVqxkdj73hTbx
DIhuw472GStKORFwTT2DsZbiXsbqq4NxmJBpmLWDIzciyRW5pLFaPENxVWwy
1dYgh+9quzE0v+VgCMP84Db8ay3Fb/ww67qytbEH/ad1Y6Nsv+/bDMg+R/tS
nulcLAPFvGMPA1msLc8WXJA9MbwqBzaVecyvgajSQZwFXP8pvZ9+T1Sc2XwE
HG1tM6VXkpKdZIxkwzKFHFBNZ7zQx9sSfoA/qm63ado/Vbi3tewZjq2vnfnb
pwWZB45Twsi15CuWihaNyLo0y8zPEnazcmK53PWMf6KXB72ssErsPJ8EMfRa
+VjoSYxGE7e/QRZvlSU3usymnHM6gEyL1Zm7FbHqEc4ntZTpIBuinPU7fa59
EqC3wKtXr+aJKDfXwmsueMzlcGzKv0MpJbuM22oQEZv4205pmsiVUC9wmWhN
Xh6Fj4uH9YhcKY4rdwTd97UgCrKBWl4siobK4Vt9x3wcwZKchiJBqKNuUxvp
WgGIlHTXwC8l8XkpxEPzASq3CmRT9rkICuA0oM+9fp2bCNKPjueTSQa8bJwM
//EEeOIzBc84+NFfVHTjnTar4MIj3zXPp/0nadorTDmLcFS1h2VdXDK1BIfz
0MvQbQ00/mN7FtFLC2VSXiBoVpyhmck/D+Z4826gCl4lNz3QJ2047Z9IuNga
DAILm194tLl8zddUInKi0CyDuNwP/2x4XtWf5BpA4hufmLF8Z4sNgmKl44JW
qnNPouYBf6mOMS8Sfg7M7kIH/8DYKfMgvQLQDKBYboWSUV3HrLiqedVQgRZg
BfeEc14jWWjfDJ4r+vbggJfZt898OW5pxbpGUNN1eudqAoCN+k+x6J9/CyJT
SMCU2eebNoFsGsS5JV/tIsgVvrGb4QDKNqyP9/R+AgcGERzTS7UkDKX8WRRu
lQkq+E0bZca8RYLF05PMngfjyXgeYQ3JhfRXgCMqKTebFvsxnEL4zIFf8JBP
puuwA9VooEMiFOORPhzd7g0OGJki6amwjVxSzUeEAy1BVodxnuzdpqyIFTew
6BMc2AsSD/0BE3/FJ/q5wisx/sR15tjggWZ/b5ZpqDM8RyAEX97Lm5ynjscJ
KWoUzr6pcI8QceHdEk9r+Y82hMEpRXOE88Lpe4J4amGRUlf9PIe/EyXnkIaH
+YNraCwMzouBSOBV+mSygm+8QJ8ltrfu+LGVtlzE3VsZmt1zch8eFb4ZHcWv
nGrijbFKzJnpdcRr7ELO27rJmCo+nB7esui9c5oFjmb08L7kfG1u274q5PwG
QLB5B1lTH178qfVOG+X2uCq566crO9710SIHjq6bpea1P1+HZtu28/0RJ/Bf
p/9O4yAT1BHYSYN55nlDVrXepNEFtca5Cu3gkJHmT4Dz+kp0QvJx5Qjyxhoy
k1dN9ynAS12tnlek01Zh/CVMhZtFV+Yhx4B7GDaot7ByzxUGefMV/xndcgGM
ivknIcbly2Sf0lQnlDs1H6alTvq0Ju5yMI93BAKgZhDHBH+GBB1mZOcP1JKK
3k4Y2UC4X1pGB5ZZP5vGV3UAwyNfhkeK0wWxbCWjdtkO1LS/bT4j/ElIVPKa
WJx1h6n/LNNaB7T2SBLk+y64/lv3BqErSg3Vc68Zg1mhxJL6F34okyEaUAnF
4GfVXrRKmBZPSPzSQffeeAD3fV+WuGlvMJF2+A//Ux9BzTppfG8/T48yH8vG
Gtoq2bcVJo+JqRncAygMv//opkWr9Pi3k5CBei3U7By6vQq942Buyqlt+yBr
s0iMGSb8CRFZZeOW9xdHEbU4JVemlbPBkyTKaJLNcEGRt1W4q1W0+6AWEo8E
toLD/OshyL6F26rJyG1+dccLiW3LrMD7LvnJw7dqrqvfQipDR/MDB4Gi2de3
zUHV6qcUy0slhBarTOUCNmURt2L/OBZXsFyXycqXVOH9olw28F/Hh22bkxVu
VeSfJ3/dGs0/gk76ciWFZchJFaovRJeI55Cf+gkVcZ3Qx+YxZ4EXb7ROq7uh
b0Qj/XrEaqT03FJqZRhSg/3wNgtDgEaZnf3k/kqCc52t9jACiizXL2MHD4Ln
obK1SnksR0X/1lGKiyDeMkmoOdC2tn7bPZu/slcDGgPUfb3n5MJcJYtyECVf
c/n6fobSMKc4aqpEuuzU5L2sxkZvNKmAQw1/L0kAoavnbYhW/pZ5+spuq3XJ
koPP9fw1VfHPNNzhgSqZr7yyK8iT+6YnXfcXgTS1Xp7JrZLoj7BTqedQbILq
d1Ln8JZjoFWZI0huhG5Iyv3Lf8gZV38LawI4yLP7hyDXk2TWuP2b6ucVHBGO
yd2TFR20e7MUiezO6B3eWiAZQ92dVlOR2DrwFLipciOKOWbUc9UTwMjjq/A7
CFbeAEvJOGXYMRr/2rf1vVlzVRYQczPgTe49w1ZeMl92NaNDpEETQocXi8Ha
FQQ7Vjmgw5FEK+hEejZ9aFXX9sLFyZtLBZCtV3azn08hMNX4xpf54iARDDNj
mw2AVHMGosnlVxnZRAB51z4pNpeUGpSzGKP86FYVp/TTz4/uQUWODfq89q+Y
WmPiF7a0O90mOPRosnKeU8QKxBWO1u+zGV3F5Byppk/oxCxgtxTkOxyh3Lpi
aAWPP0j4+lxSqnMDAWMpfHbW4eYmjaa63D6P7VJBdX+id3Hg12T0QIayx9JM
U3gHhHsOLDGPUO1YM6qAGI8uT9pP3ed0YbThbRkIQTkqfAtJrmvLlhx/9Ubi
edbyOuj4rmPnufvExoB93dXjgWJ2yLcSc7dNHm3dZ3RX5pUjA6I/vtas/cAZ
ppI++qahs2UXKjjJbfFMEdkSnPujGHzf9ZmfvysxKk7xe1XWee8QlHXAi9I6
mXVoBvGEWLXFkgoOHD6zz2G+z/ELDCbJJ7QxafQg9W5XYeJgjnqTjDYz5EuR
5P6KA3RlgB3bgq5bYweeGG+Q6JKAw2pEjEJZlSIhf8NomE+d4cRCIfmv991y
NFTmoZkUtKHkWh7eewqIBiN8sYxLyDZNg4MSwQfYvoLwGpjDy5mqPCR5pXDD
YJ47A9NTMgPH0j5q736aIz9tGM4dXykt1aVRAh+ifoZIrAeJDEBouD7w8JCD
Isg+sdRLLl1v5cMqtiC3C9gV2bjOUsZadyyoAY8cwFFDC9sUFdkAda4iag6G
WudDHo9GtzbGcVlXdnxRH7ccexDux/IvqGAou1+0sxuDNAqtplntyVRoKaPp
ogUslabiEuEhVT8xIhiRcsJpl4HYVinT313cEKc/5Glez3CQuYrA5RW2kWSM
jR2UYepO5ENbDle+mzWA4JdSeNcM1ZnODpXs17lQ0Byl12obfbSzvhgPN0bd
iSl6a5WfVyOFncRIK922KCl2Q3E1CcTGgZpcMw7ZvBb9gaN0cAIAR5RV5yeB
nVf6St80FHiGe43i6LjPrqwaCLEI0mUsJtkTfg5m0mHtGvpLdc/buOKx/nLk
6fo4eqLm2nUIjBbgzu0UjEeCZS+Ihp0nsgpSJhCe+mCeUQVFef25dr6A0ZKR
RhnSDTKt5e6oZQPtUdvfWYwBATllTZFhdyZ3phm/4IY6RH+jY6zw5MDiQfSD
sYHPg730dFrtJUlk+IeZXpkoaXU57T6+t5q5GK1O3nmSG4PLAaK4MyO3EewI
ngRhIx6Rghwk5MWgWUF4Vyh0F6heaXTH09HvHGthV+WVjTA5W5HGGcEDwix6
/tGttOjOykLRa+AT76CkES20YHY+h39pDvZNcNtvyBITy2Ks6ZYUf14HML9r
d9mg32aeWLXTG74dXQrngBXeBVMvNfNZvuqkTUrSwxTjQ57WVKdz+VRoqNUw
lQcZgmCz36ENQP9EucO9PrKUupvOGK8PSnRNxNIUzv74m7o3zh/1mEUo7rH1
zgQdrLDJFzWaBj7v1fle6nFpzpO5OOmjrbnwGSIvc4Z6jIW8i7ppBPXFy1eZ
1Jw2Pr51EJiVRU90XUUh9Wjgy/04M6gTYWq3v3C/89fb9F5zXJCD1R9lMsgP
J6x80qooqK7r6kFHSnF2FEyb50O+IawVWEVKixIKoOK8L01JnSloPSQ9rstF
m99v2GI64/bjWVC/xR1a7KkHc8WSgqMOBwrBXwaLZswqNgQmvSNlTsTVwZ24
BsatvDUl0vyMCYKd8/GgimM+TbtW/9qpvamrIWFDbxIFULZ1CrzXm3MH79as
A55K0oYCxbCVDNSYK6FecUbsuPWxCFEPCGQAeWFJaP5R47Ph0erQBMRrct5q
T2nb5ZYKfI0aqIcBlaJpvLuz0NoVhUY/urYxQ8UmtKWSwl7CyXHfBEqaHVqV
6fq9xKQvcX6DrtgZ5h4hbBQDFgs+IhUTfxcCw7Rdh1S14FQzbCtK/HnDKaaE
4hfKotSOv+M98gaFFlP0C5FdGjfGSoLgpY0o58UUh+rujVCDZbapY5HvLV33
jmTNqZimZfjKnHXw6helXdv0Zb8UuGoh+pl1Bqmb+iq6Gr1PL+SR7sWtEo4e
N4yMcA28IzDiKEijvxKlo9tKr2qNhvM0RVD/JZcqajT7e3ZDG3yELqOX90j1
pDBpl1P1JLs7oLoou6LRXwXK7lbw/aNTWGW4MDKUpGOP8J29nNxwjpJEUBCD
gRbmEXR9ZM2GRGMv0h4GmvB/eI45N1wld7ZWEPWWvV/kVBv1+N+2p7JpibU3
rjFDqgwtIB/QmfTwdV+symOjw2aYk23ny5ASrtqCPAipZ6RMk/vutCXSyHOK
iCNx+vt6eTxrlUea3087nMUzHyBCUhJdYJqCNBs4n5YOR6OU+YVH6YYIQ3Uf
lVjYHRV1geftb36y6nuFmBoQVgVpIMpJ+AGJ4RcfYveTlE+cIFW3se0HoLTl
sXliAVLUt292wLIN+h9wq4rBHMpaVCtXTn27ZKuqvOhMgwdlQFjQw/UHiMoQ
a+VzroRd2x3qx8mpwBIpTwIq3quNQ4XDZG+LV4MIvQX46tuNGQRmXtDNhmS7
1BS2V6kKGQtDVMmVKD6uxZ775bKH8bbllcdA5BCvmPeMmyg6ydi/PfR1lLmK
PdpiX7gLT47l3bMpELwDkI6DIftryD/KIiCWK4csc1vqFY03s6XlvfP5Hc7S
Tvtg+F7reIdB8tzMbPwiM9YEQwuQq4+8Z9nGF+w4M5AkVc8Z4Q97t33qgZYc
Rnd7qbHPMX3apzJmtskIH7O7OWsAduldXU38NJe+35rTwFv3Q6LR25Pltg8D
0Bc8QNqLvQ1o7Yc83KN7mnzFVBLAsA1veP3j8jNITeEd0sT7is/jZT3kfPIA
Tw64lQNgmpggl10ySHRVXc23jplikJUjUxcQGPnzOaFZZ36GAH5cXSq9k+hR
bDJMqflIAC36UPY9lL2M9DX8NyUJORN8xus7AtW8EmQJacmnYrYwwLqCHlTT
JLH5KDZWEFmCrK2IKTbwT0Mkj0RX9m5P9cu+f9xXaYzToOOIf9zGZ53Mi5M7
qER13ECyS5cM+YwFs1ujA+3QYPQ8BF0vt61XP9myIZUNglSpBl4Y7dNu7fO7
uaV/lJQNnEVn/btj2g25afv1fsWpsHVT067L0W5G0IzZKhlYUbKFXIPKieER
H4MzwjDpZ1qlMgqOuRNyoZWhvuPpMt115Ma6Qvo0HqNa0lQHGUG+PPo3pLCs
31NWdM6Jxq7YRhehvYiWwNyFLOTb5XP+kCt1yK9n2GjF/aHO3wcFAECYtoIY
S00DapEBzwu97iuv8Ix3GSZhBUFZ0FnGd0zMNvXLSEEx7LHItho8DfFmB0ia
6yuW9nSaiM3ozYJxo3P3NqcaB+yMUFjUJFZc9SN9UFYpiR08t0K6EKtPBrMn
YnGQ05XaulpZtznWMkUzWFYg+QHAjR0ZFNaQD8JngfCJ2fxdprjH9hgayeoU
sFIHaERZfdFBg4CUwipSa+XT8VJSkAQqgBtws9FYr5uza+0SVXFHIY0rQpxr
jeoODDIIPUeoRERW1nkmyOizNwy8UhX024uwXYZcX7L94pwTwse2iJPj2snc
kyiouU/Al4MHxJ2Cm0Majbwgw3mn2chvcAPjg7lnPKXHuiEXTc1Kyawwq//o
m505mZ0OMDnlrLE/c9YDjzUny9ZMzYELwEe6O/pLErSPAfD03jjj6mNcmu+G
DZMpHJy5Y+irEYH8Tu6yeCjpXtX6ts67wjLQzjiBYo/rKdqypENB/uF7VcWW
IE050bxkqsv82OZeG2owmPcx+pMvb1POZYI3XgUDIYcuAEWFkPs9xf6ezpp8
2/tj3e1X9FJ1Z1PbOImHIqKS6JFfralNmxss52qy1TbB83KVrP83NccaIMiD
5YiCM5UTXLEu6FGjuMsGrAfZg1DBGiQtr5G1+rC2rmeQsIFpexRS2b16u+KV
RZqLgldG9+r5nLbMecagM0qmoKJP4LQQC0EEnN6QyQXlGTG6flNpzlg2dgYT
w7RHCx8vHwBjS/h9fvHsmDwKqFIkPMs0fhlhGeA/TbDyQKKOpQtWfaLufoOi
m3mQj09FV9nNaAtbszgg5y7R70W/2ppwOM6VQZfIEaTexl3cK69yX50DyNLw
onf5ZCcHYpAKKhLzZHSqAjeWQVfbLdX1jzdCWaXWlCLKkqa3+9C+bNpWMVkJ
iPS354QnrsmJ2BvfSFALy2L6vbVI0QTzNmSHGrCeBN+NMrCxsuafNpA0gSW6
qkOJW5/tMh4OGFbqv2l924z+mXapucSh0ot4AFMv3kBY8pT0YJpNgbExLZZX
vpvilwk/eeQ1M4H5/wNFnCW8q32iCSfRiVPmBO0ZyxfAfoYN7DW3z27zlBuB
kRrp1vSbSc+O6z1/bt8AulvJMHryq1pSjxve+t/gXq2ewmMRuosyn55euqZA
vY4hvyIyslPq+aYSS/njjpuc+Y57MpSf4HJx+4Ey80ETi9VYyuy8bKGLPhKQ
6xtyzRfRjaY4nsMfp4eMY/9P1Qhi/NAKlaojfcZm2tq0i07coE5g3+OyQVru
X5/9zxPjoa31Ih7kBEEdf6H8Dj32nGRWpO7YkKTBAGguVs+zkT3f9cmSf646
2tF6aEdJEehS1RpBd8zp4FRUbxwZvUMXdLKAA7FXZhFvcUgG5rqSwSTP39nR
64cLKEQ7HDOrntPsJFe3F+k72sQArPoZPS7V6b3Sf9UtEuOOJhvcckQYpbC8
A6fZcZmI2T10V5J5m5rmIfQnO07CcfgwW9wjg3sOaExfZ7roHFF3cmcMELrp
dDBYA7ryaOvllrjS6/Mx11Yvy+JwvXMxQ9Nh8S2TElr6jfbCHVEKGz8nbjoJ
80ZYk0Q6L7/EyTHi1MT+8+T2iCTr5IcLX0QMa95REzC1fIeeWNHXzt+UrXH3
vkhDXHot6GZ8+OtCjJyahCbpIUCOsdnhk939g/6B4x8md7/8oiLfrfF94kAT
41IBz+jLOnrmmwOKHt/aDa6FIoQ/r3DI/rhg6a1/OiaJPmNSoM6TRRXDEz7N
NO01b/lIK3VNXGAHKbTxijCHz3lw0Oy5pFlB5aGryRpq73j7YYVFArWn6KZb
KnwFRKXJKnejrYDpQNoSr0bjgvKLgAiye6x9wszuTfuLJB+BrDypHLEeD5Pn
kNz1neSH2zdH6EVlmHyk/sPPelQQNNOuB0JbgtxzK3nNq43hAYLXU1JjZ3DZ
CX4WpLo5Q2LkGJ9kWkXDxfuJ+MyEcsCCHqNGLwB1KX9X3vDsbIN5dZn20wvd
l6IX6TWx0POb5MJllH10++MClLMQ3z74OdEds45+FZf9PJMr/403J9HtYUiX
RenKXvycpvnn+FWRZh4zvgIH9+iHBXZgoa1tV4rgLPjIJFbvGo4xibZq0SvP
zhIHozYQPhrmQU1toAZigwCTh1vgZhC1wrhzJ9IfvCk7z+YBzD5gwWrSMdo2
dRFuvGdsonwC51Z9tkh4+OPTcpNUzF6B9f5BYrZMFudT7iUAH3UUAaOXHgsh
tBBxTmZ6ZhdPcjtRM55jmzTQ4cusGLI72/95pNLiMM8A3+DV+s5Wrs9x2XGc
T2PbLaVKHeIiIh0ZzZUrYe21mfCzHmx/B130QTccBLDGe2dYhjGbA7CMurYn
w0ODLKRG0f9ZTeBOdTQaZdoOKC3/j2305atnG5PeDEzfy/Fs9nbBl99Duf8A
eOpCT/06K/M8y6qRhvQTRO9U/EX1Ct+Xin91ime/VyHO0i77sI/aiiVtS/5s
3cgsq/k3ooX8C7HcIjx4dYpwMwy/aCbUhRBHg12xjRMdvoZ0Rp2U8Q18oUWv
48QVpLidx0esWIx/ot8OkhzwtrGXTyjAo7/GN8XBV5OLHV2zBLRRX+tTWa6L
g99vYkIUTeLZaUyByMfjLohvKY8LZa9lncEVPKAOSsn5aVELwzGPKxHT13wv
EkFTVzFUOEi90aiZoZoXqt7N8gG7T+yBxtfITv2KMIhIaIcgf5QG76Z2V9Pk
g52oM36qNGb7VDtjKqT6fjc3Hn/LNikF7LLZqpb8jrM+qOL3XB6VIBib+sKK
EhLpbzGj+dv9jYR8Frdo50S+17kLnntAlHCNNoa0VC4WvwUEuwj7kFADErqi
XlNjubpUu7Empur3KQvBi/RXtYEhTKm8pO12VTxG6vaqwemtZ/Fyoow3FRwP
ogu3Oxliek2BHVPJelnULl/PrKLSZgxnm0li7fHACONcCPFK7lwFe0NeOxX+
+AL5YFUw3J55737gpYoBw2LFjzwgzrUhKP5RVYH7yvH9uxJOmhh8D657AGTO
eSgQ0IrDiroA3Yqn506pQR9Tvrn1ud4I+0Ym6JiDFzmqErEmzO4y/DIvbzos
4PyroSxT7jKN4IiWwMbebEkocroTp/ZZYp+dYaXrt3wdoUIoFJyTr+2nhrFU
Q3ZHuZDkAjMD240U1WzgS7HaJC86C8P9YEhliOVnD65tj+sWK49zo6WVhWFS
32EJRSm94nD8r46iz1UKmbYa6oEbcERnrl6ZtD4483gcJiOep0GQa/Fmj3It
3CH2qXCJW6d8iy3ctH3v6rMvCzmD/6wk/ZS+hUqe32bdv9Fkeze7Pa1ObRaE
O5ajW4rZaaZ8B6k1Eaq8h8GlECZTW/m8H0fo5zG1uTQ3gEQWw0I0MPC8SqAu
IASopc/S1I3xRFNBVXgFNy1kM4+pEsTQbj/4zj9oMSiDCs/vL10/pnrqmoQP
0jXKZnTsFDhoSmdKVDfbew29v8GDCA+u/rECFoMh2YtMdKcHJnJ81dOyuNiA
aG7dlQxomJQhI9igzh0wORXOGSHZn70apeox4v17j3Ql7m2CO/zk7M1URJL1
DqInKblf5k/q4LNfy8FnMKIwgq5QwGY+HRP7Cd4bwzSNVGE7/3RLJ7rzuhdW
ulrvAIDWXzyLNUgNsEePCAK5YeeaexCOBV5XQtpaKIBOadsd2IUC/baWUUSd
UB4PMcdqvHjCNnppkph0JoMjbzSBlfQ8Cjqq6y4cuWuJF1XwsKjL+JF+sOSd
PzhfV5lbGmTKmlNpHlYlNCtJfyg3zgNwdGm9COSgxXuHdwLjDxQwPIcr6cVg
R8wyCJWNvITC7qlSqh7NJcSkuL2TjOZS3SRVu8ruvuWI8H8Jzq99hZbXZiuQ
f+rndqkYxssLJojtgMoEJ33pTzTFaaES9BsDBw7Z1jYoEBeadPOV7mI3FjEx
d2vOEOWmVmvVAXKIIdIMUtUeu516U02NcR8sWD3++0fHUtdwWlbg3HQjjY/D
5BWAFPmEhB87IB7tJWEp17ttwdPsfEUIZ3Kl//aoGCX12urRSBUwq2xVRxiR
2tsJ2bM7UBy287UISgOOmcK2FsrOZ5qhaiPTodPsKQHBSmfxRaSQP5X8CiNP
aIWeHfozgkzmSS1HW4qtInSTQhMYJuuxMKoS30Agw4SHZsOmYH1ae1a3EORE
IQsKWdlxvnLEGQ0rBnTGdJyitH8yzDpixGyDihvM+2U8zQ4wIxwDQwaqhf5L
tnMSdxeEqXL2kCglnNkYCXIMYIx5+IeceL3TOMk6ykQSZwLUqVSs0if/ZH2H
DvjgmxerXD53Nx5kK0H6imO93P1p7tfnOQex2J6DbS3bRDyiZJV90w/SHibe
plpKFndSpYAVaBJVeMz+D3o3mdZflCEEfWp4u5URMKo2sBE5YBcSP2acph7j
rgo4NbJ5p1n6ZvYbRKpT7n+LsB6sPV9jQhCl/dUvU9zQFhAKVbmueghnNU4h
XkO52fefYksSkOJFVY39CTKorcLm0mQj7MfcaSQIciOcZEoMlXmaZKVbtbB4
GSWw9gaiu+Ue6w5+dJ9XZDqva3OjQtQKuH9cswmB4VgeXUreu5lLfwcNEiJf
raAUjxkNwJ1CSYMmyTLHowLNO3e6hY6odWrXaL/3lcgHW4ToWGLOQeZe09xR
9Bhv3NUe/7AiY9EgTGxyxZ+8P7cid//LzsrlHfNLiY3lBeaqdqGoKlVWC4cU
Av+LOHvrAW6q2kRKF/KmQ3+N3rqnPxlt2fDy3d26BgE/qh3g74nFumATcfps
GNw6kZHaztgifzpORtgeTrJoLnOnHcctQ1d42VzvGSdG60OlUSRrqQ9JL9Kn
6Q3EtdwXjnm7SQ7MRhA4EuMhmY4Ndrv8MrgYUlZ6TN5AJSX6dX4Jl5+HXu7f
BZAdYW1lmLLc5Rwi8cce1xv/TRsfsxkveILsaz7Y9sW6XLGR12WPSze9N8MV
4o0oIrrYxuYADSDAtekMaJQNMpsvgxv1Y4xSVeS2DKhiVxpdfxyn3cQXTxo2
LcRHg4w8hHYpxnq8lV8fh2+Wq9bERrvIrUY6cEjcPZUrPUIkArgZkAMRlO+X
KR3Ijt6wHZet0lUySGY7Q2ngukxk1AX5hRcrtarU+RVrIT4Xbtsqj7PP1xU2
m3mMnmLFrgbMLfq3qi2g77On/EhwnMJkCCfrqI2FWUH2C7C5VgLruRDFN34+
OLLeNCc3GweRHjaVD4u4PYVsNOvUkJLiPJp97hDm8eah+Eap3S+ORcpAt0Jr
NwTsbCA37OqK5EzXhpMgSDbsOdzJpYRmW4GLoE4P4BRjG/+Z2mA+5CemC2MW
QjzayvlCglGlSqEDnkeTxOZLygGA0qZjWxuT9V9aM31xBQ+08mRvMFI8kae0
JjGUylqilO34MnT74e5QGsJiHRE5LxS/qMJWWqrje6KJ0lV+dOt/FUJI3eC5
qGFd5KJS/+IG/oxFRLKig0MBBUOlqilnyHx403KNQ6pm9OMoRH61kiG8rQZL
JGq0GSFMDLR5ocae87PgPuzEL0kkQog5gtRvVyq/2QHhJt2+3ajGv0g3HJ53
YRkqQuxNbGLudKcD1Nq0CMNjw/oGycDEyV7ABlBUhHTSx0+h6VN1460OMjgJ
xl1dxCCpgPSejHJlbcCNiysm/7gf0EVlsl+dXBqgnlsjhl+7Vi/XsbiA8gJS
9k7R51JBrkcpYF1H1Jvt9nBoneOcn3mslquUe/qqMEEi/CfjWCMfqh5iH+21
TnCSrlk6lLSk+G7JH9UTy3BEbY4UW7Aj5iF9Y8TKEdjlSiK+ZzyN3o+TavtY
l7N5p5Z38ZBVglfExpsZzHTzAsT7yxBhhdKLHsAO37Brw6grnSz1fYzn2zry
Q0BqszoSDdq15pYXKy4sHwmoFWPHSuPWa0kucr/27yH+hDYZjsVK1KvmOUTp
fe2lzO90JIfLpTupG6P4L8FxpgEqSIV3CMgmwGJ82pZMx5quZ2DIipIOTdx6
HZiQSzQoS8uH5MMngBowjqd09/YxRPtX65dYdRgiVZG07KWSVDJ46CzSWZMW
1l8L5DTvfV9yqXhw/cyv4TueafvuE6CPe5ZKiv58oWehfEm9Q/BzITGHuO/W
veJIXOOoCUyC2ETmqjnL7Y1cnLHeKv7AiugsuI4ljU9ppodDxNIPFegbv0Gs
g6S38gxeOwdriYBfIUMZ6vft0RNVBPxUxUKTPDuLCNmJKf82XRntwIsng+zB
gvVZznqMcAEGNsPAuWByJ/kg0VnCjkIlKglqgrX4oHgwkBBPfx+pnT1A5F5M
zWrtI2KRn2Ux+RuuYBbFHMjcBIUyJO5B6E1Ln561myHD08gUjhbGq2XC67qz
dqfToJu1FW6vs290IUHbZ7XvTquVq54XV2xrUnSmhSsx31A916SkiJu/kYh9
eopR4uLPbQ+UJHa2zeInMM34oFy1fDg/o6pqbmdJNUMUhCYalFU0Pr3PE31d
n9svknnotNahmq5VTAqHpCziIq2U2NOOMFS8dSw1DGMVb0xQkUSnnpS9Yl2G
t13R0ixEEuUqOGApng/XsvtAqcWZxJ2v5Y4ymly4SxxmXUeSt753bkjxXRC+
kFv4UzwSZfY/3SyGsz4/JvGJtsJevypjgh8dqoArrIgYtp2NurA9rKM6F2nZ
oTFWR3t2skk948/A6xcelvaef+OWavt2M5tgH4qMoZFFFr1aK3NZ4VYVwgQw
lFAELWO7FSoD46KNlWvBzS9bH0t22Umcjj3pS/vOQrQaLUKuSKhKCIm7191r
yS9+lgSxHO2M4H89TI+qhYOayW6miyyG/5zT5IW/+EZQzyvvML9Ac0ZxRTOW
rcTYFYFRIwM3OUuvaT5/DMzp3WF+Y1ScdU0bnshUVm/8xiSccoPPZdT1KeyS
uSVjZstBSgX+cHzsUj2CkoDkODwarvk5beuCv8myGR//BLFDwf1e5BLkT0oX
va3aOWxitUafyk6pZIEF6Qje/0QJ1NNua0oelE7+S79b/in6BaeV9sWRmlZ9
+eKZ5NuE3aRTVKRyTD34qo73JRBZ3WsAV+psYXv6s8oCI2pLTtBoJQ4yY7ai
XAUXHPQqkt8/Pa04YNKXC4gSTUxvmwkn1yvcA7kR5xIjgnyiXH1vkn+tRUTe
Hy3wSpgBbnqrwx5Y6QM4vqsJvHOkk1m8as4qFjKRrqOBzLq+2Y5iA3nP8bAg
sCvEZpDFkDB+7L8Ob8AHzfP4OGYbdF7j73KTkqg6t4s8+8PVNBmFt5gDsTdF
HzAtTpOa8KgF7v0UMmMLUOiGXs/1yYxz8ygOTC1oEEpLmh5jTSaLMHmaB0WP
lTxryQanpSUair1gDp/88iSQf5JgRVRfFcgoh5DJYIYc4bq6EDYDpmXXHPgV
c9GkpRtNOhRYnMEue9MgTgdiL/2hWbKM59o9Fi+g69bJOsalQszkU9VstTeL
bPcKPju5F8Kos8wR6tQ/KwTUoWE/MzKDmWXgq9zAWzzoYI19WnsEoNqdNEzH
tOlWwnsLuVKUjipzBvASOX0wiy8Ida5U6M62U961gBb5yS5RxavgXJ4/iSmZ
t50yWPeHhmvQCwXIrVSR2O8/MDxjwbW1j9Dh//yPUAjO+m40j4cF3QBYPeh6
i/6Yzl6IbcYnYvbKd5NUaTigGLNl5igaflEG49fMdx31MCVqHGh65ATNWBtG
holHdwsgCxNFZu/+csIaWZMz+tAFVXD+MOvXMwZrMft2DKiNcedflxTHP0o3
nkknobTbT1CA88+F57Hth/u0JBte9uVF2lKs5Mk++zy/VNRVSKcJSHPN+0tn
WNB03+c6BX7s50odlXEQzmkLBHwHcHOs/qYnXZ5UBO1835RJsOE1923ycRIy
/GWAe8l/7PLgk9zAvH7wp30yKNKgdTdcg50Ms964wAxCO7WOOu5SEozI62Y8
OxoIZLktOyo4JwgOD45Ccd+gEyl5WhVsWbmkd838zsNdIuTBmgrC1q7tsHMz
8uPIehMnmMEMyjJvi+N3WI3pAtuStSESEO3ngJb5oONSJzyqZWvJHdsSesdh
hu42u46f4T+Vp/bKD620+WxLRfOOhhxcHWmY4KbIsGOXBeqcBEmMfcmN1/IB
mkm5rIZe1V+nlv7PiY0QPrsbBY5N9bULTGJnY4wjwENO7eJsV4BVCYm7kZDa
hoobCiS4U3a3x/wKCxxFmaBGp6rI6PvGOm6niMvPnNJS1pmu3KYZc2yL9siy
jxqogYZje2R/D0X44szGn2ypmOQTTeUNfIkYYjiOf8o71/Axu2IqSxUKs586
hwPRkedm9QL8vmBrgoNF5Ac5Nj2qKIAS21nhOkElfmm/HDAquBn0S0qh66eA
IaxgjYe41GS5dQ1FZZc4+lhDuS/h8DQHZDPWNRNYmiS2p4r8Q12Sj+x6ql55
xAB7gt4RX3Ggq9wr2kIqDEfZPr1zAv6jMlcfvHsf8rK2k6ScYsbF49mtzRVP
7FBO5IaCZrAJ/r2n/sI+GjZrGuKZLX4nOS9szT4O+Qa1Rt2UZc4JytZR9UhD
JBoZbFgwJ0P4tjDh+Xpe7wszEP1qBokSmARFuLqZZNM6DZLJ8g6/k8vFLyUB
2SX+W2U6S8i8P5yR10D2MZ5LRNIVpDwvIrue8vfj8diU+yEBmQTGEMnnCwU+
SgOiDKVUPkCbB35nBFktQ9tzFQQ2s4pLc3TIL+jLLl4i5KUpCX7vyyffqbTs
l0rSFHZOP0XImZLHfmK8hnioXItVTAx/sFgWOeOFnrfieLp4Ths61QkPMOaA
mbnfswFG33F5YPi0XeJLgQcVHQAgJ1ObaJpU3VSwAV97ugmKF5uK3SrrzSFk
H4KpDnAxVO6bSn1HLpEmOiPGoJ2wgv+V1GIjgBmeZnK5mEn/1mQ69/E3eP5j
ofeqhWX2TDTi/4dd1GOkPXzMMLx9HYfyQxHKZyvMJzjPt+9Tey0Gyu8WJmaS
jZ1FsvgKPh3vbMHq5tDJQpA45GvEXD1LVTCt0vEgu/zwRIFpoI7VsezGGWrw
fcfhRFwXGMJP7m0piua7KXuHR4UrludwUbvqoo/YNQD7VtD3WGkXhpu7bjRf
VnzrItwj7w/SQeej+sXhgyXhzm/9s25H1mB4HlpmiRE80KAwqllRW3UXnxnZ
ssskXBpTD+H082Ynbf1W3MJegdq9SSeGFpfhr7j54/JWeEVFVWmuUdRIqTgr
IFcpZxeu7XlY08J2x6GOf7ER9KJDcXNwyaW7vsCGnGZhaUbMRbfrXfc6dDB9
yZVDkZF0tD9lkfuoceX8MXIFzVFxnRhJVvOOAF0FwPYLCE1AWtPGWU6w9Lls
fTGLyAtBieooefTuOIhicdWxQ+jFhMmIEMl4cD87kA/TN+trmwVdzidqFLR8
hZQRZKDk1oV0WmJ2anImdJEue9huSUtF+tdXbK8h9aIOVUeV/+o6X1S6cgLG
mBg1YmXh++ZsFdkW3RQNrOuTpIA9w5BmClp6g+IAm4bY29Gz7d8yClSgd+aD
Nafixvp8EdX83Q0jLRkVeKeMmcJpi165sIZXdQt58k+7U7kCq8NE4CXyZSPa
ai9vw6Y1JA3jj7SJbJ2HY8q+fNMfEnlQVpb9RfGSHTAlHntZNQxv+XoBx3V+
Q/qBznj7l+MGuTAmQlo8Q5REL1lKcbQM3poEXc7nZ7sb/GgAv5EmiWJoRlVX
RPD/dL3XbSupHqAq3H9n4GmveSCWl7C5xyiRTHQzXCWIKsgOB41M6lWyTu/p
WwH4lLuFAFtDATBfr6WlEqSio9iUeWwsoGBYI0U/cVi4zW4pNM5bG1AVQ18Q
lIO/76Pt5fMC54IvLcvvz0t2A5G+QHiWUVZIzm2MGHzWaM7FAAkG+OOApmCI
ALnWtMdVrsPtSMB/XMiwKY4BedKUBkAkSAJLr9JwBw3Z7c68NiSa2meQFHwx
EpFfU9Oe9s1a2I7GChg8C4WaAy2qdOHDWqcTKTuegn/Fz5UUH7zcVeHsoeTm
u0jkD4fADT939XAl0FlnW1LulZUsGNQ0HK9OW4J7YkOUPMo3W9VwIFGw/8kr
AG0tYo3OILB2SxZ1xbSe7t5hB/nhGkbtJ8n7A16PTJEkS1/8Pa2XRWBfZRBg
jcG58CBGZOEDMrfPM5cw1Zv6wwndaMykZSC7xigIBhq/DwC4vOqSDOmh2U2o
1n4Wek268X7cAt2iHz2pdD3qjBd0iXxKPc9CvI5iNxqOWo9KBBIvIaQ4ASfa
l9VUSWKfGh1oWkb+4p+4n1ezZSvtMu0+i5+uBSF9n671uTZO/akP5Jhc2/+N
AkFZgWY6KXzU9ovLa27Eofqahvqdx/9Dry8aPsteTdXHLiZY6co1N6elIKVG
HYt1yR+nio5NkFIzxzlhCpx6s8N6aEIjxPqsTSaRClNnRRER/cxqiFaxgDyG
SbeB65hQVRSAVJxbBwO4aJWPUycw91DyjQnTpDBdo4brvEQeUtRAc8huWGVQ
uWzjR9KL0Xf11Sq0Us4HiAUvy/lX0n3jXdLuQftPVF7GaEQyQw9fJWA3gKJ2
SpTpMIBwW/wyQ7GllimoDX7yu5uKZ0f4Rg+2jiLYE+3FXgyo95PPzZvu5XaP
h6N9PlIACYBq3tzQzYApL91gKiZvXfs43L1CwqdjxH1ijx1PQqB4EKZ3itR5
IvCgWpghcHhxKDVWUxy+bo1NTddGPA976lh9L/bWofHWkCDmvVct3fa+d5yA
GIeEi4qMOkeG2MkDHYQVLyBZvWm9YoPVmws+sx1y6Mq4ZiUO/+/o/8HewqBz
7kTln/mfikRBcPV04KQsY3M2Xmy59kezNAOXbm3EHJ3L/ylLQYvq9zlE0YPq
Ifhwzswku4esRqaDN6xKlPKHc0MT8JXTVl9gYOjuSKBfxihgbQLRe3jFTgin
/I1+BBqhEVxxtDLXaZUhEBefnlswjzQ9NTtdQzawhH+KbmVoyFw80dHzlVNy
/xw8RHYzAine/KUgKV6wkpQu00rQnEd3mLPe/eHzSVf4XCl/yIkQ5EWgItqF
q7p2m/i/V+s1PR3PPtAw/EHEsq0lvZrQKvzCsczjMR1SOFyUxkvL7CZSIc1w
LODi6OkrO08HrCy14OSELKkg7YTCXODn8XWtJdHUmRoxKP6MnKyxXj8Io35I
b+a7/nzBCIMFogsBnX3hHBK4EqJGisyWVSitwaV2dIZhXrl+Po8ZhrTUEvn2
m/3Cmi3ZXQGZ5FJjkdzqlJsRsVv/9qW7NGJc2dDEppt/3SKXYyja2GCWfBhk
obMxtRdceM/568Ab8FTL26a6QGKtPGgly4vCw1iFy5tv4+45IsfK+TWjXP/1
FeWkDm3kbLAY8J14lrI5hnzlUnWGvrckJzVMwcR1HvgLit6iRI8z4zFJNxzL
8/23ocP9AAHa+bLj0VeOVCEmbMk2esE3Cs8y01dCvNG3pPRgXlHzSBext2l8
16TetSzKknwwYVwDImmiwIrin3cDBabwZCxLb1D4jRumOZBGl5o/n9m72fgC
dfcKjKBw6fzFE/UY7ZlqaF4Cys3fL0ot9bAeV3WzVJwd7wZjHjv0aNJK2HJg
2CdQF+nmII+/i+4/9hRmny59A0wLjN/81LWQI2hwoG3LTfDdZa/47CZaMxrd
rl6MyQaFUQRl4/55OQaq2i87T8WKHgFU3RKlC38uivLCw1BujGfZV+iFa1nS
imp1UCzJLhfxYkeg1yriMBLr4bigoFyoC572v+v+f78TMZyGSDP55ehXsKWe
LeUUfyQG4VeqU7YN9cOjH3frJBib2jxv6sBxj/u4eL7y8QPqSggIbVj6g5xy
yhvgdY3ZmZuOaqFKf2HAfGr7kU2icFjfiMLVMN9NKYRdFhn79pv2xyOYMXHy
UsgBhrIRXqHwTTMamJ3sp71g0ljf74QBeSJz6Dc3iE9GyN82ZIA/C7z4kSfJ
BYGKEW01tdYKYhIkvtkYyGmkYhM0INH8ypsJOHyLJrjcYjO46fhw/G0AOIKu
P9yq7+C8GDpqfydCkCgtzskQFZyOA7/Q+vhpmdgTC6QStrarrzEFi0Avt6DZ
8gtRmqug2sYsWNBExialF1iRuxJtQ+JpvglNFRK8q9cXGhKHTOLOJKFjdQaM
lujlQuTfxb8pzOHKqo26g0Z0fivTdOmdF8QJgkTnGUq99EYZZrugyjyoqD6u
KVogC3BkE1AY4rU3GSjvg7POOLFA0Mvso0qz86oUs6+Z36xevXqBlAPhk4c+
ubBD+/CzZS8bG20uiKh6peK4nKWIefniJK3ADDZWaqr9M+/m/do444F8bzFv
ilWyMkOixDp3b/AVR2tjlM469bfZcaCMk+MVSHwsYvea1Z6OnNpL4ZNH10X6
FBHonqt+nK8TJkOYLmspsMKJCywZdxZHiMk7PYPGjgPUPovPfYEkMoIyQdRP
VTpXtraBogx5c6BF3hh5nh6euZWg8be2VCKxWoKn5eSnMsiMdD8HUf2uBw9L
yuBEJXQ68q345zd9tLV5sfExXZqC7jb2VJAgqLyD9CCB30EmvZPpgG0kaP4e
KtcaAPr/ZdzpdB8PA5aYIzLJALGkeY0U9V6xO09ShxX7iCyOnfl/lOJA0ck7
UXJrtivMcvpoyMjneTAi2GIsPsjB+qtLeueyfNF97u8VCFl838O0lsLrHqe5
9ShEDkWnD+NAZVxcPB6SMZHIUxn56NKENPKN7ht7gcXrHZ5u/YyCDQC8RE4q
uO80TIhqjJ33966v0KgF4JGZiME0AKz87fGEVKpwxmchJsiGGjwhzPPgoX2g
sAsHtAwiWY6YZVqg2D4vpWKyPKGsZO2BObRWb/lRa2J9MZ9UH6CIrkv/X9Ia
+kAGd3+80nC8qLNk18HOB8UH5q1+4BiA5RA0ctw2hGAwP7G2w1JBziV3+dfr
VDTAbSUyJx8i/Sk/WtEHILHduc/dNkd7gwTlKx/QtBlBuvLgbGk0t0uToNcl
emvgyKUln40+3Nm4xOuV1Ubzd+FdPOknTFY5uuckTBx0CBW0pZnyL2nQJhql
ymPQQIN0mTohEsqh2FTH2hrSNUvx+t+KFMzql59vBTatsVEnQyZreCRk6e8V
PZrIZe8yTQ12tEd9ztGndL/DtuVtToIXnss4XOCnrdwqvKI4bsNezZLjahXh
NqL05KcrePWlaGFTnFpgr1hRrV2w0bb3CxOtiQlW/9BJfIvFgjctnw2GGioF
fJ2hGO2wWLWl3Qh0PeNE1oBHnopVZl9b1FRghMrv6pRGNJbzSDS7jsUxl1oO
sGhaeKklyzA5FDGWfzbRUXPdN0oNWHJHzosS6TmbglRdFWELVm2LwpZdtXKH
4dLkBKFhmWX46MKhySJkMyHzEc8Pvgt5p3sdAoiBbGkgTWrG0KSP+/eDXAoo
q1xIOdatWr7Mejh6kX/SQqa9SWeircBo/8MDx9dk2z8Gf997minvhbK47CrQ
a2aDewZvPyylUDsBr14lr0r3149UjsJMxRLDJ3BB0cA3Mcszr9I4TbONwoD4
e/Bry7SsdnerrsIhLHYKNf2S/kkf8NoIDWVzKHPYujOyfhBySnTkrKc8NSTK
QbKO1cNj5LRbZNe3XlEeb5bJueM+0mXFMPQltrrk4Zilf2QPf7WO2NFmoJ3/
koO8PMm2O4wd2hO6kEE32FjBYC0hkwFWp/2G44H94GyfxuUvWf/IWNGKkM/8
vEXmX2jdNl2Iwcfazd101gcHz04ISzKSncPMAvOqyeWWd1bcXcDKHsPEot9B
/TYOYCB8Vg0Pt9MpkvkaBxxNu40xulfq5wHC4k53NytrNZKkS0LT6uEAD6lB
7CLfdjngD6IegFqNFheRQMZX+CuNURjTnxi7lTHBMVGWNZKUcE+aJ5So+GpG
Sp8EI/s4A2mZeKRY6O6VG/F97aPLoOhyZ4wOrzDk7Ds1ZlyaEc4SxslM/O9J
JRIZYl6VFcZ6tu9M+NA7DhBXS0LzmWGSfG5iuOyNoLQsdX9Uf40mJ8nF+cak
77T2FJAgyFEYgPPnIvyhwErvuL9yjaZP8yttD4uwG1DUz3NMjdoeNr2j2TCJ
BjlhFZ4aGvZLOMQInCp6JQLd+4rhzd8io/FF34TPERJkahAzuZD8sFAyIny6
cprB6uSNdnQx6jgrPk8Vu4fNJdm+8oObQkZDFfFPRnsuosvIs9PJ6v77bYTc
w9BVtX92vx48WDDKZSUU+Fmx80JsqPP26D/729DZgJSnCjirDz+DGN5bjtOr
PepY2jpvH9HySlNiEjaA8x1uNc1GQ6JhSve0fAl9JwW7B+q5bKp7+yT/sdH6
Yj4pQN5ElOeAv+EhoNpKf1UbxX4oC/QU2Cvo2fFJck9Sj4vsWfu3Jh1R0o8x
2HLe7nGuWtjNR7EW6rIdfDwR4QB8PLWI2aKyq9ZnSDb3b6wQG0HkJmPxf/0b
4faYyDSbRVmK+ct1FjsKyUToVNGvjnjA+DdThGvCCKXhG0BPVLZGi19ldyj3
k/CLMbTOIF7/zqvISQSHn2VIks7jAxMWl7ZrP6uwY5X4T01psD4KL/M/Bs1R
O3W8Z1Z1jBsLtIto7hoVDuAQdD0rjhHALi2zxBK1JvLm9bWdWIexHcKCXwXy
N65HddVLs1NDOiL6l6nYdgI1r/w9ihUqryNGK5LE/IeDcOwc85XEHV266R28
g3kzaubzWMGs7KkpkAaYucaBwJiJX7mFwnGSsPWYszHoUsQDvL67K0mPLbmu
N3lg+9IvAFbLMXVl6G5b7m/tW6DZdfo92yjZaEJtWH5vOG8vW8sKyUp3awEu
EiZ4gxRFEXi/ExPwv7zCytFvocydG4tS9ffKltIyzZxqvW6kpgsBoglG6tS+
p27mGO9TyQJZ3ZV8Vz/tNSkqF7xIn7wHFutlD4dfqnac42heaBI1Ll5j0qqU
UQSSlmI7zAL1qgPWNBRmtVKq+AgET++VMBi9FUB7TBDdpGsFOpDilm29dnoq
Rxb+o2I/tg5irTQndYuMI4JHSWus66fNr+b92eidFSwuYPeO0Ar6pWz/k4Uq
CzaUOUtxP83g4HG/cMrQP1ldM48/ZrIOWB5VpSmM1pmA8rVZT4ZiQmv38dLc
ccqo7wkhiQFKEUav6TGtNGSJ0b5/oXCqVAmAs5IwExpET0LkqYnRFqM1b+br
Gl0xYDlMX7uJVufQPCXAjQsVi0Q4CKLL3cHDRMU7/ry7gftDyy+aYc6LM+2b
LS7eGEr7C5GRG8fPnasapON870N9gSimu1TFj8viot63j/6hBKkQUgHGcMGU
yMNrwASUJE/XQSg3D1zoi5yZBwJD7GwyUKgQofLzuoU1m+jlO3AU+E2LxwdN
U0FasjspZOFczy36ub944uwTi8+EVwZOYyy7/wn+rOW7tA9tEBez0B/xm/i9
rqXf5a/rqTY3kvpuTI7w11qiGMlYpU394ZkRwn2PJ+63XcEvHIShwuU5sfm9
gWbVsUQGxJGK+AaGIpyctq9w3QYGy0sLwGP0Trl3cQeIM6OOLM9K3GkVHf4a
MfVW4LXvEw7s0F7WNDznanxufQ06+KM4befmTCQkKPPciulStJQKgXFIbGLJ
pX/ZpuihsbmhlA3bkd497fGqQOcWbcJkT1P7i0CwrOZXBsns7c1uwNZ/bTtL
Ip7jKOWjJvmMWdPhHwhcstIgch1/QGFlgU/tDLIBVXNFdI851/cFnl354gkU
zUrbpKDdClb8fovCZeUOY/4D5msGlSJi5A3hcglqmKZlBs01Qbe9DbyeNJdS
YuxFL/q5QdGOu1ZEYT0h+Ugn7RZ+5Dc3lprEbcI6yeC0H8LnY8B7QH+E3MBS
k63GMTubYzbBVYJXJCduDDlyYsbRIubEATj3EL6rROQL67JN1a5ffusT7tI/
QwPkWWGLX7/gpKmfIzjC+WkDwoZut3VBLi9G/y2LJqY80iOtfXp59jTqRHrf
9PWr0Ora/SnPJz0etd9r4wCqtiyr97LCquKereYJfv6FfjG8kg3b3P2pVilN
mvgj5zyemBPsOo3NOU4ElsjgAFTtc+QRXvIlANvwPvpg2JolTk/VtAypLbA/
Uq+XTVl/Kg2NnVbyMckkraNoVssXMIK4QluNj9c8iFljpFjDt/KHILNnynaT
AAAJMfmER4s9Od8VIHLqXqdXkUmzF8DlA5gJR/E4AUFzUToCLTIeMgm9HRU7
oPTUOwAOIPQuD/pZGd+5JZ3xcmE71d1WRhE/w7yScgO+lrmEPoN07UZyHzvO
Ux/R+qRCd41wVMpigraSbQG4aUzwwaVlHiX9sAoezn7Cb3Gmj/fSBuKWm2v2
CIJ0H5xugtdpQyZRGOx3PCV8hGNpBfHIIY02AzE/3O3vZ99iDq9ZD0pntKu9
dAsLX+sy1ADmDxunikugt4WvnmLDSWU3EUmgVQgg7YLO7Z5C3U+ku6UUlriE
JpZXnaOVsodZ2MxYHYOvnNE04Ek7ogig9TxJedRFcJoftNTEDkFHw6KznIIl
b8eU8pA6zMJAewEbgdHjfslH5CXp0T0dGPRB0RgpwWXb/VscjKjHFnH6Wsi2
1e5jJffOL3vo12tEcCMqF/AyZI9negxJs2seONCwmpSP3CHl+FsbuYFDrx1J
M8z90yp+Draj27vDKlBzOoKbrPg0n8rQ1rBE0Px9fam6WW5QiYZxCg6LFB9e
qjMLvLtVtECGpPtadwgiaoMiQ5NE6cHHvmLm82JYX1mTMMqbDOrD/jt2/2Oj
RBmil33X8FZA3mVzVF4Gzgm6MoZwBaA6ySKpD1YRO2gywAFgNpORIT6Z/W17
Vxk8STW7LsrFJP5J5tV4VnV7UstTMyREEVzmmv0ZsxFW8qZm0H90QXhWdY5H
z+UyII4sSu7MHRWk8Ng2ge0DG8DXxa3ZEFxYVo1ifaTFaLQI0dnaHLWCgIhs
mVTJX6m/itum25JZVkYuZnQFfNUWqyLClUZrEKgz1BIhq4jn+FOxPsXkmXN/
XjQSXhvZsAx4kBifaLKR0BXwSAbI0mMYJVZ1ejPi7k7pE02t/rSbLMhtd9fk
7bgqtrL/32VPtdotv3YyMXRFSVJ0xTcYLsv107i2pmFpHJGxmQnb0YvoUmed
P62NsWjWC67MLne65x23LqC2nWe3uk40Z2pj5nNcyKoISC6TMQQWp5Ft/4Qw
1f8Emt3yeQyPvaoHXkAaQaTDzgC1+yMNPXERFGfhOi1oH4ogrS20escGu+OJ
xWvH0MpLAZt2gIw5yMUBo7G1dZUwj5UllxcwSEqDlm/SgMG3EOXj/mLMBF1H
42rzxg9Q4DHTdcF9PlgkXEeyP1iH/3EJoPxGlgFXMWrQGzJU2GqQekNCH+QI
QgRy9TNzP0ju+/8FocWc2UGuQXHQxw1ykki1SdU9mqN3TffaLFUiYRGYKRsz
fUDy5Ca4XhpXrUWtswyrmBSTfHyd+wE6EjxhSvtveXguEyaAfQMmCsw8fpc+
NbWgO9GQ5u2Mp1HUPVoWAg9LceGpWT2YbR+DbZ14qIjlyWjgrdGJ4zI7hEd7
hJ6seZ9Judq9WpbgYEGbyVDQvElR+u6OtVqYp2gBvFwW00B5uVJG//AFvGqF
UHJ9N8icKFedQwq/DfzDWLgemBR7lqQ8gAC/5rBe51nMn36B7kNNSwZvlHoA
7BKac3OL0CAuKydoXgjD3/qx+7PqfFlYIOxj14YggJYc5ySkxksLD9sCucPf
9ucVG6XieWtXqnzD/JTbBdc+/of0FBk1BQ9Bfg9zNdrSyHoZiPK5BStuAWHO
/sLst61GYZZed1nsKijz18rFRIMAvMrj5MgTtvGWMioOJeZTor/hYM/m+XTm
69bRXKvuRocSjVgIQyDkSd2+jeL+ITJx2tCgh+Cv5wirYIb26QysOSs4SRZ9
UWWKiaoY/aj8tMqBqyMsZDacBvtCYNoa/zvkuL4G4d7qKdNQeXKezizcLU09
jtivRXHVOo29dRVDHGtcujFGJGnowMTMmUPmTron1ZKLwX4hf/THrkOVqiTI
eQSAIX2Zlk085VU3R9AgL1ihsRNf+dXFmtGJ4h32ZTj6OoEw1pqoWivf7tZ1
Z8QCj7SSIDwJ3tCTeQIXVpY7zpGt5fCrT71PaPEsNqA8zCCdtpl2gqYPnmvt
nnKUuRyMi8PigPJus2GmHGlp7NgL9p7oHdLvIazvippr7p5avPP8NDEQrzZI
J/N2OaniZN6+p9gN6BErXxI2fdavlQAJfHxvlY/+mDhIPpPb7HcNd9346I1y
MuW64uYnUx0+KNDMixEwv9uHzIFGhibSTGBMtejLdhbZM4mWjfoz01g8FbMS
3eK8QCJnVGdW+DWGZAClw97rcfucAhlE3O0yf1wyW0CSp+suTuP5VHyMSgD/
DMGY/CsmdPIn8v9FGMTVum+oiud/sJEEZMzXOst0BTgQ+uZ6ODzLp6Rf4J7H
Na+MZU3QbY9Es4AWo+byUFSBBWMSV9f+I5Dla1a30tvAK75FhWsJJoAO8GQj
/iBKNjZFG3pGXBTZUaE4HbZ+cFPw8V4jn7zLw5wF5i8EY4ps6001X755WHK5
+hNO7Oyf0EUQd3kHyMNJBtYFv0QqWwi+jaHi4W/9SEE1HnbZxd7k+krnccTP
k1ezIgk6gBhaIze0ozQpkekZaXLUQ+Bn/nFyILAckrFFchuQ9ra00OqKFPHJ
Kwp0yEtb2P0t1L7ivW0vRBh70uPkWgWatfAeHVwsDT8Wb80SiXGPAp12Rnhl
NY8yZVzBYmXhelVb/EH0pxFzpKEtZiCoR/lciAAwrbsOPaHFR3bQaLfaRSFY
fZmrB2CKgkCqx6Kcax3yTrO121aqUbN3QUgiQeqBTQpTqjg5JR+EhHYa+Zuk
5J6ulFFAlDsDHx1I9DluJwbZ8S54ZKtGHbSb1xoChRXMWcIMe+ARbOaRg8pa
asGC3xqRAQLdtvMrye/DyoAnNZcav4dE3Dz27yLAhAbfDSJ0YogVjmaG9srr
P51vbicKgrts5IaBTAc27sHpwjRaaGzTYvRVBmJAqTu6tiKZJF5AMBfcsDvn
Wl+QoUQOp2pmNza8G0l4kp+bVGTNQuBD2/Sw1YGg+4PsNvHA8BZJGhTzdqFP
G0GpINdZiCxIawxH5+di+uiC0s4a26lGtK3PBUwDXHx5i0rom/6fvcjznPy0
6CkpveZIAlSr9wXbTau1n7R9lEFHoB8/ORdkTfbfGxCm18k9r+o5tJqDl17v
iplZg0JbekGCdnPS3WazKDIpM3wwGrQ3z0oynWvT4SirkuJ7IbbfGCtat6Dz
bwXMQW8Q5d58VNhqzps6yQhnJOo3r212eYgt2yh8Qkr8p5OB7udjug27aWe3
oBljDeiWrlW9OI3s2lO1IkfxBl2grwKoPg262A9DOvy6TsfDCwRSaJ1L8PJc
uXnH77muGR/vjV91DqI3S52xuiXMa5Gj3HCINMPJQ6dO6QdLrCRLiWYguCYd
0kaec762kTwvt+HGLUuG7bpxetEPmtrKjdpGlsYO7Oga/fZHo3pwRnOMAQ+x
31TfiBzyC0x+vjGxJo+Eae50ykCV7eXJ4+W+uaAb6j7ZTo58I9dttD4Hv7M+
UdEiijjv2GqocCoVje3wV4EzJtXZRAJsmDDwnzrVTG4w2RD9DhIQI1DNe+J6
3YhfNEgwuh7CITie59q20OIgH08sBwKNO68UhwUotNoyb+fijAuIYCVA2sl5
alZN3RoSFJea/dIdRpAVYoxU+sJcF7IiuquZqgzfegKIPgq20Nn5e/R82eab
iLIy3gnPDko/0NHTzpRMErrArzh2zVtGzePD/a7ZH9hQac45EqxtTRXkJNc0
qO7PWMR5Owc06qO6LBfVkTG1k4sxxWJ4qiJ/OB3EreH7UCGwip+orZS55n4f
xhr9BHUOwxugnMyu6Tu5xB709Nfy6ta4G227etuxdOQOZmx97Kees1f0i8DC
Nc3fzgjKTbXFOLX/Evw5hsvFbtO/Q/NqWySd8wHmU6gd0377Gj0T5xxIckh0
0yXCIseLL8gmMKXIW822J+EsbHl5FGeNOAzPER0/NLJPPfwXAkps39f1od8a
iriDNWkC0vOozW1svvjpF8HvyNcg/6nD25MgDNyI+mpOSG1VLanMQ6otQfXc
qDp2N2bokhnCC/zs/+zjKVa5MJYCqQCC5g/4fL/M2Jl816QaFCRctvvz9uJT
FhSjB5xo8o9va+Zv4X8fb91/VcpY+eMFt7vCf+XBnHEq5jl4976ZyChlgnV/
cRs39HsQO0MfVPX+hyl/pVhLzUeoITCUiK2cQVjdgGRondFTa4X3MhGRmbXd
UIDTJ4PPvvpyuTEhbvwrDFE8bnQSDFxqzNp1H7K57CurFGuKolgoKFF9Ijqg
NW73p7ij0ONgyJqkmGcOsVwVk7MSJ+ra8meq11RQGdM2s66PCK5kK04/BSi2
pubeAr9vbjH9236MODIlhl6yTDFK+V+7Ij+avgseJ8fxPFsaYN0JQL7VypKp
aZ4TU4QZZshSpxFD3GN5jEmh5gj93ahYsnuTPtvV92eRlXtDkFG3XtaELzrn
K0inV0+C3FVj7Erun//C0WDlrptxmP2wB/8Cdne9Ob9rIHlS7TalL3bfHf3v
opkgecdhV94Ip1GMF+XfXFTIOjeWb6dPInA/6uLHQ7XIl81Q0FxPDTUhsLSK
RMOJmFVaprDGRpS45NAcGr9N/DLWoVgBHFmDTZba1HWr1diw3Gp2D8fUW6cJ
Fz9pvlh1APHebjJWnDoAaR0RWsBP8E/0v81mXwpDgh6yrbQmjkkiU9nI500A
5z2FFxTa2wIGVDt4mfB9TYYNEnxLJxEw+uay5Or1Bs4V6rSNKk2/26gSoFLR
8QO8le09wJt3Njs0ZBbxONWIjE0P28JGimoqiV3QLYm1C7vax1O+HfuuW7ds
a5pNlW2GFI6oV4gBVWycXtk+Ev6ONKIKslOI7n4vJtJ1N6TfToKxfyDM8OKE
iwJolpf9/hb4se92iMg4bIOlY3SIqfGwT4bOkNmYuDIpyLNQI3MqMxLzwcLi
AIpYmyNclfZmPhVKvgKjR/VBL1qURuaLzkzEFbdVlEZu76keyEm69LVKbrw0
i3eh8OGVdIGrxHbCbPF9S/3yBtYw2exu2OZD+7IYTNWuXPYprmZiWpy7Mgck
HsCyBKraTnfXaBLNV9wxd4ItZsO97N4HdAs3pMyoIBwYqVz/Mt7mRGM1M5qi
dE0KBqDQApPeRGv36k46y6TXauRfeYaJQtRhLKuYSV27/J39ck/HwPeyXumT
4PSzmXGHl9DwRmRd9FKi33vpZS+QH4hry6pgDKMV0SJZH2n38Is1FmRxmMVu
T9WxiaOClvhRN/mlVdGqnzjtQl/X5kxbGwNQ7FjBxOwijSDrxrxU/49LhUIx
74dcQ733BoygQmC9Lfs4jvPHGz6MFnwv8ff8MmWrnMcAuGvfJ4VIQAaHWuyp
JHXhgKC3B9aE92dEWGpvqBxBkoBGeQ/kGzgSo+ojhBDR20p/7gT4jtaCI0+s
4omjZ3tYTy76UA/Wm6Smgo9XrBuGwf2twBhen9zpR2Vi3EVTdbCzfsnl0MBp
mCG1iouMrlQCiy4hTfh7WJ46JmKQFvdIprSuRTZK9hn22cWKvZT1bvxXIdzJ
y7z0D+VsVGb8/EkARnU3+V90Mk1NSbIsWecQtujenKn7G4Mt4MXXiAQcFPlj
cuGLrpRYTut2A5JoqOihSC8dMvVIu/vY+qoZHee/gY2ppAgJJYiCBlcMAF9j
vZS1mo3y+akh4LlOnBYVg3Url7c0tLCTGsqR2ArfpMmrfXd06eRX48fIXoBK
H8sN+AVyasJvp8gvHqy9kaxG6q7kscrukevdnk2y6Y58nYltsgOIhEWwRZMq
x2o94Aci4T4/U9htDcdCVc9L9NJ4sIFgzImLpfZFnU1zswJhXrk0or9B2pR9
55HpyKOuqbCCCpq/Ni2Eu5WKUWvyljX+FZRYCbdQiJRmfLwKtXrBoPPmZi0t
rVAFL1+hOCiKWr8YywqerRvgAbY6/BTvdMjN/sWiRGpy6UoeNW5BMcSkTBjC
zOfW3WQyhuzZZdRw6zS81x02rxlm6COOmzoP3CKixm1AwdP0GWm+Vokktrrb
fVRWnssj7EJ0+XZ7DTXRdu/PiO2UfhnketTjeoH3kq35zlpJz5byCNtdBooU
tH3s2HdPKVJcwWOVOTSkRbjBbxZ3wihowegYG/qqz2CK62wp3Z/vG7+Yw3Hk
B5eKhKKfbXrWbiTNkgqCYUc+SVfsfSGXWm0rHFuiFyOivMOiw5+B+pVwlkOe
7jBuuwesJHyTHMwq1/aP4mXL4uUe+nbG+7Ddob6+WwdU2lWND5Mxoxd4mfAt
+8zWNwIO6y+Kvey5FXkuhbULgZqnti/eQbMZL6jedn87ZQe4j1ziI66gjpVM
Fe7630qGSIJOVbSCFA9KQSTobXGlUcmKOXDv733d/8GY/kPhYkD7ujfuD7VO
DzMDqM4O6j/t68bagz7rvIJgvY+OF+pcF2gtFFR1OlGBv3lLzHsTEUO/lSLK
CL1oku6H6EO023jRHnGwo9pgb9BkRXQYtpqtajh4HRtm3VanZqvwP6nf+2hj
ssC4IAkqPp/PLk3U09o6loqgXzJqbZ7+YFltsyC+SLTWOYjxhR+c9+NL60dD
dvaDrH62YQcfi9RJpGlnzcaAzhxN2ihK5QAVIfk/5no9bE/V3Vvkvr1uVQBn
Q+Aq+XYwIxOm4JGnAci5f3pIYGlyThILm753PK5K4eo/WOG9ojvkUYFqZ12I
qrQHz6ax2hC7k96C9rGz8krLaZkMz7tXiumm6tzhxodys1xdBHmKELaavTOO
UurFSkkCmsIxjEA90q7TfVxG8UukHYQL6LdM8XYpun0vKtViQdGR23ZHy899
odOhZeXVNo2aCWb9HUDczFsAzL/c9fWGDTCIK5955ecc/ow7HAKU+CCjDPNs
X1I5nWUY8pnSgTKwgxYYMdqwQ/qQyYRveCv9bpa/tFhtImXQyYD39VQIeGQ6
ikGECKH9wcs8mG7hJ8Sgj59AlvU80n7n7p9vJhCtRjR5QRpTGjbmkgcGHiKh
eVTXrkP68VKDqJwbdsBFucUOXmmHXX7zeIJzeM0CazJd9PpEHHBrvPiUuM6g
e/0PBcPvZammmdxfH+vQYzoVQNSM2dlnvFEVZXuyqSRXmt4QI5G3UVCLy0p5
4bO1e/vHVIKTFkVXDTN1FnwPvQpjIJRtQs3jHET407eAzVeF4lMCVQz/m7Wo
b4EhlDUF4IDw7wyP0W6rChf03hJqbbIkHu6cqNvU+Ij0zjrzpMI6JvaSo9lA
UE+AKf7+tjJEMWDYzNtBthk9+uSX3wSIrQWja04oAyAzInMeKG8YFXRovfre
B1Nni8ijroIqhTzAZKV31LMmOZtYGc3Lpyvgj1CLYhfVndt5wBW9JHKJzXJQ
I/H04AIC8lh4DXsnGycX8WQEsGbTYDvru+l+3Tpi0dhoZK1YXzW9+wRzomNR
Wk+tNcOumBm3StwqM1sUP3HCh8nq4vMGVkceT6q9t6n1y5tYv3S9TskAcNlq
o+O6YmneEGnIhF7JxIE7RzmPp7TqLrfwfmoymZvptSq13NglNMLxyhegHPN6
j3sglL8Xxmo10II0rj5Iq7+VFHh95/8iIDhoqMqiQUWni0vdVJSuFZvV6s8s
zTUeFWINJIJnP4tVWRZiAemj4cqP8hpPlXBlOWBGiKNzkSrSZYMarM9LlF/4
kPZ2CrRsfthQQPN7ghQ2bUrqUmjn9IomlejR4lh9YBkthLdIPdHYh/RGJu3K
YIJztk1KJKIz9rvMZ6fu88zhh8MIGaQTYgFYVX75W4yYx0+G/T8rSnP0TywI
QuwR8KoqynpjEEPE3GksV/umd15rDSq5s9Zo4eTcXFEgUK/Fi/9cBm0bw04r
zR3SY8yoVWdiI/HS9U287RlL0do7Sc4oWro8GCA9VcS8MO37XUqq8ezhmqVj
hoHCcl1NtXoVH4aJy7rFvfLOKruz4BIkA8dYazm57WhuUVjElQz/5aqzOnIS
5nMdYjVKLYs4ONuN7/PyRR2pN9DCLcxjy1PLsVJbwGPZQedVwdTpP9nsbYY2
140Kqb8roYLkdcMe5IH68j857oxy9aVNpp416E1zSJJsox1WURIDOECPkjhT
1rm2Md/lb5zjqHJK6QvXFxzKMBnIZtmFzaOARWYcpnmyMahoR/TVgOyV0dxB
sYbuP2ctCFp5URLOoFlg+QQRCS43LGjzGKjL/0qSW3rfnVvLUHJTJQU996Bg
/WUs6tl2CP/zZvEpJubI39MPK/VBXxyOwfYVejiwjEUSepc5llnNExPrUAYV
ilYCJ8MP4EQn9XJc5E21MQsSqQLr4Fp/X5kpzS9IvJsnhWYB7tY3eHtI3SV+
Wya6A/QOuGd2YMv1sMwDa4Z64FzaUwMm/ZX3Q1zDzXlNrb6Q6HJT4+sPBLGk
DROlfPDQcHNTnV7Hs8O4WcUX0f+hhQqPowLhJUsyuhq1Jk5fW4xM1uYYFhzu
bnnA8PHHzMVJBUr8L1YQPTCshS6g5A06EtAYgBdYo+iR/Pql+NV+nPy+JstV
3mMaA7fgfH1NN7pSaTYVOvvtK5yHI2gFueu7lZHXfKp+R1NiSYawR2HSU3OD
RFG3qr8InjGwmxAWfIkkMuvxLG5VCgx2qJDOtRgBhtRbRsbA7ghpzHti47Kh
jSqNwbhVZxICmgL1ldcdHif6fV3mzWO5O92ZwzaEsxvqmiinscuiPvt47m+8
ROb7UwcZ2Pn6R1eAy9YF89FegiYMoRNBVSt2I1N0z6B47VP+J5odwFAhNKq1
LiaRc207khbCci4OpP16zCk3dX39Z5b7od+qAfT4mk/Q/nq/k42E6HB3jC2y
P/mBOlpyGn8Mh46wRkzANJa7xKFTsWqDgl+XuOa1jFoH+EEa+LLhahgPXN5o
jt2scXkASBf/k+4CaP0r2ScHd2LX9l3ED57OB5HTCKgnsMV55wAW1yT5ULJX
V7QyXhtI+WH7lOgFzOQXaWvhElPMFNjbqTT9cTJVkT1rcezO/pqzdrYuHscG
OTQc02GBFwHqnfjXlYI3uakRIEbZWew0L8ZaWWTQ4Mjf8jDWG8c4GwDAlnlH
v18shrVfsbSqoWxUCdYK9kOPjGX/C/bKvwqDyTS1TypCt0nspJ8EPW1eIS8y
mDXGmImwpkPClkFKC3c78E0AdQNzc7yzjNheCYqbsdiCHBl55neNLNnlNG6y
BzPuF89MvO5cFoslBae7yiarkt3TGL8FF7VuWK8L0KY6OmoaEBMnsf2CwYzO
ivdxy4vI7dWV7UDzDPQfgogpQefUVUZ+qElsRBk66+N+IUy4uEVc9BTGIpSE
3A+NuIb4/dbrsdXUt0mcjda13bu+diDt8G4Wzy/W9epL0sK62mvN11TF20lL
UG6GMdFZ9eYVkzX6hYhiam/B+Dln3IQ8Ofm6J/ph8icwXD6xe1kFmwGqr5xb
rgOXRGYS8e53ZR8QsdKCnW5pddT42+9K9bL+wu/oQBUlKQoefmY+2UoFHhYq
6Ydx8GiwAD4iTLH2huy9u+umaMS60vMjE6kYsXjOcJiiun/I8Lb6cmNyVQTp
Mib/zk7FECkS9vACff3+EUWHmuRpXk8/yNNQVBakcnAsUJMgD4aKmBP23p44
4NoEjYZu2id7ST3za3+TcPlfk/7Lb+ZfG685enlBnKaixS6/Yc9RAGKVR7Ed
DQ6iivLNMAgqTFnjXGG+/KYvvyPCjwEeJTA4MxzijpLOXlMPW/HnxvscBvnd
btRukflH60pzTgXTC8jv4SnMql/z3cN5Vram+BCXKF1HNo1Rq0zsjP/OIvVu
jTOrJW0KQrmcraUE052JPNW88B/UXxyMt6gY8st6oqOI78AcGZSpVfiU0hVN
HzL+b8xfoua9W8/hC3phee5hX7m+JXVwx10mex1PkF81z1GMWvryGKJDVkcc
LHDTmlpVdatG/ELl2/9YvuDg1rRFL11JWeC9PQMN+idVZ5DEJsbJddAQAOl+
dGQ9XjcQXkZ+cOy8UZLZFPPEsefP4Qz7Tupi6EoTlZ3Vt6Z68piQOcnKFz0R
ko10PvyNj4hNwYhpLBWAa/neUuYdMtjscgiGox/Y1Yg3UEnz40RVs45iEgqI
aIVUgP1ew7bVHXK9xnAd1BhnZBkvQjuB2xFs7xR8MtXk4H3QHYWRZSWeFJu0
wFF6vB/EBfSL9DNjUQzoD4gg/GWIVgljBaaM4afuqbt8M/DKhUBaLP/THXHZ
w/9khogBDCvNf2kP1hqmWl1Ru+i0CO2rC4vyC4Phd029xB2mwyyPTq6XEB/Z
x4K5ibdbMt8STMYEJJcfsSieWfwztEr/RxWT7QewbZkAHPsTZ4QWoX2vJwK1
JFHC8HuyIUvxj7X7+K0xzx6ccjesroi30mBDxFTdO6+UJxWliRkqakA/R6/4
Fb24mU0q8kxnZ0NwFd/Uq7BXWF3cBHEUjRoz1FqJOE7QujjF0x/j1CvFV1vD
3Ig+YDf1Frd5zdBmj9EBto+/9GeeOiSiTNfIwmSbHBAAhuulb7L56OyJVnL8
eujGAvOgOTDFMTZcIrCsh+RgvlhNoJ7PwoDUlBVu0BAEcE81M16dgsaLz0tU
LyeDAAlhcMTUiDjBWOvzEYCoFWEdZVThjHgqYLDaQ+47KrE7k+hNtT/68VFW
cWL0CA6K+FJ8+mpXx65uJs3f9WvE1qEVwSeJnBmftwxud4rVtJ8NU+eTQrA3
blEgZe9tdzsTCmx1jGKtftvr8ZjirP6P/0LzvEiL4vjdTKtKQaw+UW3bJkNc
NFY2+AydKARfE/BLS8Gu9AaUdp35W0K7bUwK1gwcPF59cMntgVu03OhshI9J
fR6q+Z/OgP9TIRBAqED7XnQDQiTbIObKqwypcX0wu2FJ+7T3hP16ilYhDmnX
VWQQT0ap2bLj+oWPtcKW29sVWsjQimYZe037rg2j7QPC9xkYEEiq4URvzK8t
64AWdp3CAVkjOU/yfTihXqXH5fmU2MNXDe1zwvkUDhjWNd5lDNDsyI0ZGU+p
mD5z80UYrfRINF/D8LtFDevQe1A7G63KANlBng6bLSiTeIcKdV4FjS6iNYFL
pWkY4x0IqIr+h6GEXRKnMx0GsMpL7ZStCfqjntDr+Dbofwmbv8qAQDmCwyFf
KSXZFc1rki02B9J9QpVDn8rmtPZm3YAL8/GmBZMTjth17kn2DDWtXuuk/+iC
uhcdC4zW3yqE0InKxjWtwfC5k8XH6aWH8lwod+M4mmFUP28ciCxvz8B6wwoH
rvU+/C2i9AIFxGy5XSc15IPGOKFO76jJV/4xlEUELF3eW7Ck2tPB5a9R/m8T
qPboDl5uRevD9KIA2V3Xh+7cyzj7FBIqC8z75eVspsWuMB7TTQ8giw2QHLu2
aDWlUS9Zg7HdpGPRPadfInVMUEzPJgvX1D2lP+J8NP7WX4YeGpLZaAyTTKjf
80BiRtiI+p9OQ/h6sap7k3zmfHxnsw+n9IEcX4AsxJ54hbn17gzS0nxfqxgy
53LNr6X7EjaiC09kUvxuF3VhmMjW0m1OblXjNNqJYPIrB+3/NBo0qR6hxWNA
OZZr8Rtm9sJJYMOymd/4Xqh6vXYGHujblL62Ad3BiCFgwduxghVyz6l5/HAg
6927ZBbiA5gCwm58Y35NYfeD+wazfImXUra07Y6w1x3EslmYFz+O/M6wU1ko
lc4lYnv6oCAI1Ew/ifCiJPR/tpGWdY9F69Wj8klkzV7V1NoMxXgWzrgSsVH+
Xfco5aQwe59WrLWDgdFOAnP3aEtLti1QgkcOZoXstk1r5DekI+7cIaOkHMgZ
tYa5dFtmr5OlLXO4AAkRHm8xTXj6yOUmdPCVrq8CclKu0cIGvextwbHWEVbu
WrS+xrPpwttoUKdwHaIYF4p+TwXgRMYoXjJUt+wF6F3g+CfARAp2IEt+/UMU
Dwqf8cu3FBWADGzO7Q1od6zUlwg7ahKEMEWmPwVBkQEznQ4sqmk+P3pv4mZi
qXqJhzYH6fHIYW7W0YNqyVQGCIbop8I8vWdIlHXsh/oIyfg3iFurHYci03AC
yh9wtjohQKU87462pKpfcD4GXljYTcvVx/f6NEjTQ29RnssE5le0trk+AZD5
6ZqKUX9YmpV5SsnEfZywrwinvotuHXoqBIU87Rp6G4II8Y+SaqG2KVOSo9lx
FIVYg/iGZrB8o1PYmL0AlsdXp251+NYNEw1/dK6zUxpnFom1l2x84vFaAe+3
smPa3/MLZVWPlDtVfdcR6a4qcfO18XWrDAfRX0spAVoZLHO+tg2NYjqJrlOz
k3E0gX0qWSVNt9CooJ2ivxUyJ7f+kBkOwRuBtNzgL8vaFv3pstgvHGN+jE0P
uxouwDZ3cZ4NlOrRZciz9dnIum/kKtGdjSh6H6rQTJQLJDC+5Ge8wVUpFM8f
j7P27nBFM5/rQR4ahG7BYu/4NKll+a7XOHqc5xG8U09XTsloklg/s5jrRzCz
34yvBER5abR3eIZjKr1oDDOmn5dHj+t77DpbR8RhHFUHzm8Ro3D7PFGrZfer
jZS6VsocWiw4bFJY6thm7ksd3ZOJVobhMXmoRRNSV48FAyaT58UX+TiBIw6X
1Zdu+3sHUOpJBSNFxBq1wYncqLOZViohD0XbxNPjUigdpHgqcdtDFObZyS3a
RNq/grNTnNk+66T/p9VT61R0VpKlMYD8I7OJo9sv9kIIC2oSCc2Iu/5OFzrs
Ljzp5P5pzHvaoetFmXA7Z/VdJ4Qc967Bc5PiQ3yMvQZVcIrr2/nxqG7wxV2w
LniYb47ZIY5Bpyqq5iCmfMKa1yGjWhft9GqpC2sbKvt1c0Aws9h5JCKS4V40
EMTZ95YpZongVWYImfr+7QVI6vYYn2o2RgkUMIIpvXF8crYWz4dSY/DDM99m
4YaM5qvmmK+h0kESIB5FSv+Sr0FbFV0nVrC61YZ31BVFSqx/rw7BC3gIPJvo
7baVQezyP3tlYzWrrezDlM4yGXWjm94gLfXZj7RK95NX5X03GPBuUlz95ouJ
LjKvBnSHF4ZcyUFis92H5tptZ7xAFAus0Ae0B+Oskh+8imkahH3sQ9AMR7+7
xF1GF5yPejjClDth1vECY/RsejLOi3pYQOsTwb18JkxOOFrJzdRKpLlOasJx
43M6eofnFqHrFgaKkJIWvyVrrtugWGGCKhFdFfPH2uJF9xWJCRwJFktW/QMP
kfANZxd81xhE7mq5oJ4Q7cp+82eU7T2QSVPBWGfncJVgAYnOG0K3FyVdBuIK
66vi3HAmTqJLiatvqc4NmmphRoSn/9L9+HvI4SbqG7KvG33TAdJdQoaS1Qxu
ZkVy47BXAXk+HqG68/JDn9dxIfCaPf3zLsbhlbEZH1BH2OZRpD9blkjYF4wJ
JEwKXYRRvxRYmWJL9cpXfzLgGX/F1skztPqgqvvOLydZWlCmxBkI6aQAQWv3
0MZ2sdmNgwwjFArnx06gyQY0ffjheKnI0LJpLhdzmxLpN7uTfwVQnF+yqnns
KWe97H6vjeJh4uYmHy9ICXljI2LsG8BzjQGut1j0RNHATPfuQTatHDSf8MHY
Hk4fAAHGYpL2lxLzL58HvdpcRkyTqzxzpsFgjWEn3GsD4IeLK3lJAruMuQvp
cuyN1W3ZnCynE+E9gWsez/AlxH4IhM/tOpuEdeG2NJGhR6fjU/l5+kQIoC9N
0+Zg4T6e0FZiMjbsZlnIgEJJBtpVwu5sKsOXNfX6GJPSaIVfdQzCDepfY6zI
f9ZBY9bJY73BcZMsEKxMBMOvaKA0FxwItPCl4qq4CNFmYqYWkNIxFDKNK5NZ
IA9XcV6+25KgMUOfeVayoqirO2csf4ZxPGygm25TdyycyUyJTvcx9JmtFp/z
K3A1XhxIXB8oJkGuJUjjwZcSrJQHSdx0yYGG3UhhUgqV+cioV3zeF5eBDlGb
Cl2bwFRYjGREXJ6b9scRGTWXV+iyKCkpojTineM3gzzGBpsKFMuudNqdS+xB
/873H9HJoOn/C+TJP+/0W7Lw9v8g/PYGWi66abK/Bpkxrmziuana/FYKdW3x
GM9tf4eU23CKXEh7PWmoA0cDQbJjH4fojEu4AEja8V09ulzur+VJGpzEqy5w
7Krb5L3Aojv8V4xMRgOgxnTdPmiuiEUwdPk3ZljnHeQzL3EQ+X/IzHoALBhm
yuSftF8Fw88ERGE+eyfzI+bIkkTO6BlRq65c/ejFjl5EllM7n3gmGIo1r3Hl
5Y/xkwb58EPLQ+GQdHKV5DlPzuMDSDsGcYpoyC4k6M3B5XhK2VRemQm5nlPf
RZMguRQc90Tj9n/pnrR+F07YPgwwHFJAiIo3RBmCYi2K6XiaUtkHGYsUu0nw
5l29uaue656bTJnS10+wMbIBL92C7rkjsl4bhA+ZTFIz/Yc9yPM/XRHAAMVn
2x8oOz43fmviAdyjEVJkJpIkrUW8OeNcVtJZDUuPkGCqtS4eShjzHzRBZvUy
XMHiYnw+l4EXO1hv3j4LKWs1tUIzvgLnk7lAUp+MkqyAkD6rnsG1nRpLhynI
Ts1iVG1asl8gI/YRFCq9BC4/cl71kZpPLrF2z4ldHugYUc34Zl2s+hzheIy3
h5jr3q7JBYqhJmcAOwGpX3okwRaKQLs2zJeBhDv03xpOo0d/MsZgwh/Q6VeB
GR+XEDFv7zfWoHBXLomJEgA4gZU1VJLjeTrc/mFEGpmHBWcOIk/VTUyxNNIM
EWbarlmLDXDhynyKBlyuDqNVLV0xEZcFhw9vBQkeglwHgj7uDFpJa5C2bJVk
DNdU2WyEZA1ArhIW4iymblsfbN+OvERX/h348vAHAtLghsgj4bL0/4QJOZKh
IES9bvLH2VC0MYl/8i7iCgOa+PNg2U0eNWkFtdry+qp10Hd1EUv0OFWy4u7l
YuTzhrGKSCMU1a6n6uaaVNHKuEwFyPZK3dWFyZdu2rALxqnX5jyXFfEl6mBK
4cYbcXOF1fO1AlDIPVIKFKNfRqcpCtaRp/ZsCLcHx06LnQCJUFx12ZesSyVW
7hMn/I9zngYuPQ/Te40Uk0RlEH3h1je0DWj4ItmVV6tg+nBkAviiYlkVLLzI
xeMYsv2Gm8guYbiiBR9fdeE9zfFtA8xF0tiAy6jCPZORQk8EYytKMEChKoBY
ttwgKXPHiCWiD/3+Vu9JwCynKl38te8Q/tPPoaulX3Og+onOCVIhCKBrmgCs
/lpFvlon/za9A5tYitj2Q7cj0QuRxRkuCGt0Hko/8+IXIZqkBdpyJq9ivKXW
SCbkVhixSMUPWcBQOynYRkYpFNixDX3Ryoft3CxjF/bwbnB6l3JYz6lCFhHE
QlmSj5voDlBDId3Yqj1uyp0LolAqk29jIjCwRCXiU/sSgePvjYDMM9e3dWZM
a2l1vut0Y+/03Xkm02h9KkN/tu9DqueOOW7sIvH3r7Kh8p9koUaF8fMWGQRi
RkqAlicLdmmiZVFzjBORAflslVbbLYK488jSWegw7hg4c8qqozzLPqHjwTsQ
nOWXf4IXyoCuJ/7+4UbGecJXj+VO7YulUalq7fd77jm8cjVZD82fGOEr82D+
w7tchMQxRv98NjYgNQtmp1FAhfS525HZhluoQOASo8j+YeY6z69WWUoqEv5L
bl4XzG9RCypPjGXT7I5/9qQwp1jfBqNVN1t2iAV0oka/mVYeyE7gncuKVu9l
aW6kDtgC7i2CusAD5qfHqrmw5ykmQ0qYkNiqBBzXpWaL4V7RJ0IjtqgC4rGi
swo2MakggMsJm8k2RVRhjc2VqSQRnR+6/AHH/kP3hDzA8ObuMlAWEfWB7GeC
C8nuxUaVE208gzlGqhfN2WGnYhlpWlxA+Xm74NifaIxi5TwwlXHkFSwhVShk
6p6xhxHC6/9NaCVDcNmczREetoQ0TU93dXvM3BqWVV44ykh5NpgAU8WS/FoN
jvyOYbSBq1sTM/cFHNZp7t+jjIlrJEYwPk8JcKiQrhAMQ3ekR2DXCeyOay73
u7qrEV3kGD10l3OjIIhsrGJpw6wI3Fy3PxLrP5rQuuGT7bDFxAAXM0EGeKvq
+5EvGMfRnBcVCfyZv/kqXINtBDDc22x7arliFw9bSsdo5h69UE3miD3C0WSd
SDVDug2yM1gd7uxsxRqMfJO9H1apuQjqMGJTC9qgEwuwumt/SH41TbPw4P+T
7iPJOiVOX6cE7GcN1QQWY+LzAqMTcCmcqz1R/5O6m/mHqn1sHagYoL0iVG6M
H7TbNIFyzwlBUajLOvPCOsUxw5NvavUsQAYzlguQUqR3uJatTggZay0NX5Ly
+JSrvrBecEH6F4v4mUIbIi4Xxbyh74mbejB4sehOiyyLB7U4U4nXrfCPUHiB
bZXZITt1fMdtvGC+C2h3AGBdDZQF78pFsrsqssqJ2zgF5TrVdi6s82EOYB4y
sE1bZDBKUj5W2Oc89CcWZkzPDW+eNfM0fzujUiPOe+BeFe2PLHwssgaFbrTr
yf9UVNksrGczGGLayyMSV7wrjgbPM9nCa9SC2nrSWH8ZIV35KVhWrB1dILCb
NIKKw3ajICZtfxcIrvTaZ/L3HUtyvusb00nxPv9kX5IP94i7u6kzOCA2DqjZ
QImIrS3GRQr7/8BfkN5tzE+0ltYdOT4UWahQo47xevElq3p+PVkX2iggjFC2
/62LXqp/efSWEntKtVoxLwkjr1xwSNjdKXzrhtaBpBV7e7+gZy3rHRoPHSBo
wj4uYFQPX6nf0nWUL6J0sb8Ybecrc5+LHHXLUfRBQqTo5n/YkgZjialoTRg7
f8zOX9vcAeSCB2GDTeKsiHrYauhiN7iUA6NdOCkt4iZO1GHDRF0P7ZU1Z7fy
iYJ9HH/xqS1UHERQZLMu01Jr78Ky+DmlfOSL2OrgvCiS/D0WZHwFcUiRTAj7
5xcoN9sdUe7xpAFyNvMXa3SghoVQ7ip6aYTCsQzHav3CgxCBu4OVsrmv4ekG
6IGsUMHZtrJ7v8Vus1w18N+I1CD/thDwR9PDlZEF0QbcldlBXES2gBzNb3ZZ
VEPQvNWeBAIt9mFqet0YTJ7K9851rTeL/L/u9PXe+x+YQ3G4gP2WLxysVMlO
bampDjvH8P/5Fu1Z9TQZ+h9m7LvUNv9c1MiMJWiJAdqjjZNES0QwmqMg6J2e
rlFtq27DUSdcttwyeVodKvL0+kBiS2h3IqwjSvzWQQDuIMwACZSNzIyqlVDd
+BWXLpINvsN2TKzjQVnnqAGossOaIHr7sXfR3pRt8D94fY/oSBN0sC9YNEG5
w3hghrn4HvFew+J7XrLF/5DoSBVWH9ChhfdMD1LJw2HgS/f23zCNdznyM9mN
BhwVoV72RZipkZr8RF07Iy87Dq8EFm2cio2mrb4f2KtE53f1lkVI+xpsfoeX
tMJ6vyj85/JQK0F2EBwUDVTCdGl462+MKbI+qVPFW3V42VApRYPxGVNhFhZs
zzevRJEXM7UViydUfU17JoIO0AbLjp3X9RDpYnJe9nftl2aSLSmRPxDX5Jll
WSCQmmOkAGYqrbQBhfjclijv2kGyO0Ek19rj10yMtjza7V3mKpIB3CtGlxZM
fDsO5vLRm7A2CkTfWyfhzTAjGzfBdjb6PYWyYdbWauRnEY5y5NMVaC23wZlK
jL2vMrVzvzSZdhISxgScxNhYXCK0zlNOdaq5o9vN7yt4BCkM9+0MzLSXKBGI
4kf1u2e7iHk8W8OCuQwTK4g2Wk0wOk1n71nIEL0CTptvrWi3JNzx3rzYlJMP
h/EgeQ/SDUeZ1PzqcOkuQjXbiiN/Rxf7h63Ya+nlSLcvyar9dqzBW0WA5dSz
lJAaYsBy5jE4XAa+N3z8/86SiMKEBpdT3APyqoUdwOSShpSgfQj+JxR0baB6
2cNhTVD3qWr9ulsOcoBnPGqblVhu10K8VJrzHbhzMI9moOIqe2bl+uf9SxYb
TUVQ2/O5zB6Y5PzXInSOzlu4LMGfMZP6WgJURsxWudaW65wG/Y0gpG+kgq38
HfUtT5TTLMYamS3l9Q8rN7Ka+x9P21McIggyHjz5MlN2NQYYot18vbp1jsjf
7HCMiwRGp5AADtfI7D8btUpUt2ZDBs/wAA7t4Ma+RmCQrpj7dmuX5K4r1tbd
9xVl4Ruxi0dqwUah7CPDmD4iwyDFQ/E5fX5Wwm8yWWWh85RMpqEejxCsq+Ri
FJTdVZT3k6A8PkYd7wUb0xG3wxJ3tYJm2Nt4+tDbBjEseZu11SuWwyuZkIUJ
3wztbeUju5SneIAIbfRuo0RB6BKOQcL2Lfm5gr2cBg1esrQmF/vvnY2vCvTG
TPBuP6ShZAXMTwdxatsoJkEg+IB5SiMn09zV8ZGZYi06JH7/7AZ5JDZtdlIO
LTS7on7yGl8V0kdSqMWCnqQFcU4tYSDUU873OgMbKeizw606gGvbApUO53D0
6wnBbNnTYqAKMA9wtGaTqQiYRjWSZA7E7HzPeYjl27aA57VGSDuUrLUIAw1t
jHukeCoUk0gUOyOHkCUw59JtLv7CNrCGNADdJNtzG0N8IUjmhEwEHTAdslHu
y14r+sgU/kyMdTFIBbm0Z8gP6nveo5eB6Yz9Ib6wApdB4kCQyYQue0wX1HVS
XEkJd8S2DCCqw+mtl15Toex3REhdrcUXYUoh1xlD1p91lS4xQ7FE1i3y43x3
0ISKZ8/1HRy9R8SPEhDjEABqit7yupYXMDqkQ4nlC3D34S/4MGvu8KfE2B8W
1kZe3IJNO/ER4+iZe/iBv3Fm/EJC8tSBZatEF27erj5ijwy5wQKjQTbgFJma
bzDyDOISnwkJOQqvp0rPM34VrSn27c8lyUJZtadngp8a9+dSVnfbz7R/XQer
sl0c7kw/zRsLE1ChkzP2kVlU2sPxdPT/whhkr9VqFm3uVFXWJAbzildI2hFW
6+IrFcfwVPdts/GCp7uGOMxLP6eNErvp6fcmePnDmbFSnCBlQOA3ExmSCXpu
3XUYmhKcLGCLDhx3kWkrhvGmhvFPDAXU2oXJg5xzqKudlamqOLNPbjghxvvO
TuZZBk8xxLjv4PBQfOpqGd6ofwLIA/L8JqGDLqQu9wbzh9uR8IjUFRBgsHcZ
YRvO0X7HyUi9MKQ3fscXQaMP2I+4zujhg4ejQ8EWhtECyezhP9PyYghqS5ZM
HtUhsTnrv4mNNyc0eBqwZcJcYAQix1EleJkUtl2OdVkOoci+Z11oihCdF5oN
TCaPVtnkMwXycU+ewmp+p6GwcJ96mCAs2T5/F19UdgeLQRHK3LE34a6GbdUG
CFJsGmcSd2AfCrZAzsBVAFROhb3qrp37rtAAEAYULdmOASRrQe05N9bm3yF3
p7DJVEluSuHcje+ue1+U31YT8G4t0EGSe6YBVexTs/TVAvucNG/POk4EW4NB
9hYv40XFiTFg47ZOeFOmGWQ3J1kxjlyX18C/eY8I5voPAQrPh50lpJfjC2Ly
Fz1B2fNdJKP/JJI9y1Ty6D/KeHTDe2IRAynvMsRGtsIUf4+axG9etrGRnTKs
MvgpIsHuZggRZQop1AqzHGwipI2BCDJLFT+SDec+f+yTPVrdNLgeervB4m4c
suSHAAn8CSMl5WlI9RbPchvwtqDOKnTiSkKpwjOthWj69AeR5Yaf6cKGIvkt
2GMRtSlGRGqRTGNkjkIwp83tXaeoWSpWYlEHbPqIea5gUG7BeTvJSQg4bFXm
QilsbWllSh0gmXd92NRwiVlJl6uTUmDBexPXM5OnrglUvSEJkPHeQ2OBg8Vj
clnyppgX0F6sqDES8FlgpyqOrVpHBLlZbSrF1h4ZvoLZVuxW97Gv39oAdhJ7
0kTYWYdK93tdRHgguEBuD3vDvcPsUvHP7F03sb17W/iA5lZEiVsX7GELZNPf
1Cu6TkprjIO0wELNRBezs1My5l7T2wJKUCrLMzd4ITyWgN7rF4mJKsFrMe/p
rLF8vYXZlI/PgttITGqvfIIYhV/i9YYc5V9x1tnVeRRlxyMb/hAI/XDwm9RX
O5/0SLsWQqiBDkqzMsAIlKCh6VVfZDdRgizWDpMkdh/+2fPbJZh3X+Djvet/
DSgj3gMEcLAecc1lh02Gl+x6OMLbUBOw7VeljgGZdx271cpjAdlMEsr5pZy9
QcRTe47vDMAMs4kJTuTllkk6vRv4SFhGOeTGbsUR/6w1RkdgEJRietnbjycH
/mB9yjWHm5NXX3MF3RvP5MNCDk1ioRgUFVv04wlSnBy/DWFeMVLtwYTrtxPF
pJa1Cs4xLs4Hm8pUF357cx1DpHU6qYwqTWX8xMdLNaBbkaAWXKqrC1rubiwK
scB4lzoMGVOTulhgcHXCEQKM/WuScqAnZpSZLXgfL96Pq4ZKAoWRC/jfzLXS
O45KSVewH4Aa3NBBXVMvR3IzsgFdUNj8ofCZ22MzfXnSQiDcHaNvjhRlG3uL
ZzvM3EnWsY9r/Sq2uE28lDicy0FsgxrQl6QOhIvrWnqjQug3bsn29JIDKu8W
jT4391k+TJ3weCg+0rFLpCRiI5PCkv3dRcEk+B3SHyDZVZQtFtthjmQ1WvPL
JDksJ1HB2woycWYMoAXosSh9mS7shI6EGx8qGaMNSEREEFg300APzclh0VYP
T48m+Lu6cRx10CkHmetGPLIkGeCPqT3vIeH4hLpqhJebRLGVlflvdLARGKHg
lJtsiwaQrRzrZ6+w7sjNVeflog5KwybrVAluz4BhOIC1Wx/CfgmsSwf4Vdp5
OJljENimsCBNWd5nMmcN2EqH2EiZ4hw7TknQKMzoRXlBqu09BbXZxuU8iY+H
YP+ksyjO/8rdpI89Cifjx7kUeZyJ27syJZKyBrOTDbPLllUvNChVXRs+L/jH
6dNZe3GNSi68C1V6FzWDlnoAEFjC7tA55tovq4KQLu/vqwnQdf9vJrGpj1Iy
U537zL1IZD4TSO6B7z9qXasICb/vqb2LhxvP/dZk5YgzRBsTd4vrtCGQmxoC
TIl91kglq+tOUea91YpbJnkuoTpuojwL+ThtFMM4Zn1NBofWA8vA5Xj201b6
sRk/JXHHsDoygEEqPCZlcwN5Tfe1KxENBf8UK4iYX1ZLSfQGZfvqSqMcdldh
dFabQV9p5nb+U5sgonhQnRGZD5E1/Tr3yMiDDuwfH0imtFS0nQntqpiIitPD
XWlGqGgkyjBFwveu3E8HD7PSQJxp4JiJrT5HM6ajcHm5ZAADsJpGUb/+wo+K
OXXo6fhi7Q4k9OVinUHCywmaopMgpeWzATQQi+wQOzQ2HwPqo4TiQy6t4Abf
e5Tyn+syMAfMiFtZ0VIL5zLmyHTeSLAae9ya4QIi4pN1W4EU+eTWVEWXX8Z5
rWRDQ47iTKLKPeQ6fNBdM63nJea+NTrjxi7CDE5FgGjfEKl+zolAuBaaR57s
ZraTMAlaJPjEYe4gqxQxSVWsye1e+a5U4vZ93DgIiA/GdKfNQsh9ZgOOMaMP
6KWCPSCU5ZMt3D5jKUoN/7BMQD6m514XTGLee5pywuPjJMWX95nq8spB4N8a
jUhMHxhXwj1uvFQNSzoidR0gRoxWJHC2EqFHm9j/YQOO3zAfMdxJxdWPI2+M
8cefWP4Zem1t2t6En70SvdGpaZQWyEzWQbp2WOvThvsruHvR95FkdoJ9dUCa
Fwl3XghXCOCi8hMZHZ2Ape07BLzObqByF3RXSpqhmu5qUqJfXd3ugPZbwP94
dPFMvaaayy1xrLa8q8npzrZhl+H1HJSzBW3I+alkvPCChLzXuUcApEBEnIEU
LpHYs9WRDVYy1liXA8pjqZFRZ+ZfmyLC+Bxk2dw3KaAsQj4m5n9yPYMVvO6/
3EE/1KEYUVVeFko+MylhEsOkU3+d0emLUDx3xUJ1clQr93s0kr/jucBiQaCt
EE3cpIsQyxkaOYcQxYCXOku+EOjWmcORHHg3urMDCWFPmCLtWFnRiE55i211
lwD2SZAe+RazM3YFN8dkTqTpeWYVnt/EXhyqnF3fyK5YYJF4jZOdq89JOsBl
2ISVThxUGxe6atdSekX+NQyLA+gnGiCXfKwNFkBCTQoU+PVCC1Eg3Gne95/p
KgzJO1LbalzdrpCCHevxVWkTFDgN9fUu5MZaqmE9Lr/y+5kv3vS1vnbZDeFC
Xdxt5LgNRWvakVKM7Mk8NS3Lg3NNe7YM0IAb0Q3d+9YvffxKcI0J81YuqKd5
7eYS3rrSikT8/xJ3iUHQSyw6eWXltgmUsNVpYfPLEd55qJmL0kRCZTW9oAoS
E34CRKJnYxbZHsiScRcBjXr6DOeStSQt6//zLQqIcD+6pBVpUoNYe7UohC/V
vyV7Swvg+44KqSMT2Kw4CsCKImEELBPcsi5GTmHW7BHAuVLGFpeyghGo7tFF
uRDcaypA1lh/KKMIujOL6QmI+vOb9XGmyg47jSEixfsHJis0LaO3Yl0N3XLp
2gx1Qhmj0dAAJWIALTSxTcraC6s7CKo66pH2u3efLIFuQhDHT8eHRBta+4RX
8JdQxKTXBjQgnFtKGTIADqlFn8keOllF0Mef/6oTZmF1+rf3uM4G6dG1tVev
3U3bLwxyDaKwalTlo7DYq8WqvKUVE0ElJK5M/S5l/QJzf+28zcO0pYIu+Bh0
JRn/3TzU1YNdImXc6CEreWE6G2tie75qsbeyb4cQHezsEvz0xRVOFh67bg1y
8kgSr4MqajUVqi46LAz4AmYzyD7IuFvBuwtP5RYw8YAmv+7mosLzMSVhNbaO
wb5dCkRFk7RZCV022vtrHoy18KABQcszAaitVqa6SKfVmSHgHLHnMFNnTO1K
U8y1EVrZcPbLMBr0V57Kq7ivh1p6VqBG+9OllUlkBvPjQ17FfuLDN1E9ooTc
YgQ/Gqv0Inmxx55RK+2ZLWKVLIn5E9hJuA7EmDSuEUIAvKGO3Wn6N27LPfme
yH7Q3Bh/oR+m6EjNnHFizWo+01epK0zDRAS4ssgNNJ2mh7YXGRUsBKVqAnOh
51wBoDyFOypjry2qHI4OrjOVXARwPwVQ1rmUTeIlO/WROsj5s8dEpUMdnZsk
Ey/q5aHiQNQBbXc07dOADmBIXIwJLhF2C58d7MCJNx9kKfOTJYEgvrlp2OpV
JI0m3BcRxnK4so3tX5zFuTk/l87O3PeRtq/eNWTRvk57w2TgJbkOh1kTfa2+
1OMVu2wDeZG8tsjtf+3jkN2u/WxVKZ4vdjHYJs3w+hPCbgu+wdEGYMqFa89D
tYUNaEowXJZVPbUBQ6nP6lOSYPZ/246XM7Cmrcgx3GYcw371hsCasCn23XXN
pEEo2/cXiKy712fDQJFDa4dQ+Y+niiX/DzC6DdMymQYlpW4pANyDCZ2U/NJc
zpeIwwVQEjXTrX8a+Pr8pzCng+GtXrD18Fom6kWg3NgLL9yePv7eQDHL/rzf
ITuUZMmKGdQDsBgeuX/7a7q/+3GVKhxdxLP7I4Qca2eaR89qgPk++xrG15g5
kNIUT1sg5u9XFf/GoTdRB1kVLx+D2gB3KRm5ROWRFIinbZcR+NKbLJio53X3
i8LmeLQq4tdDRBsQTVoHueZVFJ0N+WDXGPfhqYh3hT5Zq+DEd38bUXoXULp7
ocA70xUb7bntVv56cvMiXYEiV0O9zokAOhnq2J/Hhz7Ka9YmJN4A/Vc8sVmK
y38IjHXvOQhVw6AWhS+Cmh2lJA1ufaGmxUU5fPTe6TnDlhNxzqvCiFegWuEu
Z98ILT8tdAbaP9ocf464g7B4U4UR7sAUjlj7mdJSKrh7sLbxv0KmANuWxz1o
FIt2G8CukSt0niSElXZF56deQmIBcJ0MBAbyP9yapiXXDXEIn6f+aqnQIID/
DCrO0Y9Oa5tX2933teRcyHhbY1kJYTmg0EhLHDwB5TFdXYTCPrJyDWgQt137
YUDy7ZDCuTqKU38kJckpyz/Su8OFUCCux9w8Kv+zwAS3qN+thIYEV1jLCFDg
55AQOm2K3d9T625jwKs1z1jr+3yjfnsmZfNyOCOR9L2sf9aU9m5hA6nFggHn
N/k1fBFPq6NlUxuKotrgyXYZGQOh0hUf6cVh5b5qb+aeny23U1Qrl/N5Cfj8
4Jt6cx479oqQ88iy86gwKTN5mIYbZovzEj9OSwQbziaW9X4J8mMmqvDH5wKr
25Pb9Q7+NjC/dBfEiMlAH5I7ctwkHN6NRNlcu4OVLoT4pdnJtISR9dwRwaJE
htQZtHbyqDC+6fHGQ8O+eqT0GYJ0PJQMp30eRD9nPRtsI2706BcbP7FSHA07
Qgl6y+jz7ocm1058C0e5kMH/mUn2mpsaMk23JI+o9dtNYdnxrb9wUhLRdqFO
dUsSCnYPsHwwSL2j+024mEJfriK3RDfHd3G9gQk0fRDrkBFgvmMDj3Qfi3fA
+1EtJ8/CMcXvMVnOY5G5egagNyQXVmcAInm8et/CDIG5X6gGshnJ9bpbc9b2
vJ9s4JwCavsnWSo4OG9jJipjD14jfLQz1y+vDd1fO68MqDGz6/qO4V8XkMga
SIyUwLFcCkYSfHpG8Utql0EQNI0E7+giZnvpAnUbUAQ3H3JXZhKGxDQd++kl
LEHUuFn29D6FSDt8yjePK3HV8IPKq+4ayVmlLfATJLOnqGxtCYu+z+1pTrKg
xxsPqTgs+WfyryGYmFE6kPQnLbZf9e8u5+W2rOYNVG3JynJm+6MjiGg0rt/0
xFO2cFdQTHpO43gSGAVgNiqFJgXrX/0XF+0F6DQjlphmEuUweicJfE+zsUqV
BLQOL7rYKMzNy6uFBqTmDjq3xQxbEKp0K38YAv15RQx7Wu5QS1oaGFcsdXvE
sSUSyA+1xx7/AXPgN3CE0fbzrCDnt+HHYTyAVme+vigOwr3CoiNysASJ8RZj
Ez8BxgAur3RR6n/77+P/VPrJVJKUzX4QZv9Z2tGbrC2X/ZzC03zxHzqS5zK0
z2Ts2noh/5Xj+uR5WyNkZeRqDzKsLt6qJ16wOgUnTuxeWWhNO+xIi+gLYRIB
vbPqiktFcROTX/jeIzcC95wuerG9RZBQSQOqQNLmXedPFS0n8P+reERRIjBF
XqEAvc2xp+R37Pr+gkZobJNrzF/rYwUOHnHWRR7+snsk7d0I7hp6dPiXVL5M
9ncZ/oP81w1KERj5k+8Sxf+hs+HgvmnvAQyo03EcEINh3zTENrHox+0P7ucN
ILGHz6janfWDR7wJx6LethfsjWh0ZZls4dSNmZm1yFftbNZqUoU9oFTJStZ9
R2k+iUQLZUWW0N38cMqFq+YXHzBSRmy+ZYd2PYigcR3JXMM7xBnWlh1nVLph
XmTu5qkzlthWOTEcXE2nl7J3rpKFmC9cEBMLWSrAOnyQ9RDFLKKG2IfSedFx
v4pEuMcI1JZ9rRuuQWxHDUJ9642uWD0Qh4D+cnecqzIPRxv2AcqomDoimQAP
zdMwq05ONQPu25doT/hWLzwP8fRRPzCLxXMriMfRvUDq3cR8Tm76DxLidm3h
kQ9s/7qK0Wm5DQe7tAkVMWM+3NG2S11k2sF3+Db8vh/nfeaLcF6BxWqxxb8+
M7hsxaMpuXoeNO8FsBaTMdquRA8sja4xEoqrb+PngX17OL/6gxwjVPwXzNFG
VN6B9SxFoMkWJ4iiQObwr22bu07jttttgBfs1RkFtBUXQEGC/1raGoD2+ywF
Ux52nfYcBp/lbCRteMwpGsW+SApTs4r87fAjNppBoo75KS4+si5aNosMKJy/
7hBBe8DBKZ2LLNm3M5txhbjkKvJfpSvHywmbzP+8q8oInAsfUq8rTxAba/bu
JrNRdvG0oo4osoaxzAwlytR3jVMDA9XwyTAH6b/h+N27LTdkT57OJwHuYz7C
F8BVb+sLbylGn7WCbAJNAkvzABCkoNpgAHnP0m/v8AKZVIZON8xmg4TPe5fU
/Ack/IXzdjAo30Rrpic8Ork4GCI+0u2ZRrTyKFru3UrpFYyEsfPWsb822fYB
TqVPFlSrVqVSeXrURzfK2YWCTCabyYW+ySKzdV+4cNCXmk6euk1xcoK4Gm8k
FbeLOILs6BFU871WJt3MKTFoco0J9waLyzlxLRNy3wjC6HDZRgfctJOQKu3V
enHcX9n/eoltG7ZnBxA2gqRgyJzLfvbX3XblHSYn3W6/B+fFz7BbOHAHcNZx
oFaYr2kpqv/HLTNx59S1PJ3Q1BHEdePWF6RVWtVupA8ZTAQv2D/7ZMcG5saN
X4lSpgyBvYH5r0ZE1R8XDmwfscTrB1EX1oQ8hGrV5+rxGmXK3oPkoBpj0mk4
q66CksYk5hWVvvDsLwuebC0NfHZeDVXmZk9W3PxNTGAdcn6K0vG6+rimtS2v
IfxhBYGNO8QrgtkMptY0A0V2mEHJLHSeRd5j2Yc+XWt2O+Y9zpq0XI8oqyuY
cTjP4IYxTyUo6izjCb5tsohxaI+ssF0xyTahTcUmsCVnsBnkXd8YIr1eUkwV
cvoYT9IAHTXZ+JKvCxTrt7nBzYHUHCwo+YaRtnoQcIPW9v0r8UfNlerMyWYt
oaLndJPjBgUpKB+UC6uIvjRmVd10oDOReyJv5xxwRBJPRu1ujPUaFTrd1FUe
Hc1+YrbJ5+AlcNGcnQcLf3gaFmGh1TOxTVBMCQvaoG3vbUbi7X8gbyhud86a
+apknZ56RsJyBACBneIBBHr7L1N35VN4wvMYmbkkn7Py+aCBAet/MfMyzCR1
C/rd+AqvjSu9OaMzXpGh+JCl8UmgWF4ZKKdspHBDA38u9YHBGg4wf0TYS17G
kh5u/p8bR0cJlkZFqLljVsnHS4vDfdlq7WlWYT5Fcx41oaGx/BvYM5VGjS8v
mfL9MNnrLiwW8AksPtIDQDw7W02jXNDDlR9Mm++UUjgVljKxoE914gOAnH1e
wQ8NGIw060DRtnNvFq0qibELtTlzqa1/U0zlh5rf7xb/FzeEasxJTazBvEC8
EcD4gjkZ0/y1xHtHZGO9oOSj0NGEqShloA3Anj600Jb4aRPFI4ZV8e8REgNU
QHn3IIQuGXzR2wzsTo98nfCYZfn/HHSpm2jLZJ6V1XBcXdqL9qgMYMcBxviG
NU92xfP9xpe7mR7xUtHf9Zgrg1yq7qJrp8dUDEjBCGckJud8Aby+fEKCYFUi
0+kNLkTHub1/fpHqRscP8roiokRXzUTAmC0i9ZDwEGdbOWpM+82yQ8YvwTGu
A6eIyraawnG1JTjIJYAP6apbzfjkPrZfBTanP6uO6Fb+chnLEWAELFof3F3i
huQAr/0Y9dvhrQx+ZtoIm8KfcAiMShPl/l5XMWy79hxtbwSbfhysI4jzuVAu
nNR8SjZJ7dQPEql3lm1/c1ND1nk7jg/paggZ7k+JHvUtBVkbVkkvKmndNXnq
suWOHQ6UY8lDq7UMBi2B4NiOxx5s3qYca0kcCCPuA28m92zH4uZEwD3CGS4d
1xnP2tTzrQzFD+Nbj2MZmlVC1zlhikCldrTK5nGkst7rMNHltF0QsbupdSrb
CjeT+YLOptiKZ0sEqEulZdGV0qea6NXG2G42zUGki0iKSiBY7yNssOmgbpAn
jUM6ytc1wlje/vxwANU+2R05xxY9M4X64uUFlyHgELX5K5aHLC1wyue95ZM5
/GZK+I92EOnLye5CKu7x2ez1ziML7l68DHUNYdjSLl7wLvOcgw8gsgqAgmsb
yQRQ7oZsnBY9AibQVopn/X0O7FvqBpXPJUXv5nEt7JDi8jnvWLM3DAC6k/9a
QU/OkMeDP/6IbOBTWAH+Kjq9Hem5E2MRowEyTYgcOJytuLAoRXPBt/pvaA2H
u3tAk2rF/rXDMOeVLu8Wu8staBnNDq0k2XRs2FWDqfoNpVA0W9udHa2uFuMu
MOOlvHs9pvbGtp32jAZIklTRmwPtWs7MP6pAF+GgMq6kl/EvdrP/gRkrfIGH
8/4W1aEsJ2dJ7m8FmmwdLUy4sYcgSwBezrtI0dSNdDxCTMt0aFX3+WjWkNIO
Rn6ctIzFR4Yeas1uyJQozQT1p/yPsTjCwJK7NeY/+pM4t0LSlOLDhYhAScMb
oq5e8cMQagmxxsgt/Ng5Ruv9iOFV7pUxwkI5IVflLVTs621VS32B/zMpCFAt
uD82b/Sc1YvTBKfWVdnTfC3OzVnO7LRdks7gI0GEN9+Xb0JijMGR+cNHhKgt
wyA3pFbCrIwsPtfj8LV0NjrZlhrFZkyZnWwSkGfBGYAOZhT/xOdGVP8/0zAC
M6xVb+dW/zvgRagpPFZ08daNx5pJJ52w2iHF+laxotwIgt6cHqtNkxCsQdYd
9wCSShYSGAlleqRb/tM8dcUHnVYRlqkiiixM0XUd/1vvWvhvVPmJSZJ9xBCl
807q+ejXehiAffL3Ya8kcZvq58sWjTTr3PCFAxMt6gtepEPVv9GmBeZjaVLv
7why/TEKhj2vGvIdAq2yv6+9ElAGUjZXU+ZW/tHvs0VJNq/YP/Uux0UPUwKa
fugztt98kO1U2KqbXyxyCCnGCvRjGq5YTuNXDgJrfA5lDzIUIfrqjD2d4y0a
eddhFSJavPmdL157i4VKFk0LgDcYWR+38WuxqpMwnZ3BqfeS1Z7uACw/KkMQ
8rjXGHQYl2CJmCCLf1iCjGoeD0GX3OMm/vF6FD01qPvAA2VD8xIaoNVbeK5p
PBwnhces5KN+XJQ5I3bb9agT6n0JlWgKz+MSbLXXYbfg//vWN76WidjxMhSX
FTsNa0jCUmP2ADnsyOaZJ7q/aeoZEo0nGStCxodpT8LDAZ0/cK8c0W/fWyvi
h8BIvLGNj/q/+lIbvHScKPYO7Cw4SuoR3v7UZQ0UKyD5u1waNgMmx1VUoApr
xtK/ir8ENn/5u1vU5GGqiWNwBYst6hze6R4FajAeLTy+UCG6Qg0qt6ZYwvcG
8IjUSuJScat7IYapVY9Igophd3spqVdozx5XkMx+z3dKFPst1yK3q3JbHWP3
MFyrjpxn62P/7o9IEDoasJuv8pQM4fX24GYC3WHWiYfw5wBMZoenq9I7+BSQ
GFuDn8gFsaQ53amACFHbcBoChQF7BnHGRm02dirdaxkTaIyTRpddaKMHfQYM
mAutWlBtQ6gNICEKwrVA5fyZon88u7CsFAHW6mT3bHpuwxD+aHOwVr9ZsTC/
RXC2oaFemwfKTzLh3IedVLVcdsBiAUlpX7V4uRpNsWJ/uRPNyWYBr4lKrXP3
BzPD4fp0F4cldX0ex0jgjGa7aOLdJTx6MuEoc4kxsifXc1zXoZYGfNSY5HEu
gjOjYNHHWzU/lZkrXdPqwdZuR3JOdmUfpWfuPbnJVrQzTMUi2Fpg9rlwB/5M
u9LzAqUrnNWkPhZbo+iLMgMMc0aKE6FFsM/NZRc4DBtlUPyFaZJZzA38XUiH
Ekthw/Ujm4l0b/EAdQQLUiTy6fMYQ27Wndr9zLYvXWlBnaa6HDzh4b4qk4vk
wXBhuBYFuw/xdIeeqNN9DqVML1cIETnbUx397tts3ku4XwYq0vaDsb8HYHdS
zkeSatRWl/rtpytTztpMF2sDBEBZfEtzqZbzjuMB2GoxQorNBJ4j8RUCtlGx
E8rNcT3qqiOV5uLOr1ZY5qPOGmn5lvlnC9rVFEJrGaDtY+4FQLb7b9z6ji6b
DOUCx7tWgxHCRqPgp1aYtU917DGQEdd/kpOeEuzV/oaSc7ReVm2wSzoKa9tA
R3Qf+eE6j6o6CXtBF1gw4IOhdqjzQlypBiRrC0UrZ3F1Uf4dB9OvQdYADXtO
0OStnIe7otdoWsOj7MQOOudWC338KXyorTWlOftlV2ASbT6dlUMkj2NBQRS5
9kZWLOzXPdO1m0iu9JWEyk52pyl/oVuWea7HSrxNJan0KG97f1B10lqE2OBn
z98FMTDzpZOdz87otL2ig8Mfzu12cnYZ6U23oQguOjwy5F60bTa8wrRSuQE5
jXFOJJRndlcmr5/2l9VHKke5hRLYlz5K+lAi+OcyjU1PJgH5nCyUX15uS7CV
UBEj/Cy5Iinpg7Hjo5I5YRc9iXMho8+XmTPtELlQlSpJuGB5HkL1FCIGMAam
rAK2U6UEarkaij5mxHp1hghO1HtVZyMcNYtPzwGAQSLUR9R9N7yX//+V4GiT
oxXwfdbjOYunz1peUYJWJw4tgoSnAS58Q3O1APPXhEYGUzqXQiAQXG4bGinA
gTCug6FfFkKYht5fyR/lRD73//1+6xH1ZKK/Sa3mgALKDpYCIDjthT8ZLl7L
2hj+Cvoq3ZL+isiJdHyqTSIXROBftcf26FIJbBzBRYN05rBbtSHJx+2PvFic
Eng3a7Fim1QtVmamkBzb3sOeTJsIpLsmAISvZvAYbjzWHfDeLE2Htn5uXn4D
We9OmRxnVj4PgJiYnIsEJ3rcYUFUZdPJPowmzo0Z/g7v2J/rA2tfJyytCxbN
Ml7BWPZkcCp+4AMH08QfOpqB4OmgsdFpl+DX+AODcGKj/flV2PwHZlsb20UX
Mjn4wNR0wgKFGDSIyWomDZEwP6w9bHBICPlmcGR84UhnowX0VUM012k3c57p
AL6B39V0EGQw3e8yrXXf/skbPf+S7Uj9xJgqfQ3IkJgMN/hifgfm/XOZCy9K
W/0KzE4nbJSHfz+CO/Pu7J1TJV8WPjPilk2/qgnxFu8Uv4EQe4Nwq4oEn2f5
J8HzIO58QFIVH4KHfgpZ6B03SqUgoYHDPJ/EjXO29ZAKUuNeV0VbMG0I7c4k
ja0ttB8KtIZX6sc7cilvTuddWUy8pKune6m2t0rCzhHF2cbizLnIdOoDXafi
7bY2IKOmBEhkAvc5doHByVx0IoizPUhN/kLGDVOo6LTapw2x+8LJTZmhcEun
SjI7NoIwScCFh3Ys4FH9tR/U3HrABxANsFhJDQ8mLbP9t9WJ3OolZ9bKZWsv
gW3ggILrDOElTADbtk13YbtNmdGSMhnetI1GkhZBpo4kg6B9UfTcYcLgWLwp
JLlpJFukrPO03Rbw0gi2CiPRgWfdrOlcbVne0DhGbZ533jFyYC+a6GVf7WnU
qUJcqKp3ER5dua2/75ISim0pocsq5zMuA28pGFSrDzKktQoDFbS2gsU2CqzT
KYZfnC99BAGxXyH8i8t5wx7schbr6WSOifgaRjHV9WrZaaA1RQtXgV+1WFzM
5yM6BggAmGUcfqgazkymLP1PaMBDfGABON3hD+w0p3eaYSLG7cTOFS3zwKy8
ipqsmL29eCeFQmRUbFcXw8QsRTJCFjZ+4NhucY0kCH3h2j30ViDFoEVe6ZU5
R+cbQbTRYYvVwnPCUgOGOnAkd4RQHqjnLbGBxnb0PTSteg7RUYwjuWkNlGG6
LPpe1wrXh0hTw0AKPLxsb7aC9x1XUCmxtSBglitllVXsUpI9KB7FGqk1QIHC
NfNpQV65p00diOJBAe9vpFjHawCnfsdRtuqKClhwCJ4SmPHyTiykeIL4O5rb
6XOn3agRckzPTapLhw79/fbcb0/4nl4BrgReoIAKE//enaKejvnA4sO/0D+d
wJrX/HGUU3jR7LvDOgSNymk3gnuZr4Z75+9y/34YAYbqpn2VwQ8yMrMExU/I
gTpl+ZzSoWHDjJHUEwJ7JcMbQ6XDgrwkY/zEgZU2IY4Z0Uw5RoE80A8EmyRc
MDI+Pvtm2qNiNxjrLwx+WZEqHdlL02Qv4eVIJ5AMfOr3mM/q+aX16ifALlU8
cd55G2ksSqe1YWqXDMTOJ9CTKGUvYnPhUs0Js/+vlcNrbBoBwocMF1WG4NMA
AqMhM/NxMSTfj8DwFQgWmkoAz8gevu82v3cr8tgCqR54MNQcGU9DJL+B61Pq
ZHSlQWIgUXEZ2hvcg5SotFsBwBHQbqGx6irmd8D8jdxxWO3bvnMhtIJtBYaZ
kenbVqQYzcCIqiPP99c0jduHV2Qo4sN9FVQufrBENIbtD4nufkYBsw7ejbd6
yDUE6uT1BizQgbh+YRRJiFS/u3I6k5adjmcN2Ol3rgaTjh4lpSiXErII0O/M
B9bhvzMo6aKGJ/8l7Q9d/ET+4WlwNCEsM/24oVVEcAHqZDiZiUzwvBVe9Y0G
9ZI2WiJZr2AubeG5hzCpOxeGMZ/X0AwuzcqBv8QhV8a9tdhzOQ/8s4zjUTt6
oxXTcy8Zz7u5JneOM5AOegmuvJuV9lnG1666xhzhzxh3RAyFWuFfIHWsgUpb
DJiMdU5uWLEXNUSrpsyIXvQjbeNVBkg1YHlHRrbTnmEnbmPaAmOIWXc7X3ax
3jxyUJVCF+0zgq3VQxdWjHexlFH+/MCoSZ4oC0f7bhZrI6U8zB8BCOSKg3K6
FoJjfwe0K2pLYeZ9Toyd5eQBRSTKmxGnnszAUv+/g+eoTJ3buXkmL5yD3uMP
Xy0MnDCAamfK0HDmS6wC5QTjWKxz+sg8XaqoPwT+yjGZh4chnFBj7+ERCBxd
nMWrB+vU1wH8ZxLFFEV+8a0eWzwSjBIymwEeiVcD7qtsglHSzsx/knLQogdF
SUsFrQUz8qjsJm/x/27aqaDzwHA5IuXU4QWVuhG/wXFdR5+csvFjKSBDvGJV
HeOBR1dNSr+VEvVLYeTq+YAy75/x+D2erxdPoCldjRMSpnW31qaS1anhObRl
g4z6EDbmlPZcm7YSE27vV0RqItThkD1PzWomVrzntjZQdytltYOoBaJTN3uh
OWbTXvEK4jqhgb9qTiLzmd50XMxTFqhRunzOFDDYTmRt2Faz2r40bsHlZc1F
MVJPrf1Lm7u6N8rZTR5y+Cqx3b8U+BsW0/q8ttIyElRISJd9LfYLCpFGBr1j
KR1pMmikde8RZsVH/zugMvv22HQXs4jvFwj/sQvPhVmWke74yNVcCER2iGd7
dT4/z08BCcpUlTChhPvzPKUra3uEr23V6+3XESOIxvq2KCfdKa4epfWfFTAx
nNFIiLsb3tfTOW3fjYumj1Al8hb3rIgIahI/GHk+zKYmhofyYObmU+Q6F040
D1glenYGhuD8hPyAxZbinFDwxupaq01KPR7uQu6WX41solwt5JFloSYWrlEw
BSWaJwdC59tP3M0EhVEozyYYRzm27WLwpwZO6KTqatmam0cPE4+JMhQC9isP
K1K1MbjMnbZPABfAblF39dlk033HUhtXNzAcDO8qwlGa9D52mKHvKz9+i1X8
KPycFqsODNX4aasdC/Z9ed7gzrsz4qduqTyrYAdmVrXmVAnaJ7B2+0flxE98
MXMHTw9xgYSuRl2hR+em/tCgRbmz9Ve5ryLN6xvIMyz4ARVRPDAvRTfxaLES
fjpGbLl2djBLFm4kWAc0N1wLMOVYK8cJWznhuWcR+AfLvhtg/XQTzRclTQn7
Z2YT1FaJnhEge/MspLNTdJS9nfX5EpnugyIRqi8E7N6SIO47rlLprY709JbH
FHO6tXDQkWvCP7h0xZ/aL+ygdHTApge1Fk2ewfhfb2/IQ4dmB1R7b/wPUj80
4VCuLgUxKJjx+SJKDEPvkPh7pl/WOOYoMBkTuAb3Pqm02dJc1Fajl+Mnn9HP
Jo68K1F3LYQCqc5sfQUipbz/d7L5wknKYVmFZLHO4Gr7QH1qfLgxx24UEQkd
NrNlYfI6YElq9BIHD704PMxQ4rCgzKa0RblF+IxmZCOzKXDHfCoOOh120Kts
kwrNU+Pgt6f1hwFNkjovTr5sgqpGZyWvuofnGhk+e45mubh1UmzZRl2k4jKp
l5hk3TnBoZ6ZW5V/iGh1dp8+h5+oWdLnoMZqD7YcROks15208nVKdymlA7K2
J2Dx9u0cyNO+lCm5ctai7rLZY7GLRIZK6JWpHhMzLihgDoGVTaoYB0VoRiv9
I1lyv2cmWp7F4fSVRWPWEepKjndbx3rb1u8/cKqyIBdEhjL1ds5dDSHQ8HyR
L15nOOKck8Z5VkYw+fcfU+UQt8YDLTku/SsIHGHI/oXd6tN1H81QxjI3FNiN
iyeYSZuGWCSt9cs7M/gEghYm+99SVRldh2Bx1b5xpvv1Q8zlcUWq+t7LQlj4
BeKdSShwghKF/LY8igvxFjnp0WZUxXSTxNKfcig31d8R9BVZ2gKRvGe0NsVl
0Mb5OmDwDxluTOE9ynQS9w+S+Xq4mFD0d7fjyJWESgVkU1p61O+qV8Xwg1Nd
Lwj3X1OFQzdaglOKagTUyzD5Wt1wcO7skLYXvAANK5VV4Jwe9LBcz+Sk4kz8
ztU3yuMTbnu0aF3Js35FujzTKlinM0secViiOIQ3AGxeyGTD9Rix7w0+/ugA
IMyzYKE8MrZLcKcW49ykx/AwDKIRdKg6eIEvPt2m9etE2qxRUokaDQxkwITE
5+QaUS+T3uewu+5D1FzqLr0SeieBaD5Zhxy13yTMfyH/JCV4IahW83Z6pAMv
Jq/lkZsYs4T7OMDp3iMYiO7Vf326klsDWA9ReYPFFH6PLd5aIIFy93ptQeF5
05dK4my+QyfBxgACAJCMzQpUudJI7cq/p40fUW5IeUHwUSzvawonGIH3g8DV
iRYwMGx/N/yRqEAfp9PWVtQieJqJQzk/jufJlvhBUceMk3RKbc0Fa4CyKz1n
TymkeQFxWqQnIFvGM6Q9J9RGD0Y7zTVsdTMYEzPbRVuPcSeBbDFg6xZFd6nO
QnmsTUZs7HcyTbtfKJe1kRrdQISM3Z3hyxz44/jfvdgyZ0AFQuc+/b8rgXXK
zMnky9rQkNInK9pwxsRnHnaePBzzJbWtxddCMPNWJUX4OdAzy8oQf9tfUba8
L2Fgm4zoNBjJ0E8fLNh19Yud/MR86DKo07tHcOLYZn4yNdJLHkGE2qxzclyJ
svQ2AvszW9M7I5f7Brbmlhzeq43coHLtNzoc8Q4FxrbXIgv5Kf9uX+sZt91B
IEUxvQ6H4XODv8b0OXlrXbYaatCD82HLiO1jshxtNXFmQC3teEI3BCfaWr5F
5n2FGUWxvmsuSAYxNJYv2ywZC0yRigVOf6LZ5TWQGjL0b6QVHUjGjFOlgvhx
nTJPDTZOk9GAaiZYCqEn7OG/DHcQk0aGnuUeGaa9MzGlnFKTBcxNMrrrylvB
SWaa3VDQAP/Cw5nGoruKFt0Fy9wcdgRxBDWM7oQUAMT2RN7Kx+FDXRNkP9wT
ey1CT00l5J5dGpBK+UJUJWN1XxmoHCHDAchHa3vLAPdlOZscGhZBFVvbLq/G
rzo0zM9MJI9k+X3zUU7GVe1jANIYmMhNAEP3aBpjG1wa+Yi8oBf5gSMjz/tE
LbKjj7b00Fc5oT+wiY3dNO8xHfN8mxtYcAA0mzKkKWmVEOq2WtqegOEsZyYD
sT8QwaomtL7hE9VZfcippVtXE8jN/qBRmbggec0pKD8B+8i7EjLwvx0jdubI
bWLRglHgiRVTfLuzDwrI9ZXjOfIRLtXxbwR+6Pb9xVfsVbe0A/iVOKtwXxWZ
1CiHzJ3lkc5MLh+6BtgVQ0b2FGqUAEU9FJgwoJ01E/WK7qlkIj+zHsW1kOe2
y0dHv6zj7HAGQUkZ5FJTuETHtXOBdzVkCWrjrXDDkMVOia9uRurzDoCpGo+K
II7Ci9m13ThwZtWJaLFgEp/mOeqCB0ww2vo3iu966pCj0xcVPcRPH8o0364+
zUwTzrYyxZcIzQHildy3LY6VmxQ44fUf/0CurQj4RV9z4DOmYwW5qoca8UTY
US6KH4YaEtW9AGv8bXvuYtEu7xhFXbzz0P/ONIc+GmyJ4rn+VUmPzGCXvwbS
+dcRBxS9I7x0TjqTH35YfisYslBV/kvBYLx/CQFWBGhdiHTGBp4FxOzucXfO
+9Ad61AocPcwf1s9sBu7EzbfYqsdMwyi5ucGErGYUfBkReVJQE28mOP8JJfm
5fcItt0wxP2uto7MdIaYpI41m/mbHgLk4ownoUwboIH4B9gyzUVIophkdHZF
RShlUloGttuJjjBJiz1TQOwC/aLIen8yyzb+e2K/VBnQfFj4LBsh7BbtLz0C
jX7Jhr9CQthJoqCgTNhg02Aj9kZYNoIr+uCZbx9hPDfxvTPkFZsbrYdAfoSJ
Bhmhh7JYUtWZjTxR4X9OJ4knZJz8xBc28FlPPXDeddGPhT9xv0ERaqrPFBtk
r52kxre8tmLIUudf2S1fPQaNALX3cp0vJOL+mXwjejGAYxHSypKrwk8NjYbG
1iJKVNF+quxKe7QxgMVcMslaiZJUywjySclTDE2A9Q67yiWQFTud8lIo7ohw
tvlT3tS0hfRAvQb+uodY54X/ZRVgdJ/RG+MU/26zo+a89sDBToLcGNzdjVCT
s1mWuDuPu/J0U1VHD5SGlNCKIc+ufsEfU1OMGPdtqsNoTdPUhCu3vOuEA/H9
ohzt2cSbfD2XAnAGpFcm72qcUCvtJRLRDjbbHkO2OAYPf1Yz5GgdNQ+L2uBL
OPfEQ4YmL2cCvYgZ6aBlNtW3pJwKKi4h6Q0vykkiVNAAQDg0I8oG4oSGJSA6
i0MXFaHMdSfyn90DVqFc0+FK2VwLB3sg5MGtQPfOzfEKg+ktEyVP7OiDQFJU
abI46CTjdWBSgxxoDukSzh/UQSYtF4tcBJ5pUws1xNA6q1lJrMWmxF0peHZ7
vpZqLwso9QkiLuknUYvImxgMIKtwmQjvDGIwo8GimP2lkXxoRkWhxFNyJoP9
J9Ia1qNjvgQsIdwsyjFgKpAjuroEQfcwF9hIxuY0wsWxKdk8GAkp+9HwSCIj
eixvlwO2H1LyUpwEaamVL3sobJY30xqYuI4cEOzBPbr8PLlYAcTJTWkNfMid
w1ul456KKg/P4nagaHKwTtL6IfiyzHVRABrNNIb6XgPIV45/Z6fwpzSDC/P0
mC76ESDwnSR9UzacuTfscFEacwHrStRrz6tc03V9kZrWLx7CKOuv3p1EwDRV
MaQEWMHIQPy9X3VYpkT9wno2jpZ7SsfTA19VDWNK2AvVdCZcV6Swgu0TBfgk
WTvHW3LbNWngbdT8PNLXL2pgZS4rD91D6obYQKjAzeOVrhEEI6FB9eHpSNky
GpXvfhHbT16HZmF9Q1M8yiFiAaszO9FzfXkuO/k48yp0pu7c82cWHuM+rKZl
U2G1Sg0nJ7uzVCQqcdpFadFHI2iH7m7nvTptL7jlE1fbpPUXDkJQfgZWYIrz
F/mbGTTiz1V73ahDj19NEUOOyuN1WyZ+GKuhxHNTtkwHmyO0fMd2Jyq6B3q6
YFjBVlvkjuJHav359Jox8BSwso0UX1EPjSbpiWEDiRVh6Zg2aI4yzE1F30g8
E/aI5QYCWzKY4hJ8IZK8jRq/HIepKMNUOuvYT0iYfRfv4xeL30NiWVRVo4kw
ZWluJcWj4Dro5Y9V/nUA8DMw4E6RR3eVNp0e/kqeCtQU2GMqEaaTTFhmrI7+
sMex95pwbsEye6Qia40B/kZRBGVJs1KQChSB1EcwJLTEGKIEjXBiY1pp7sIO
w2Z1aLPdb1Dp74SLxLYjKbjXhCrUe+//mJmKIKlh3Gr+wvOx04RKZjUc7QPW
dIuGnuc6nyi73jJZXUaJvQ6EN+ZtPIWK2+z8OsF/JfyMvwZLLUrVcYPRxjSB
WK9WF+c6d66s++NHBhUW2VR+W7dQnHns/7LJgr5wQIF65reKO/EGTWN0xri3
WS/Tt6tIhR5jbmwYY4WBNfQm+OvcwboOIM+uSJGPQd6kLjpHq4SAz4m+dk+O
ScxtprG7/DqNyR+5bdua8PRGYaTBGfJoJ4mbVj2DK2rJsvOR18S8f3ROj8H8
6k2TYIWhDN3UDbqyG4vbg1oKw0q2+BWFf02u3yEAZMTxCWTNAwCK0fXv9VZn
6EAmYeMRlK0uGXxa8q2u6w1L9emaSy9E2ltY48L1NYw95sNJWf2X47lP1EpV
ChdteYNgMcBRcldCzBxDXzQy8iMMtgzJT862KBX8SUZNemm8lS8viJumiMBC
g4evYUeFiFRR7iPZNUMwRPCQbCVpizfOpTdQxcAJdhu+RNhczVkBDPZpWCej
gIyxRf2E2Nk44KMvrcdPT7Dw8xNJx0ljtC/EDsmHIDFmN0ja7224zPA77xqP
OhzmVtJy9iuZXbeTrWD7p8Itq6RGa7dTGrl33DKbgq1X/Fkwr2hHi4wCdMcK
mj1lj9BW7Q57tqg/7YRZ61DOLbQZcD9h64bFbTv2WGn+wMrw/8HgzmkIZV2o
4ZfoIn1+U55ZYJoNdyB9y/MyApBOC50gChK4TIp4mN8OrajcT2bghogJrCjL
ky4/hXqhQIFIi/HqgGzEu3KhltZvhsJSLrBeuBsSdlnTiojm39+xo2fKkG+i
l86t+gdA026Kef9ttZKGJ4Bd7QbmrCakujcR+UbFQpXgOn1t8nce/qLC0Jml
7z220WW1s+AQwd6rOiWD5hvU30t2213WxXrTmR+ZO51iE/qXzp5C9OmMp8CB
0ZmrV1ZTJMOIf60+Pelbv3pW0/mg1AZFgB8gJV2oxKMOLaP0QegzIb3CyO12
q8iZz7AZ4qHg1pv4m1cIuI3UiJSevYy66YQuP7N+wgPa0z80qGM6SP/nbdg9
wKzH1ZlRp/dQhbOSzdTVVKLAm/mDYwo/Hi0V05wveL2FX97HuvG6hljpIOuV
dd2q7MHrpsKhZKSeX6E1HIDvO68visGGKxpMHz6++6FAjsKMjozQkkZyXPbD
3nGMaxbnX6IFMOa79IMfdHJQZidxcAV+NTM9ZHn+d404l69hDKt7fnvMIhDI
sUt1ffKtl5xGOis2CobGP+wpM5PlrEbKULpk8gvsbDzy/2T/GSHmHfg3O00q
5EIN06QRY0I2RF2KPBSC6E6eLndlYpSOBhemXkGuH3nGuVCFOekQHbRcfQ2V
BWUjbvFYq+rpCD6kIEbCJsc4fakRqBX26174qcd8eMKVPzJv9hi2aaTit1t3
pMIc43nMPTtdusY8YlsLFdNTj0WroSmwd+TPxc5TRGNZST94SofLVVSOdtwA
bL5humP6BIyNhkyDaH5db3ImEmZrra2h8fHujG5FFXKG3QwsazEguF4NfH49
Y4s/fBCsYe0yx/Fe2OQBt+GDIOowbjbRGlhyceNYqpnYsLTkW46WmKagOPv1
yWOpF5/QC9Fdyx5vcbfVVnr8C//bKt3JRSjF0ojywMrT8FjTbWvQ0/+0LkFr
BoBhDkJKQPN4B4KTHHCzluNI1krzv2IE+y7Tx1uHnXOyWAJlQmEx/LNCs2jy
Cio6XQpPZioZPSfdC3W+61VEUCXJqjYHdriRInvEOyd0WksTB0O6LJgJRXh0
2X8665BQkgbZm66v0IPskBsQK2ZTo8/mp8OG+49JsTTbaXXOaE5LSYpVehcu
TpBJxiKRvf5OdPg5rwXBPWYRouaDekdjLscTZfsvcZe/jv/niOvULpG3s9ja
KxeEJLV+WuhLnPCC2jKnIFl7VQhuPEGX6Uu16lyMvMfp7+1vHIkM/HrCCGIJ
ZhhfXLcuiWgwHglKj12+LfaJIeuuygDDk+uFBZeokdTRH4NluZzLWV9EyvvJ
PO/LPqr3zdhavdoFp7TgmKIQ/QvSXAOZQ8UFDAzyq5k6VyCn2yDVzQ1e/b/o
/6HAzwPapc3Pte1wcmnynkfK7OlyVOLqj6fl6NwQWsmzEFbr7NhtaCFhpzsN
8qJ83vX2DEdB0fZ4yEhgCXugPevvCCGI9yHnHl6ZQU5fP+XWLRPLYn+BQOqh
Lrm+BwbdbornWIGh343jfmdyTbs5T8O1/wri3TPIZ+PeE7n22fCsp5FCxnvb
OAbrfadFJRCIHYO4sWiZGlqVFaG5vNmuFu0UWCDbQtUeDdQ1gNCQs+mUj53e
0Z8K3Cr6SW8Qtjlg3PJSTxSqWUCPU1S1lIFTaxJj8zUJpZ7roKA6SJBvU5aN
+12bUO3kswACSPLVPBN1a0pNqkOUWOvIygmFrCUqa+Aatz+s/HtbfgqbIwuJ
nYdrmqtEJKIX3lmh5YFoMPApkzTHqw6ekRQNfRdlC5KqS0wDV5RcPZrCrKhS
olLmOMr2SMKAbvdLLFZ/dLbfaCYYFgP48tlcPPoGCugEeT3hb2mxrCW36xYA
IzcvwFTC+Qgjf7vCu7+cDRq9hZIXoTpfusY83RujrBMW7bciduoyg/ucldIz
j769LT7xTYdidhhUAhp0tk4Z2ILGSxCRciv/YBH+XVHSNY11i8Lgt378s7Hz
x74Kqxm//qkW7EAGg9HWqYpCynlV604e4wVAfC+PrZyxuYmdPhFI6fju25QB
qIYd3wPoR2sk5FUsasjtEZeGazFx71OFOL7VB8bhTZ0Q3ABytuvKGtbjCY0S
A6lZa2+T6Npu2IT8CPCF4jT2mmmk91ZasaIkovS52RzD/BnVHdYCt0azVQpJ
m7ZEHDuAq3j/cxh7MIM/MOMrYQKBHbYSRNsUzenxJCmlAodixcfs6quNL+03
5e4J557mi3H/0xKEWS5pq1vQFmj1wOnQq23NfWJNK+S2nB9FHyu5IN3z76IV
NX0I1l2owpnSYLgvGFvQBfhF2E7kYZ1jmXNB035X2aYs7/IZuNDWy31LPEgN
LIQgMkVo5nICKM+6xHMBCvJ/690BHFdBYFkOU8pPAxB9Al2jYLXppLCD8n5A
CR8dEUAdjbcUveQTmGxid+hjm7NCIrUJnSLgaZ/VrI20I46pg0L90AHQChRZ
MxQGYBQNxxZs2zTvVwrjkLCLH0WU3eHBdDQVM/+04KzxXrw0nXa2shGAAzE2
oIW/bor9aczuojSRz6nFAnSqIvNm7/wOtGoCxIWnCrNc7DXBq0vFgSVn1YaI
FUJND++ON8ZJ+kMC3zQY2R+t/LtC3Zh/FFEUZX74tkHBUSEyQYwiZ62AujPI
TwprVwSe8GYmyipVkFhsh3Hu68l9oBosHrHt75apr27v8wp9AXSssvIkMFK5
Wt50jsOfMffSKB+Rj+saWBMY/yyFvBVWZbp38g2Ozx7rrzw6k8uZzMeYsbgv
uUhMM42y6j7hMuV3x5I15tZjNtaeil2DhCV82U60DlYZuumf3dJaWPd/0mkD
e3GzJ5yJaPJ70uVzfJOxdHX10fsgxCJ+R2oCYbKch/B5iyWTQPH7zxixBtGl
BRI4uIOzMUioRCt2vds1HhLk/TTD+SjTkZjy+SpjCGQPcWO+CfXZ8KVNr2hX
WGQ8hZj9DYOBlv9dyEGWhKnnla/y3Ci1dg/TUZ07YxYFrO2f5lMMw0WmOfa8
gNWwyV9qRpVrsVQu2mt3wYT1Rf+7ZINt7fRXWrPvCmYl7AWVQSpukEcS7wyH
V9dsjuS4iBiNNo/rnsEuMaNchbTq6oBkEjiDatNYW327r3FWhwYZOFJ1z1u9
93jjSp4ZsQbhSaVtWTCksZb1II930UYpIqH6Ybma0RwO2Q2d30OmWOxPjv8q
tiGYyguHcTh1ZzRZijtRP+KFLaLP3nC6DC/LSj0AZd92igMbPH+ApIuqB182
LxdfX/sp9GEwAx+d9E9SBnZfFd81+1jMV/1ckifLkQsONpekk6e1m3404ohi
mnimzEWJ/wA5uWNFc8+zEsVVNi+iFk1RAbfXk0ub/G0v0UZ3Ge4f/6q88Wvp
VG8fMKWACUzIW2xz782G/GK50zmpgdtDcCHPUPgqhNaxW/vZEj4LKs2PONBO
H6TvcnCsXQ+VuJyYfvEQV4WZgD5WnQARI9+VYl0IQcN2Ve0RrzFRzx58Tbzw
Mo5YvOeJAjHeeDp5mCdM1zJRHa2ieEj5GWzlfWgQU5Baxq1xTff3cPY+iqFP
o2+BYVZarrIRpKWAK64dxgtOb/t7zJ3P+oQRoXOqfTE6l6BwBwg8OhCawuY5
arhKgGIu6Omb9TvZFbjH6cKxK/VM+icuPX/Vl8oqtmJciRjxqRp25Qpz/Bn+
x4VRo+IAXebXaMoKzSGE1RJt0mCnIl9aUM9brpeSMEJORWTBT/H50FdU+xq1
+HQrVD8elzpjifnCLOltDTUNMnEj25BL4lEE9/gKlx/glJXeLiaoUdBeAx9F
NXMBlWv/naSNAhvJnzrEiSWmacCaNC/qbubNdV7aYiYxROoudWd3DxqrJLP3
LOKa3Tcn5Rs3YNPZ9z8pm+oCFVixN34ap7ZGCtXtZTmTbGSM6if9eMkQDJLK
9dn1ntaty/3jgtEtqBQRpYB2wE4+tg7ipwYdgsaDmQvlnrOyfze1odYOeKs5
s8/+wb5oqnhuYK9vMrRk7HmWY4YNrHTT36/gAY9jBND3LoJvmS5FuIa+3PxJ
HNMuW5wo3ECr+Xhh8PTeAZkWOxM0G8S7nmoj8V0H2s4SkUZ6maOedJCGOjm0
rgWJTs8dQVYqyXHYZLnLzT3169VvomfLrjWKlQSgqyZN2RtQ9YL33GY2f5Le
Ugrl3039XQDyXl66u10+fvMCJAH8PH1So3nKRyiExvO0DxTtI/Qr7tKqyHqG
7BfHDM/ZLaknrhjwFmc2nsAuwb9AAwQf1rmWAWqejjqjpDvyOkT3APVrzXzZ
Q3xa3tkIZzM/zpubv/e5m22PRf3iIQicdieNrLyZK2gqXwshWUXpkAZSXOuo
SNfB+5XevNLPZTL0Xv7Ur8vhkd6Tr3xL37CHasP8wTptRLB/NkeI7fA/egxM
D52DP5kahG1OVJXnS24QN21PrR7hNrNeG41KCsi8bE+iF7zfAw3vX1yDeiDJ
jfjH6sNNmUY6pTOZiWU+5OMTQRNnCDj42wUtPJ+M2i3On6HtUNdXWNFt2aU9
nQsr8FmcApYUuM6IZBNieqjAmJa6PrA42IJKV/JHCZuiNyxdQ3lJsjvh5qsP
4T7yG22fw63H+2jDBJrZ6SSaBGZHy+OTHKAkn7NxjkdHGDG+voghkLk1T06N
7A/FOo09eL3+IIlBMmwGJ/3xlbn1z+MXCk08uEuPyo+HNBwAlR7u7gVkXrRj
NS5AiIaLTptCpQY9pxqXcfr0YPuvapEvyoNt4+HdI8n/JHgSmuA97nc5pIYo
K55CxXEzJ2Y3G0AggwV0lWI+1ylwSubrqwReZ1sXy3wDNjvaSgrtDsE7dHaW
rmng9DRJyBr5D9ewFfDvTkL61X6i/JSha8rBP2LSMrc0fLT6tLgJ0J57NEq2
EV+QUKhtpGhP6bd38ZvXr/Yp2+GNcKI1ZCrrT3kkWqnIXo3qVs3ZKxZ9FMNj
xvRwF9dy5QT6qWSXNRIkcS9cQ0N1QpYnsJoYCcrELy3phq3BaXk3KuR4ZaOR
Y5pZSO98ckVHTef/GIAxNellC7gYB3krdWI5LGb0XdAq8zBBP6oNuMVUtn2E
L4yIIIhlbMVaXL8wzA1VV3i2mD+XscqMPXIwTqYRP2ZgTHXLeu1tH6Enlchk
vhbOxpetwwsOUXl7HCqC/KKaMgi+gAvOh1f489PghwJ0J97flAQNAtQCGtVv
flnY41bgy2hOUS5KbhnUhkLbJBAVPzMFbPodohYCV9vULhChHfMCXZkTgkmm
ozqD6/6RgdKRkQKQsFErzIvnw+boVr04YqzKO0DSN+/Yd68owOI9ViDdOGuZ
0nxPplTlNX1XHR0Pv78I+Ar0OXN2npRdkUhc8fLh07CxFe7Y/LGTwsp0xAqb
3lmDfM9DUyCRDeTqi+14OXWy8V5SwxPmAKir99Uk2X+Cl10ZvT9/S1BPdNo9
CpWiM7UdMw/I5Lx7oOxBPTrz5wRKgPNXO2el7lsQ14E027/vcMwYJJCHImde
teshCtTgUkvgiF8yo4h3FCNTRLju55ansIha+ihsXZVxKTS8xLP/jIisd89b
Thj7cMAAzcfQX0pQqcv/lSCNZLbIT0oZB7Vchn0qNaXcEfBp9sLg1l7grBw2
atENJYO03gSdD2m73dSwJVFkt6IKdOt5Hs2+9BjfSzJvW1pVD/hYm88AYVbh
uhd53xNhXb3fbfT3l+kX0ga5BripQ8b24E1/TMuxA/8NoIHc09DE+phK1Yve
vVPxI0fYbtJLj3G8EIMH7kshcNBLrRG67je3X8kfFPoFNpKzFuz24eUKYw8C
QL3QQf3a1GdGZLlED7BjHKeiul7BhiC8XWeOcVj2nUU6Q2fdK+GjppkJhzl1
5BXt46BM11BoLYZRtbIgzg7AdTG9R9hWV+D3odMvhGJI2KmcH9LDXvYmgEE6
SFsV7AZmuq65lGBvt1qret+tJueOCMqLhaOD8OeMZViUysfTwiKFYH2OYJeh
OAT0EvbI9zCJMGf1CmpohTWg3xVqaR8wefm6rUj5BOuhwU5HGj7AJAZf0vNl
53ASxgyuuD3WDO48r9BMPIvKzNtPT5QtczaWOnpA1DRIbnDWW6IwMMc/a4sd
wlEBtfJghJa7MfbypbXkxjtND9GxO17at3+iw2brqPs0IvaufDpwedP7kk/o
wu35hVgZFg2vOJoWiZm2GuJc2JqMU4iXACQLs55nQwcTresP99wNZj4bglRa
0xZmRgHGXHHHSvupyasGtOl7qMmnkXGU4oRh5yvYCNaazTMyqwzy8HR7JIke
twRTYMUOVYQudzy8ctkT/9NlEwMnYIvkgRsWDnHpr2oRnKHfX7EZJa6p0apZ
OTmAxzQi7PdzzNtteyRKloun9RvzIGuz2KAX40XlM2flB/Vkihl1voUbGwWc
1AYEWQX6F5LBihWqiaCQa2Na0nke0DLmtbvInjLIUKhB6QfpB7UczXQ0n9/l
QU/ygHchGhnBJF8O5ywzhYDUWOpjdYKjg02rFVK/jv4DYVb8lPaITUWyguAy
MVwohw4P4/SG6Us/D6f4uQu7Oo2sHhUw2R3Q7S2SBqpstLK3PrFjuVP65KzN
LfbOkjnzCp4rEX3+n/tS8csN0HZGecM3O6ZhP2wxZtD1H6YunxhsM9c3qtgO
X6MpzL4lOjWfMsxP4TNSYW6ufwc9LsFw9AFstqD/BXVRYTlLmHxMQPQMGVtn
ESO5mimBkB0Qq5PsjMaOOsNkxI+GE57YJOFp5HGTNUdg+sQ4sSMa0JCdqJ8o
d7ZS+gbOps6E2cMB2j60e64FFT3Kob6Gwq+0Rrsr6lWu03Kf8tqSMRsZBuUM
E5WJZF5wBczBsp88vKQdBWUsRADhPolJ0+ulkgUyqC8RKNSle5QUZIpofBDD
Rb+Bxu/7XlQkH21V56r1i4thxTiEh1Q3fk1B4HvOEfHVX8PiOrL8szYc7mF0
7X1I+yyHhr+lB0LdA/E0V+rA/xTfmdU5NiaUL7RC90Y4ilAdgm6ZIFmX2yMC
VaFxpICDWchsWPr6cNiwehWVJTOgJlgAhHB5tO14g/TPDCvSISvUoksN8/qc
BFw8rfhnR3G4zm2jg5VWe8SDbWXQFPziTMsNlm7YGDY/Hm1r+mNVNl8kL3QH
oWGhhe7HzMn6p0MCDmZwVgqU2tE152+budQheCHQAG/S2CsoiXD0nCHuQ4Xj
o7lvfwXGuvmWbqdll0Kd+dqTNoLC/ZDM9aNFXmBS46WB6b3aiidYKtdyrtMC
6bFFzCaYqEA8l3IYPBJFk+dZAQ1ySzOpxPDR3c9eanRK6ag3OrppahQ7FTBT
DXC4OumJ5So6IFwZJcaTyo5LMR3+hua3jkR/Rwp0rcuDZOXc7bGNxtCTyk3s
uaydf8ZSmDuu4Q7L+KFjbxVkx2pdwamdG+HHzv9b6q4mpM/BRllWteJAzaGj
YtBl46L/sMpa4gsOCfltilnUX45S5oPJCxDA1NIcXbXfIGhxHnJTyQCBmYa4
+bS8om+F8OP97BludNifZUsAFew6NfaTyixuFKbH79ELCBV8vuNfwjldTVsu
oJLO17yfzTP4DTVSaswwQdC4wi8hWtTmEXvSVzLJ/mOWBVVe2NPEPPnA14a7
AZxzsMhIjbDkuXseu1E2R8zM595y077e+1eKpIya8S1pvziNfBP+BdL14uoj
kVFQC5fqOFqUvvAmQoLzV4u2CywWk/phiZP1KalwkOjGUNPKrN+i97KXye/s
lhUB4AdYUgKBdhMjbkojRgyHr/Hv3ZkZa5KtCEXgxV7JSsLahjBRYmhng/Ur
8GBihu+vKZISaqXVFtXQkO8p4dFdlbcrjp9GCGw3vtTk9lsZG4P89oU48upJ
ijBpG8kFgSR2mHTJT3LKDFvIxYjST4Gf2mml49SC8ENPAoELS1WjoLZ3QXGw
tEmz3blAGLBOvqp7Gxz+0dKta5ikXEDT3SgOqIM7syr6QXXXsv7jhMhmQz8Z
sXONU+O4YVA4crpg28eTJXA0P1NrS5V8Ml6t6ne9sI3h6LWdGft1UzrNAUow
PBhla4lYVGU+ZHlAdsdUnFEl90Fg5vfVncgNgLIh5/rAfcXb9SKrW8Lus0dJ
eL16zCV4yfWv+7WNnGWBt658KQ8NPAJ25jlW1iTauE6p3cmmB+BLNQU9vdH5
EFq2qni1E4QY3lq2GqVHAHroryjRQD9UNJDKldtP09NMry4VlrsW0JHDPX4K
BV9bgFN+iZyayufYQxI+1ii8kd6RkBUo63lQBf4YCWKQ+16R4QndmzvV6XQI
DfTmD2RdiZ6A6r1tiSSk0E8BsYIE7NzxbUPnZ5ljICRB2DqN9HBDCAWeQPLk
HTKQH7ITgI+7Uk4Z2c5pv6QHDSK0nJGsKG0gG4b8UgtmGeUUV20MlK9130Ie
ICiMOvdVAnEBJRwIF9/aVyBx/9Y0Yb2DiECfrwTQdtQd6fc8tkpAicoLhu6+
GlTSONZTKBWV4pzUW+pQezFS1fpWoYOhLr0e1sliyycf/TKmSRGa27LvBiPv
9QACMU6nCh4ew/7Iiv6FcU9Z/GOoFG7VXPZBotqlhI7c6bzfT5HiDTpojkYL
g9sSUUbCwD3IfrdhaCBl8g6ZO9SYvjzLSSAPVfohn+gIkdFtOlq/o4IB+spU
NCuhAzbpcct2cDr9Mwh2vJI6qzPwNsKDYD+Yxb5dbap8bdpwu7HxIr7ZEykf
5MLgnn0kUOMzd7dnjpw8rDtKcQBtjQE8Vjw5kEb8R0tyPSCeGzA7UZUby/Bw
FoEmpXT8V1vzXmzKuRWPh0mtVs79z+WMjkezV1i01niugi4zFgc5U0MjgVC7
9/4impQaa3C9C3WI3lNj3lHqQQlPlMriA8B5ASa6/d+GG1eLsN4SJhlUUfvL
C1PB/GlQlxj+ZcAyncwpj9SL4Yd98G7fWqYDY1bS5FetVtQHm8yGd+zTecsQ
0qW5DFF4+knCiLD03AG0vNEbn8n8LuCNU/uExfPNgOWsISn9/g6nZVmNnLE/
pqb6OFQp3Q/sPM9uX8l9GFI8TAakFPYpZn5pZH0CKuPNkv+OZxdN0/gALQzf
5WwsDh+awBxPFnWYQWiDupoA+lJqqL9G4PJEQsTeZyK2feB3R8nFMRWMp9V+
hdQdw0kJKOi5eI7lziE7JFSQtHk2UtW+o98NCvnRHsKxls4bTGJ/a47c8tbJ
sbuNmA5lyuJ8OqmadRzJcDNyXGbu5cPnaZWdyVw5krER+NfdTKei7+Vgbyl5
dvGuCgMrX5DafrZ/VPt8wvITSLM+KSBEr0XDkcaC6orv5fJJcG762isahhEE
so0sd1SbHVVwCxgeLSljsDvSDf8YXFRU5xXqVvt9UaYl50vEEIJwcSFn7TD8
JMyXCiwGr5Fy+gkyE3FOYEwRJHyGonoiTZsb4K8mLTG5HxeJZR7gtsOthrSB
r/qPJUZdVRGLiUWBSS5cBqiznEcdLu7jPboTbOXR4w5J68uweWJdDrniTZte
rzC4fyND4rEUqjusZFmkCGNZHdh6u3OSIZv5RvKnpcwIuQQEkP/OpcrCwv7P
jMc8KPYm5yLDJC8U3IsA7ONGYJCJAcVZO9GmjEMw4cpcmNijlQGETgk9gE/G
8kUX5YIjfy+NlNbEidtO+YrLkGYuI8PSUSuZ0M/9+jylnJZnSqOF1MhIuwFf
KQlP4brsXqDk50icvKVgZb5QsOR0H81P5OHaaXG0JmSp3D//tFJMrARaYDj5
UrB7lO+4OAVVr2Jjt+/iPLzo4P4xu7WLFRdfsCmcz8kc+bv6dGYc6wdcvBzm
oy5UjrNAS9U+yPx5teoMAZpNVzTnDWCFpMehiGhqWp5IKmDiL7+Pkl5/K767
zejif+Ql5XiEIayQn3j4uIA2mn2hpMKdfZO3f01RedZo12NQGckulgRhp5OL
mVHPWuMB+3Sp/c0KQSfpUenOVYT3vUThLbuRluAeNVphh8uZnuS0AK/P6vDB
17kvPDHyozoSNbJwzR0P7ym7vM61Eu/ag8oA6RVHCpbsFNe8ou1GsNWyuv/s
F+pNeRuoqNsGdJU/jyWPueVWU+JRSQ+rTztUGN6ocVEG6+EsKDBU49KeZLcT
KSkWz0GSrByYvunQ8W8VrXCymXvYIlxpIs7GIH08VTnC0sNX3QrlvxMLJfc3
luTesIi0hixd65PPTejhdqN+56DlUN+q/qlGQF29qAoBSNlOcLJtHsPatF+S
aX42/2WOhfN5QE1RN5tmP/YxqpSDKF1v8p22tb0zis/LtbViRtA57vTQKv6L
tok7nx0kOgIFtFEjGAF760kld8ruDwuEr9GjCKtv4x8vK2CTmGjuL/q25hx4
9O0JEa//jHVewwcLnf7xgTjWXHphHvIjzYvt7+t8WUap/mYuiZMLRx1mfpxG
ch84jDzPFhYTF9YxJlXQhwOeCW76Uz8SrMdtd6blXOP1zLtpwzG4n8NjNm/v
+D/lWDVj6A8VPe6ZI3IMgiK3peZKKBhpogmeuIGJSNj3sCIexemPKlBotpJM
DaHmracHIGtIKRe6uyz+ELZYrA85XFh/ymBT1giqq6TGFKoZ4R1CMyLX19Ww
VyUxiqKel6ahTdqyUPnPaH7Dmt/xF5Uf/HskJRaXSg7X4OAto2E+vxcvncI/
FIDnkRkyynymQFEQbKkLs+hHNfci1U3G48IpU42KN+a2GKEGzj922kjxL94h
BG6G5GOo+Q1xxoPjqAKdqiwdG4TX6kFzxM+MPL65MRUr0R3WlEfkPhphuFKv
2cPNth7Cst2ZY2KFL4FiVXvSSQagrzvifABixkpSrdveaPkp03NG5YLWFVgT
KrOZJxv84c/yi6VN5Et3Y91+jNv7qxP07w2Jck9oPB+j2lb08f4aoBGCAGXs
pPsdb0eI8RgG//PwTMRlejZILmkj3ZF4rMjpJGdnVGeJ3kUDlEJmOprNjgxW
7skSh6wEbvsojUKJnboeBcqcA/embZYdRlG4FMnwmMJt4Qyp3qZDnusLc6YD
fLMXfB8OTuPhHB1vIP6d9wj4vVRVWZjbyO7UTFlgEqcPR/2kmqoTbakWOKjp
VVyLcaFt1uMDc+d2RxMTfk2u8TLe1ylbTDDfHm4hcLEVG0JBLG1mgL4ZPs7R
zPVYLR7IEOFgHYnhiojL7dS7ixtjoU1J+BCyoGlnYXY+lB779bbXI+WGs8tH
N2pOYRB2/FtqwvhoYItjBjERsmJYm4mkWSqr6yMIhN4h15mOvwYrW2NlGcGj
4vZLMV0i+Z6aX6utyqvRy5pk9n9+vbLcf5yFpednwb+2EeUNHS5KgTTgVKgj
1J8QKex4poZs3YDahvp3JuqsZLjy8c+VamPU+9k8oQ82aCdUYT25ioZaDhP1
hJjH8xuerTix/3yNkS5LKDlQxykakVRhDtx+L7W23uXb/dld9CBoNd2tOZir
1DpsbHs4yOhNfblIfbSapODQXBKLVoRpSFbKsnnERC/9f77jEQuQ2nvNeJix
U63pTydQu4gkS5xYWDrvcKAgiZ1fdjwClXWlLfXAvgE76wSvjGfBvqmxGgUZ
kuKqdmKkgMJwQbW89pfXBHbBGlijYZBVT/lTLAJ74Xq+9knEMs1ynPIjZ5ve
Y1BeD7l2G5xmphZNvyPEIyej9PCGq9XCPyokA01xKGzDtM9FbxHGkAHhv6Go
c4fQPEQkOfRqgHSdRvfKKBvj/aYjhgosXvCnEWmfwwyH1hXkbCWO7uV/hMDB
EPB+dFevBeoPPWCXigF2Sqyfc15A/wwQ0eSEpED+9h+HVt4/Y/vYgd3+NmDu
c9aXy5CLGFJkN+5mfqbwGl15V+G/dEe9VsXKhXWGKUGs6Id2Ew53nkBIxOJr
Wz449l2mAzhs9cNml1s2iDltbnZyr66qbSv36uwNxIsZLlLQ3mLCMVJjchpn
Ua9kTmFkSImzDmUxN2rZbXygUGEEmzS2D5Un8B+bBtwgNo4oRp8p+P2YANMd
NhhC5zqBNK+L4yliUlBxO5leh2kdomiC9rtGcx9m4rnWLetyl0LI8Z+Jt/0z
wH3g7viZQ1M4gL0n4yOdrrWvCv1hE3QwqF2QAOZ2zb55g4Z4/CnbRr6SgEKW
H64e2/gYykwFdq1lhwOvOcPN5IFBtrAguSbPwwNiBuPOu+s/5yH752QLevMW
KiAHU7sWK9hyuZGeoJl3DYg+3SIjixSGKX0irvTyLiZndhjFVL9687Mo23p1
bG8pQwmGzKbR9fz0ZtbhxSyctkvngEPkpoVDjS/Ea4UUsuOx/n5flRm4Ii+J
ioxw8PdLQrsbNO4VHNT19g/2HNZdKeDFgWwnONpXsFlc3eyJNHBcXDXvl2nE
sRcU4u6TVqL3T95KrC4WQ6X6a/BYw+n91zadtSr2N4oCuR7xgbY3oLcbFRV5
doGXKP5zZHQUrVPVpK655vnhlZXqn2qXAzUB2Z0V0sn0doYHls8xfH338pTL
d/bdOFOm1DRu+AndSqdlbaTLgPDP8JQfOGxyqfYiyVYHeJGSilt1d/5rchty
z+/UUzk=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3HCDXTg86NhPu2lfUe37XhIUUP4To9dTHB4ZYrpshVDt3kkGIF9VJKnkRhSP5B/Xe615/pZOdjzO4TaeYkVwOAjLO+E2veRPwV+BpkEm1IGYqtwJmT7pLovVvAiHvR+q5ZQAW7H/+ZA/DMdYbHKAg6ilIllyTJ5pGvz8+jJv/TK1YKI59J1YLlfQzH9RwR1xdJKnYSs9hFq2gMy/NVk1up1OPj2+ieW8X0fCUgHtCFPKJhzNm+I0M1vWGk0p0OAfGXCgXgtSh/dzusxuAVKhO64taKkf4Pq1AxebJbrU7Rqd3PyCtPoNyE8ChZOFNRosUjmx1ll5Gu8U//kBewOaoupBIS8ZF56xjKqoDWSS1GFRGze5P/0ELGAjMIAW4/mWY5PNmqqdP8iAlqKq2idT2FW03orHd1ZjRA+c0VrNEf4smINP36uPLxMfNxgVPN0417l48c/DHt5axPAebIj6Efj5DPXzljVDAlQCOcPaYg7iuC3KyiKMGXJxVi8B2vOX5vlMG0CSgQqYYqgEu5q55MXtC9p9PJuRVD4K/U2frO44fH0Sy1Ysnc+WPssNmxLHPewEuScVlVXRFayZPjRfmAsuhYCDqVV+H9i3Jld9xqLDIHqsexr6gxkdtv/m7E0Z+7RuTnAaxoYlHFqNx2cRz6opnrvcQzUwZ3XzMtbKkHRX9SvWtSXxtWfPQtxmyE6B4lzMjqe8G0+d4lCJq5OMcX1NcE5qvpRExhPLdQySIGVJkiftdf46NaTh+Rp1HxxxNzV5cGnlrncAF0s/AYvnV3G"
`endif