//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qqaiOhAqST5k+Lxv4/sKjm/1wLcjcuQLmvBnaOzHzx3u8nPePyf7Y4xeIWMF
myUzGTDIRl99XTyRpc0g3o31uR4HdLIKLkNTWZXY9RI5CgcKc0iqHSCvGEKn
SY7vtk/AgIZCfUFOWt5bvla7i7iDbtAnLAkRy9bleRdja7hrT+VCvoKphdP7
JT2AMdPAzBe2iWs8ILJUX1YrDQ1xn/kBOhu1OBKEARObB6wWkTZRX04ONeN7
NGP1p6ioswDjuST4Qj1R9fxYHCdWOtX1ISG7ikiF7WZFbuDAGB6FZzaGM7kB
ss0cLJa+HP/srfg/q5M+ta/6TgmfH2zHOcMFUDFvtw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
b28Gz/qtDPIry2i8mUCP5CW/G8DVEtgma17wDVSZ6V3uWNPGU+c01fKy+QWq
63ToUfkZaYs3YHR/cURudCHprmgRrUx/VStUdy83aJBCL21KKILWZaiOQ5gi
g3Jp3RTf4xb8pF5ApNR1xniAslZ3ZEuUdIPfmRxsgdkxeP0EYWQYaIl5S4tS
kDoUzDMz+3toHmpxlhdyldH/WXsFbOQB3hDPuSQzDYY1BH9oO/lC4KTTqYpD
C9URGnEFaykiI0d9BOEQLwyweqYIWzWJ7apoep00NpFbWtuwo+2glunaAd3H
HlitoIK/Vfm4lwuBDY3eUxT3uYwPkqvNUdTw0qQfYQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PMp4CDyWEwYhzwpzoUpeFLBTJiqi+196ZwfoJPGdOiSscY2WGT5wohb0tRVI
UuEaCcR0DrScsL5gXMM5WdHofg0pHg5dsZFdCrISqpF028ygd7cauaebkOm7
/CPX9qc2bqHJdC40mqme3ulMWr9YphJsJP5JBo8GjeqkPc8ymbw0NrcP54zz
uIL0exQoCaBWQLCSQmcKRwHknLZjh+iNPrMPwwCAOKIR7ChIkm2rrQzLZ4Ie
LoBm4Gupopo0LbuY4mohWbNN97TJTShBx6BU9n7T65gZPJe4le36/9Wh83gJ
lyBwOTpBPZvC+9cxVshJ9dbdjhay3U06RJrjHMZ+4w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZYyxjcOcN6+xMQw4ZaJWcAaxpLlgrdIV9UgmAfZLNEllZ5iD+G8JquMriiB4
oqmG9w9hmZaNhSSGzhVmhXRFlSoyBPXbcU2uFMPZaXDuBCSKs1a8t/JuRnwh
KuHxG8znyJAQXQElyf0G3P484VHPtwk0yuuj+wuPEYNM67F0y8M=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Q7C9+uMFnKIze5Y7NexJJ1oYraoSswVsS8uAKzbB91A5i1PvTBPabBzoBJUH
UziEsHRFbWYp//ZTKAHvNKYYpM0CbpqCBt8yrateGlhEoGjo79qvLaQaxDiM
Ib6eJpUyJKnGpiraFjOAOKKp5g5ha9kSobWm9fD3ijyVGd2T4/oFUrWPFbk7
NAx5fePB6XuSlirgyyuT7mM47XxaefAicGSYxQccUOQJx1Q4JNBAGhUDCfbQ
HkZld1qL3XxP9wRL/8w4ZJ/uIimF3OI/7pgxWxjqaM05RPzVLQrBUEP8c91e
qVjhGSD6DIxWXSPM10YMKPEErzbpsyWzQQhTVYdYIZTdgL8v4TsZeWcMEr4C
M0XJlLNHG3I2yweVbaguzo8BXUx4sQuO6hsR3pte8jBV3RR5uqaOkCB/2tq4
qEql44SPauj1R0kTbEBGZgwfA6S/e/ZxoMW134bswxG4Cd/l/34YO6q1CoYA
AadMjGxHcVHVjfITArQRqZqLA2zZ5SGZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Y4IClZbbmR2fjKZL1PIJF+zKSerayYMitPk0whGacZkbuF5kOotsEebUw1Cg
6BowlktMFKUYKnHJmD4n67r1FR62ZA/U39pn8ekaTxpksFxUOBjqNkr4vUuS
CvfK23cQ4PVKaC5+JGmjAHPGp2w/+IK81d9mvOjDsVl8bhz6ZCY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Se6wdrZnQTJ5CJm9WMoJrkfJ0NTH9LcXBS+XiG0c6rgdISWq6D02iDHTd3V6
1Ae07wDJ9XCWpg9f3mA0iruaWkdeSPy2vCjDQV+b9YiFS2BbGwEg1ZO68TFA
D8YKVp/H2Q6COvQ5hQVAjgdJGTrWjKKqkZU+sdW8I4utMAwX7Bg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2064)
`pragma protect data_block
mFoxnYOejA84fZ9+UwO2c7D68eihoYxM/EQzMcs3EYhZS4vf4EPdIGAClFBE
z0pAT5Rt6AOJPHTlfm2DqOkiSFtNk6qX5OLhkq12xzAVlApkdccJKM1G1SP1
+MnQuNs6hq4r2lT71Nid5OYkr9eEZogVyoAikE/BxsQv4sby9JHEJHZ8Vsea
e87EvYUXqGAnCngRr94s62CCkU74VTe8Lt4tA3i6oZcDEiYffaWv3EmRgZN4
y9O2E6CORbqe9+jNw74FrshVmnuQr/l/Dmw/DCxjLly4VMdL+ExlRDjmv56C
q4cpXCF+pjgvx5GQEyBOnQvuoefHj5Hqw2u7oXroZPDDPu6LC3sY6KFz0vok
b0w9gsUsZOC8Vdf7Adt8CbRj2VW/jwUkrI43ISR+Uh7MoH9tzPBvlKggCvuc
MV8mHWUL+ZckeONtqgJWj5mnBsRIlxJoaT9ajOoxO95gq//7+MGy8iHIm07x
+8EHCuWUPnBUh+T1fxHgLjR1Xcf+hetpR6w7y1QynurIOEYNEAnH03rc7M1e
mExZvIONRNjjxW3+jtYXnsfYQmfoZGTBnD8V2TOF0Un334yvRd5o3izQbQoq
oGZKdiMhIBt0RYD3/co6nHBB60T0NwQNMWa96d1dtrdtezU7jjc4r/xNj8VF
pSC75LVsq262ljn0sYA22QWWprUUAHPAANM3ARVENMOx4E4LjKp+yR6Lwddc
3o//JRLBrRkqUn6tsTXKWE8kveaXM24k5FdSNSZCTaXYNa9boUqFE7rcrj1x
w2dDkI4G6c03tv0aZ10LTtpC2D2+KkTAB7yYce40oy+E4iIQBGaLwt+7J1Q3
Qz+9a8RPlPbPC5T04ekWhcGEkrC1Y4DZftqk4OCfDTIo1NXk4DvtJiKadUkZ
1B28cDoSFs/pI5sjR8QfZxt+p2Fl8bhWbGbhQu9fxIzGrlZexZI2mAKW8ynf
rZBatt9J5MdTCpbf4Wig1XRCCogVLniussp1Rq8ZRjPGNR2UdqaPF2meroU7
iFDUAdOG05XHdA+DWKw7MvkL5cWbfM8xt3YVH1+xDs0adF09T3psvmBXXPaZ
BHZZQ/tpBDSQRoGOmrmay3q76w4mXYOSjIc/NqSFWD0MhflaR375LMzbCLEj
REihHo9ItuE+fryIpF3lchmVo614BQt+1LaFXlbzA5zh61J3PWX2XdmJ2wsJ
HKt+NZ6d2envfc17oqJS6abnFLqZekdCMrxFJSmak7XUfy3ARLTKZRv6YjTb
cGc4e65zEcUw0XzHV8RxWshGZk7F5StRQsPAzDKPAK/MDYZkdOf4fyTRWZB4
4AxEykf71XqJBTZJGYnFpy98PsphkJMyoO1enKJM9E3WFjh+0cOX5oU0iKkH
I//qoFkCekNYxFaOopmE0pBkwugq66xw0xTizrZLM/PnSEEozor0TegitN2S
aPrcllVMf/95pmjrWljh4X39Ovt62bjAaAk+ZUzSImpC6t25z45W0iDY81lh
LJUkR2K2w9yRFAYOzHCPQ6EqzZiq3NRfUcRd11Q1N0hn70/AcR+ooSke0ERn
JyYAyDXdUD3LjVh/yOXwjoryc7kLhK0M5sk8OV2g4O6Ib50Gc40CIKo1eioG
3/KXVVJzTNUeghb/+eJTJKRaYK37V/2s50OxVKhFjcEt7ECcHiTO/LbZfnXh
5+92QRrTb33//bOzMadz8xdi+Q8A3dfeHegaQ23+WIwfE5JpH+uDpn8SqT7C
nQ1Ob8gDqMFdA+D0hXPWXvHaUrEZZ5+jMMRT7XCkfo7sSBuhP9RU0eUX+5Xp
8pmXsrjZcuxomX4FBzUrwan7oXZhnlvKCe+cPR9HGvDubqLy01wpq0AjC8Qq
BlABc5ymX421VfaAQlc4A41DkoJ+nkE6OoWp5niFzIxIGH46AXYqshYPfBxZ
Zvd2Muh3mFhqIo1HNdnEoVu3B5u5JO9B6UhuojngfS08pOepTnNLaN3mCpm/
3OQ3ua5lGU52EKlxvzuT8atkA6/YtpAyxGFq/9PM5Ac8EDrewKvO8isDNdMS
ja80w23Zmwij6xhTsO9WNHxBCaX+htbm+R8mESFLRmWOmDjWhMeFArR42oxl
dQOt3VL6qFO/HvIsmPfhz4XQLxHQ4V5bNpIkVVPYuQTLNKaEhcvdp+0Q8/S3
VyvEI/HTGpMHHNrHmlFFmlUDZKr4J2YqUD4IrVz/hzjMEOQzcv6YaY6HZdsg
XEORT9NEDmqXhaIYckWdLAnoCluW35nhce8YRxZIPb4/X8d4VWaT5UW881nU
OEKBfAo2NOcB+8CC7VOsI+qsooZTgXKsM0jTJFcdqlKKqCjyT44p4EmZsT2F
fORhwveD3tr/8vqKlqgxOoDXHAvQ1VQ6xMwouPFZQ/9ikhJS/eDBkOEDWMSr
stk+PX5c5oc89VbGa/7PT0IGa8NjS//EWdywDWZKkoLmsH7oq0dLqhQLo6zD
xU9RXhgdr5dkdqttg0G3AM6REpN4bWKyiPWAMk+YiizzGG8UKBgjXnt3WFd+
boSH11/Slu8S89p6DhWmUHIvB07DKGDwmqkxhSzD3akkTBB4f8/AWO2aimuj
hN62GqZbANuiIce9mnkm8HNFsSMXW3tVKfZphoZNGJ+kB1MYjvWiW4QKDlYT
5VpoS12/x1QGgIlwICxYB2UIchOoTHH4CqcA7/p/U5pvlH1nRBz0M+GKNJFv
W1jyQcTXEAWFPTWWNWBtTGKMWlpDHvEInyPMfNUJgCt8dRLXhzyM

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+njU5pMiV0JsCI939s752OBIRzxCwUVSP9uZZ2C/hSv10M3aQJW7MaxcfJkgdPKeudP0mir4U+KK5OJYjAu+j282XXzuo6M/+prBSFwYdjER0F9aT850k22OK0SAOJRu8aPKuNct8LKEKoFIcIZXbtPWBHnYQ5YoTY48wXRHqrH6zYU1mWK0fuT30ilyIikzyMDfiFRumbR2VYHQl9N3DOXxYy6aGo5eravqbgd8AXFWlloKtlTZNypydzwd8+N4GxKH+KX+Y5wRPuhhBdMY/1pa3hf/vH+MTU4R+cn9VHo9RyVWUDyxsfvtZYzOBONzUUWi9RZIYOKMx/vDDTvLzJWyuwAU0eYsYaQMInFgwQDz6bJ+719nMqQDo31Px1GUZRBidjSrfpPT2v1Si4yj10N3dLFBjxVkGEH+xzdyPGtl0avXbku1hCHihtYSHBqWjl0N9l2Nm9Vtw1MUrqvQHYZZYq+pFIXife8auFeCNr9xlFMKXdR1l5Yo47+WZqcnk1ZCKrxW+UcPzhGhlkgNFesXun9G+dfjLlHOJrKIskGAmdZw2OnsRatFwlCzAnc4rngYXCPFFnV42RVLAlUae1qQz1VjXnxwUqyG8gVJiuNrtRKZFfUX2TSaAysZAI3QI6+xpFdEHfsfGufnvjRDMB4lRCnIK5x8+SqOArEBTizfvIkcjzVkUTzsgERtSyvpju48Ac3B+Ab9Vn3LQcdYbPOz0sYCVt4lzuSHhIdBmW27T6AOOAmkiB4Umn7f71+RYAX02um/XBVOFGaan4Mxfz8"
`endif