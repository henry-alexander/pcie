// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
w0If4EzlH8vInB83VMCzHyHt1jIgZy29PrgwhDTgOAw2aEAsIp2VOokG0jTr
Z/O9PjBReuoQNsAQjF3vsXkfxWDvV8ReSE4uAbQT3dmDC5M1CB/HdtTX8QRU
aBZBCNkWg58sYXoUejtjnxar6QsP1Dmo10TbzvLAvQvwr19tysF285gG0WsI
9U5dxw2PSNt1KFNsOv79RQIZEqqzTZoNj4z13OpjydiC6fnPx7JkGTvxyNHR
OenXY0thsN5sXbAQkW329Znu9DcY2AeOLdk8Uie7KerPGA5Lv+THAgTJWxSF
s/gvlwRr/24F/cGqsmWfoLjHTCrOMIpUC3DMg2jImw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
P2HNHG2Hprw9pedA7vFx7cHk5+K33rerR7jI9vYvQsOk1aauNYUOE6Lfc3AS
tluzqomk5fz0YzLbIGmMiW6f4vuRORoqRGvx2i7ljlvzOl7NS1R9RjQnmTxI
+mlBlcEgqAABQ2ulL2CAnp5ZL9v4GOqxjQ1ZuPbI9/gtFaP1yenG58u7BvDG
UKBjQ/xssQZG+7REvhbE4q2ZvA5EDbmLCh5RE3LuC9SYWd5Rk/q7kz/e0Qtu
K6xBMCStfeX9q/vdPpcckw+Lyi+A0Amly5ski/I+z92fcDZUKQZC75GOK0aC
8uzWqpim+fcTZZc7m1oLbr24DoM57UGuNZD5pGzTOw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LyQlS5I+dQTFEP4bIp0dlRWabFsRbaADnLfv+fQiUYLIY0Xkps6wJWL/KBv4
gnrUwcqwF7uFZeqMVMJtGEwEnfIVuYH5qIF9wcj8tAJWieaAHk+BVIbBGaQ4
vuFSqqpGkf/JBvrkiypVJaC8vMjZ8miTplbGriGV5b6vbS+4VyFyV0W3hFoE
atireVTmKygFKWd6u4XISEaBHVlH6pLwnvUkmBz8LoPF8qzjogOumZqwyN2X
97hjkqoR5gPCAcrjqVvhsOV2hAbq36R1j5I/A10pC3Wj3UA44bqNq4ClBJNn
zthzHSTEkgaJ5cD46Wv/X+JlL7JQe3yjbzhAoWDuzQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pq8/mJVfxRC/KaUC3i/+Ir75NrwX3nPFHGviQbdWnW/+sFrprBibP2u1bP3r
Arzo8yUdTGtH7rD1eq1XgvMILL9FKylKUN7vdVmPomDBrjwKbhseME4mBBk2
/MksjKppouVKpyNXC12rgd0/M/2IwLenjKX8Kyqd/gGvux6EMQY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GdwSmsSt3OFA+qqEs1enltP4mtfCsvY4wX69mt3vYu9BI3VbVzN3HFsRWkGV
XG2upFPKBU2/xNu86NWK2WCGh98RJjVVX1XT1ZudwjS+LwhfkZHM0vaslXz3
XPIEHvJMZiQSkbqi9sYCBLAMCzoNBznhqVBrVrIRKFEj+bJKKJjIHPdoypdR
Q05552OGgqHQ1HYS2DjhuSu3m9YLpwoBHOp6svjgbOPO5AFzmV0K8xyV4S/I
/bLy5sCzYNAn78LBpi/HmJLfNztcKk2DDkspNx6fDpbcvPiSxUwMi+SJzehv
MKj+660dqUYM+AjGIn3fNp/0e6ikJdPsKjQjFrZ9xIcrmcbHMljqqTN7MyZ3
3g38cvv9JXyx0yR3uP5xw2Hd0CjfzUNbkMXAqtL/n4bGOfPXiSvluTqU9A27
Y8UYWyJWv6o6kJtBxpGNtdS50cuKAxdeK4s+ZcdRH7ci9DxNYlcu5YTDFSkJ
vq11qlp/D6kkbOZVd9W6BJkOnBLB4SHZ


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a2vt5WmvyY3+ZOlf4h4s5IIRdQshP1XHQcY2CwrsDyGQKiVUY3UGsjMNgYco
rpNXBwcpYk24KyID9w0S7YVySkkXB7xAuFAHyaSWLGBxfk+zRT2AXIN2kGhL
7Dck12ibIu9yoGFQHya58xrgvLqcMsDWbmcxaxmc9tfSuaA66Ms=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ORXZrtjplbzw5dYhs5L5VcJerHnG4diG3EW2pcg5w9wSIX32fqYPHSmcINJu
2pY2wYjmOvIkwUqS3YxjYyxb8XFYCzrlVGZ/dhB9mjNMXedyQPmz5R5pvUFj
rf9cTx8f1mgqeaNTSB/fu4YG+oPw4f0vlgzSHcQM3p1cA9KIO68=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1600)
`pragma protect data_block
oc4f4CeMQF2AHd3WEvErB8VQrfVTE/eotuw/ec3PBex/dkHOIyjX0pkUXHeO
NQZQvLkVZHXp1Zv+XFcNrOPzh+wCzrejSfOqmouRsQ2Z0k60ac8Nnwhk+5pI
swHn4oFdI83gTn6/E+HYQzHdnkejD0XSP2GviWtkMTt/c6szlQ9mBoiYKqEa
m07TKCY3TSkn/s0HeR6piiR5k9kQDmqXua/ffH3W0H3RTZrIsg2fas4KU54N
uOJ1G4KnAB3iXg4lAIxvoU1aP4DgBYCew5cQ0/QupADke88K/Q/A8d1NvIoA
LhBz1APmQ25K4y8qwcGlfqH5cYFZd+23AoaKp7y79MxpRMFdzZ/3JnVUHGI+
lloV+Qptjzdj+u6eIexMyXwED8pOQXLWpgQpk640nDiO+48q6PYr4lLyLKRE
MLvSccL+HZJ49pNcYT+COBdE1BM06CfK8dkOkrGnN/ufpcdtdEWADtc1KtRd
3jpgqYMotccn5nXLh9AquaG9nTfY0aH6AE3joVX1Nh5b8wZd8sMRO3r1tVdS
UZGMcsPdXcZxIk11aJPOwBYiIlGs0caDcbeyxAsHUqEJ6i1u2PMSMQ++UN0x
4pj8DOJ/4zU2jeK681qWdA8QO+m18N6CcWHhvO3DW+7SmZQXjncwgC5CXvK9
hZFP6pZ6CHrC7ZLxIzexao2nc8VeoU6jP6dLtFqcvES4I7dIdqkfbXIco4Wf
qAjHRxe2LIoFXXh4j/XLIJaATP8StPSyAzBuxjWcFuwbwHvbmQJ8Ly2NutVd
ao1bO4/E0AYMD+gBaLqL2aocarb7VNvODypZqM0/izgRoraaygElrd2XLUog
ibAeukyJpAMlTypuGpDGL9AjWdpOGadbAyazil0zUtakgDYWgs6lnlnwTx1b
EkpxHcr6OSAmuk25O6DzLsNgm4dDY5DliEFFqYaowc0r2YLla7NeWVDEiC/G
jsCNk2FGWPnxdCKruH7DE0MVjggE7RhWiiuoY9n/p7ZXl1ZGxbvDExVjiv1c
s5r8BBcj6YMauYBMwLkt/emVyV+S0nm7+1q+3S45MSo+DHbX/U0HpLB4x3Fv
uMZrVNYgZV8TlfLTD4wR78zdC9++/eQ/iqIJSCvmxx/vq+uu9oS/7pGcnSfz
agFjxKarbuZxVGB0eA4DvbqSgC2h6e97qRh0htuD+IP/rx/OyC6ivFIL9YlO
aShxRYUabnxeuMMYNnlBW7CwLHarTF/g+vjtxd6/Se6ExdxFICZibGvumM1E
X312HqTtF0xnmTuSwYLgyLR0bH4TJgF7UENtkgTE3dGunJ2qsbstAVNV+Yyg
r29K8uZw5CYJ3FfL85yThGqLKR5CaHXNri3M8rVVoic6ysVsY2H1vmbwV1HB
CKLW7bUcbw2/9BqCXWpKzJuwdvJCY0XEMMh7evQqrIgGoK3d2IktGQCn8iZd
pYBQcZBdaND3ueiRHYAkY2ShmA9GrvvQXzje2FbOV3C/7sMVstIAsyMD7szZ
Xv7bWAagA2gh5rhSjZtozGTH8B3WMb8h3eGiwSmRMxJ+5dSgKzBzWzz9oSRk
4T7IE9p7zvPZQ4n1j/xXbTsGEBqZprH35vc6vChund/K9IFelCFgc4bDeKus
QU5aeg31+RbiDIJ4FOH82sCO4HkPJ/42cKiNtO7wcZUlAYQ/lF0rDYLA7DSe
Svz5s0m2mpzGAK8SBaYkDE0IjZEpGH7bjcrZtFLQCAN2CfcKUUYdm2rwZKwe
L/ADTyK7/PE6IznsvqdORoeVLsTu3kH5XPnsvRWMAqySb4cnqeB8DvCr8It5
A+r3JJJ3F8KGLi7rJcwCec6bjYEmKHQyPet0W4ZIhPqMpLgJH7dSHMRuxs/D
RtSR4p4Frs/ga9oVmJlPQQ4wNY71tURZs9ZxP+jN/oeuN/mDlFTBaZ7aIrf8
DQBqe4NXCjp9aM8b1JU3SRA5lLX7w/5Rjxg5fgdl3a3PKCC42jJeFBz9IFD6
PwC4tV987ciD5qJ0ieGIIhXXmZ87NqL1E4XO4LhMVB7SpsCNblSZ9XXCAi4Z
6rIKjZL5ZaWKjGkuhbtNVDK8BnkjlHxGUmY7AR8g5d9PdHRj3EIF0p8Y7SRx
8mT8XiDlVUruXKu1t56HR5hNTzUoa2fmrw==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q4aPi6Jx+4K2Fl+iv9idQcMd//X33Z5BTVcGY93VH1hSUnwkP19bMRoCUFpAxwj9hjhBIIXhTiviMxIPX6EhhdffWkcRMb4t3TCqdwbnSNJT/9ep2GVQUsSYau+d95hXeUshF3YsLLW4t/1hUUSaFhdTA0EhYKX7iaQ0oBWqyWiR/5iQVzciQLiV87lfy0iHHuQ8GswdVvjpdN4JZvofaI0HG6dZYZnTA/7i+RZPICC1mwkTpFB8lD/Q0tvEMHUwuEaHj3Z7jEyDvrD4zYF4JOvdzU6CP5I9NoIS64dRh2Fk7QEVhWsmTMWtypXr/Wz15EVtJ/Wx7XuTz1MNFFWPivFxcPD+kJ5lyJWgaQZAT55mKMKsMjxVRCAI9bMZih07Bc3cAJNLfNDhzBMfkZXAehMl71WabRFN5eP4zVQUwAvAGsxa5wd/TG2beuXIbhoVF+6XSLbtcn9FoXDvkAqhzJ0zgGj+NDyY0AtPj1N3ZgxO3KxlCFDt3QS2OmHLglxRqyOKTHNtpKjkZaXPIC1WqV6t4TqY88G0paWAxdhTWUNFQmOYFq188pP/ubs2rysZy5wDZe04Z1bvLXzLtJFhXWbiPxJZ1u6exz0z3x/Ygm8ILD64jxLZNsdURkuVssz6TWyGMfWKUvibCJ/WJRCB/Klf3EWYawW+4Xyy6cWcwIjz5n/d7ucsezViZAHCz732EZHtY1xHOjJ9L2bsJy7f5T/ixyxeR5Wowa87F7B2X8o4NlQBqCRteQi+E8nRXG+h83eZoBFKOqmk6uF8Hl5YeYM"
`endif