//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pccljH1T98+Ns63PtDoWm1PVCzQ7t10+Q4Pjp7eJVPg6gwUP1UEgA8kP6QdK
/eLYgrLCNuScWFxbnlidz7gbVd7IciPz2F497VwC1vjZxuJqVoqwzR29hekp
/l9cGrgl/0h1TsKRsBufJorfLpUCt/o42bmTZgpxHrSBQeu3rZe+HwHfvY9E
TjBRiF9gJHJxfXLMKECfoiy64YW8WvH3V8e4/95tFYiDzJCLHFX+jciBDMRp
XeSIDA/JQKC2+Lc4pDkhOHPoBjpZEgvIJwV8wmut0XF+NkoVY2Cu3XXmsLYB
gXto3EVTdk5GVGGAsfU8NV3XGMY+t6MuY7AQ/HyGaQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
MWjUkbB7PzfZ4GQ3Y/EKN+lz6sy1UDxPGfytgWn5hRyF/+BfFmz9rRZzDVip
Gs2h1pHWh8mQ4SuXWdKzynSLhgwYKyFqHTj+H+hJs5v+SF+uE2p9B8T1zGBP
HnMgyMu8W9mbyUAsSEpjhMoNIG/OoBcAsdvIZryqNSsOYn6DiQl4m5RFbbk/
6R2K/VBx41cbRpT1jJo1wU1m/awQyRzvNZIKd3X1Iu1icPSwphyq6bzONvZD
XHftx/4hAi+GA7ZOaOQNwpvGrIa/7AbjVtlXqDVgHfxRaiKqMfo28sRdqepW
RMvH5JmmsNqre77aYTNFg4Pp9KfOn4215otYbqRdxA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
J0P69+iZliagxVBQP3nNdmQ3WVfnISlc7j15VdPk9xQuve/q9H0pFk4nLU2t
kkpGh1uPx/VK7ly0iiHU9CIvDA2S+sEBfo/zopTiMGXYu1yjlGPo6zYqQek2
BfB3zZBIeGC9ys3sw64WZMvwC1l1Ze3g4xEvi8/UrdWov/Em31Z1JXeB9alm
4cHFBmJRnqWiyKwY48yeY8PPTAOZVpW53XFrXDeNnmNAV8TXZDGY0z+AplIY
WcEQGWRJfxkFn29Fx7+v06ffcbPcnxujVT5JGugBktvXSnbKi2/SchCtyZxY
hLxqP2wSjSGTNd8MYk4FkddSGdjZjCYXKCmzG00mRQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Fuy3QB8hJGks7gcUZfgPdFkxnj98+/KqYI1EK2/cflNMQoTbpN1Hz3QAATZc
8F8J/qLSNYK1mxXkTx5SNC36tq4dWbKQXEFQ1KR01YrCsK5eW7F9nc3aSZKV
42tYmyj9PK0EcYsEDx9F40ucvMUfxIWhSo6mCCzSivEe3pMuUAg=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
LvspQpfmA9mfVjLGPVKYMfDNyCKMZFcYIR9kX073gPYVcKB+Q43xlhOAf1od
gTlKlR6vb4AIjXdvlQPHAY92ilxAqyXxftPnxgJGrVJBQQvBGYei4GP/h/S3
FhDuGJi2ugLtKFrwJ1QfO3VVsmZABT6vpyY/9SXhSQGbMu5c/A1oxk07Dt3G
wVjPzUgmw/7dorwlQ8nKvDL6rHEYG2HOzOrLBQnblKrnDuRRsio4A2s2jT93
HjVwCDKxk4dMXAr/hO0Z+4hbEDRoplMDMKdcqrazDzQ6w2XImopkhLEeDq6L
J7E40IUXcTYnP6Uja9bPWvVhzucL7DWlfxY8jIualqU3VLwMgu1Jz7iwC1se
XQup5Ik70alAN9XXP4zwMI/F4H28EfY8+CqilMfo3bC3Mje29VWKCiPIIko1
C9d68eqz5/Fg6yQxrv2rTrFLKjvypUCgBs1HhafVuBseCEJ9vQsRhVJShq5O
R7Tp08VHwqu3cU50wjae/ioI8fMSH+h3


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KAnmZqssO7h10xV1728r8vB1W/yUZe7V8EXV4PYvKFKDoIhyHVAHAd2Zodoz
nZRbO3xb4bSMcF+f7bKO8bRCmj3XOKi6e6T+TYzend9KcY+2LKehJ9OBfrL8
Blwt9AXKa4GVANC0l82itkE58R5vCGsWC4bFwhdGKSaL2hA5W+E=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RaF4oTfYxEw1vwez9vpvDhxsNDD5Cy096vHp0kT1NprJD+AUitNw4hPXIHfu
recqLenCkEM45LQlThRrQ414iaeLQY91UCq1Zj3Fv70RsNMg/C6uOa9/ao0q
DQ639KIZH4zToXG+DCLz5z3cn2b1RUjNQYXot8kwUwO3rqCSqB0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2672)
`pragma protect data_block
Up6XyBp59Q3CcNudw9siUZCQZ1ud6tFpZf20+y7oUjcDIs2CTGek8PwClz1i
tahBoFIYHQMjn/pBxv5tpg5yiZWwxT9SKSmRKrsZlfiZ2+jhZDfVz2kBhgAE
5r3qeBcWdx9QAEo9AldCyEI26Y+lC0fPY20Fo3/ieXKPAR7uzarPbrI7Eh2d
Aq0hMcspcwDUJBZncGN0H9AZGRTmObuYwGxE3C+NWi1EEWhPThBHB/w8wN32
uN0USIeuuDAW4e2seTNXJE6v/tvTvG4I3ce8mci+0L8fijKCUehowbqclCUP
D4FCAI0YsJHeK8sk3aSEqQ1mlX1+hk54xuL6zkQQCmhDVRxRdmMzCEdNcRmT
Wi1fCHFGVP/5sxBXw49VYZPv+z4Nc7lTdjiK2Ww12xfh4+TBMo0w45gVDqh0
TfFi79p3hlCnjtIWPecnL30FMA3wCiEoV0G2cyOY6wCFXNR5Tm3huznjFt+j
JqM4LggIBiU/3yas6tSRRzUCv6A/UuQ9n6Vae3X4iwaBjee1KhSDZbIhI3NY
Nag0dSF+CTWFg/1yXHNZYVFlAiuNqHSGiMeKtr4G8qUHKuR7C5Mg68h3OfJ8
HLTPQxhwS6pa8v/H2+jIv7ijCZ4hefZ/wa+atGeODZX4zwlUh62UqTuNhmiU
lj3q3VsYmRtWpXlSlmF4qDpLRJd/vMKtM9YYmrZXgqSe8mMZeIVBGArFTNxS
EGGoREviaMhlzEt8w/26IVBI1xPTqjFSPlkhrd/zcCespp/RVKPzhTr1SIdY
58k3LM3+8ILiGgcABuu9evzK3DlwuIcgnyFi76om42RRIV+8OLosTVFHafP8
kPx59y9glsVl7070IwmwBAVRf1XSQXCl/TU7JKpKdfOkfYQy6yjaDUMzYiPy
xKGwsj6fx7LyWW5czF+3rvUSbqOo7k0rfsukf7xMvVHdUzl6c8OcMGpqIf1S
NqSlw8dvyC+Y8h4XUYCRPKN0bNQavVbwDR5nUdBKeoNYCygiHf06pBN7gXQD
WGXHtdWu7SVyDgihbHjtKE9eQb8t8nvnpvzSipKcCBGzfjOMCO8QVMyAwQ7M
qSQRKhWpV9NwqjlW2QbdKaamCS36UVzintSoQNHBnGM/9qz4prAcfBhwi9mm
iUqA5QkCKVA94jGw36S23PSv819yVh1BWfcBbuKwU2YBSZP6HB83jh2O2RgL
vyoL/Zy6CzEScgf29SUr0UEpEs1hNJH150t1cbFTSJweqgTbhO2HznyNv4ug
lvvUK8fuhCNR4QcAl+bgxWucilaozuulvyrFYE6S2o+M2dlziAS1p1agATHY
SqJh3IXBC/st+bXHQ82weDRlBEirAGwFHeKi+QTJVYdjWef1al8ZteWALbhU
8SWmIooaBnL1VlXyRNkHfNb9JUOcCXwoDPRtefKWmxupBeDAWfKdtY2jAbsH
aD+qYz+kSqX1W2s0WZrs+IsPPBLI6522+DpoOJlMbZfJ44y6e79BUyOSge7M
osP3wCdw6DNll5pkX7ynKBNs/tpQqhUYHrUY8MOqV42dqU4he2/FUt8YCPNu
FphQgSKXGOoPnqLc8wg4deFm3Qfp2xucq5aBZhKButD83/2naPKs4wFeWQSV
TMC2fCtDXdF1QNRygu4qTTjjWJYYBH+hINhFqXoGQhrNsdiHexoqRTKewCRE
jUSBQcy9CGnWjqqI2N3Ein+eL6/q8jHHyX+T/4sYOGaUjfu2zcpnDMUaXfzR
mzmQdC3bokWg8XYuT+aJ2ojRS8SrusR9i5loVwpT7sg0e4+0ATJaios1iGiT
3Jqf+v+Bsn7lkguFebiPSoQKsX7eOdvPPr96grU6f/Wqt2Sa6AzxsTha2sVX
680Hm7sbsp9h+hrLvn7aB7UJrjQ3AnD7FwnF6dYR0snsUCM150HmH1t5LByf
TgivdyXm5IowZMC+coZNJg6RK/G6cBnumPns64//k6tN7ODnsvuBBBBlvfYy
gC14FyaaKaIgSzm2aj/XfJ2xebDn+xtnMo2QR/IEa+HOzxEhCm8ZSphxpT3c
4yaZJksOj60cTzEN7a+VxIjAGBAF82w6dDUn/ZO+jMdj9n+fTk7BGZGn4NGl
kzGnYkg1qqt5rk6huCABXfydxxDbFLcZxeV3Zx8AxausNP3+kkmNI0IzrD9D
OlCbDxkR6Al5lDR9eAmmYcohKs4D5CxEoGOd9NgdNzW/7cUnEkE6TV7bax80
Wf1VqQc/fzvHmD9438oJninPZTpK/3YKn90UAHSBN6Lr7FHY5NZcpzr/OACP
y2Sa/nyAJGr6KxzghAyTyZo1jGqIHYQ7zG2Hl5iV6MrGanisIjGi9JgxMnaC
eAgQc/vBodREDbaTz4u2n/Sj/qc1QnthcwiXJGz1Xsp1PCEg6kQuDxOGLmI/
4yZD4+4v6NZBgsQjojEIfsD6bWCJENryej4ZpxKBc1Dsa67LUsc+iogbAPIC
QFR4+/xJBHPQ0s3CfOwbOPb3ulOMjPjai4FGkVBktdaxKK420eNWV2mOzAJj
xWiUbb4rfKIfnez79TCGxhoF0rVCSK257FmgXK94l/ZhpooHCOe4ITwR2GWX
ThliyUzlP7kZhm/DacpV3SQ3TrXMxrjwsN9frMPdsA2qkmcvc+BWNdn5ZAHy
44me7SxEJzTs01vDDlTA4Ly11px1D41H8j/HojxNeMWiPe7sEyYtsldBLJsn
00Nt88F/6AVstWvOZlx6nrBlbe2x/UiDuL85TrMa6/5kPGMlkCHHsRiC1Tcg
3v4aKfuvdJwO8gDG0/YmUBfN6foWBMQslxOseytHtSnNcTcr4ehW9Z90S4NG
KhGwJt3mH9+n3dCv+enugYAd07Bc/ozFfXGaqNQ8IK6YIFQyK0INUWKq17Am
tlE68SODvjHfpwkcPkDEacnBrFhTy5ZflCjvNsCBKWJU7ZbIabAuX9L3vcZ5
giNm4ANjtU/IQkSCrOSV2sy1S2atIUCJ5cEA2AMOfI2trOfgjjIbT//5mRuT
YJclAlWy5kO5u4ZWpA9C8r5uvs6Y/qzzGijZAj9OSVz0NUrKYFUY7wUuqj7s
pfipEGtkGKs18qaGuWbZekGkdT+rhLiPXwkudp5BkEVKvgwLb9GUPFx/VmAX
3AB+WnpLtEbmRO7d+HJKdcj4pWrBs+AvbxvtkPSQzLaXHuV+AWw7HDfBJyFo
F++NBekC6DzcGam8bwFOd7feTQo4FRm4Mm9rKJlkNqDbOE2EhAjZ0a4Aomd3
L3S0JQ9hmHrFwLAKouhziDO2cT+nlwqzQt6vOG24s/rH6o5hTS17ru2HXDLU
SRq/DzSp/tHOImDNiPqIJ+HF2A9/lH0WERu7+8scjvGDoAtg6Qg4Kd4+7nnw
XJOpZJO5r7c34id6RYF6E/r3CRlEj4moilZyeVn2aJz+EmJlR5hbQtT5sptr
e+6F5O5IgcQuyVPrIe34Pjw3K6EhKJX1Na0IEGlHJtkjgW4GKkQNZ+emNbhA
qeVLIvBpw/Qa6JoVR3P0AsfJZoUlQmjJ1Mq3nxQVh2Tc5KX4CRgIhusjdEjw
0SDflIE3Et+eqsV7J5WlI6I=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+mBSUAt5WWWqrPzXRBhRGpGeJXfL5UYrPRR/fzJ3TTYC6hH1LIePJ167hyWdFl+URTdLvxLvHqIFH4JyQNjHhnYcYAbN1Tzz1/BYn/N0/nnRhiHw3L6SXub2KGKApsWqTKqyxKC0+gm7VAnwL85CH92OjgaQj7Guwxq3QG6d7f8uXb/1gO4+z5GoCRnGLhws7t8WKs9hkp3FDMvFnTtnhhu7EBhlVg9x5xVecGjYQSvB5c5QWHACTinZfZbrJTLCRspUR47IEMKBAwW/JjgsbWOkOdy5ZcKRTsnJVk6jcX/pLMVyPxtHYmwUMbJo58Xpg9iv9ZIHmJEZM6MyCHn3tcz8se4Rv365Zr9ftb/ZaXRZa7t37lIqhTpAfmNd+0MbjaHL2ZDwNKxZbaiwt4k11z4rWg0kfFqWcX10wwv/aMbCHdFhg4O/cpFVK+sOrxxMl7HR0b5bIO+cUzV7MBu/LaM1bRvO7iN4KUUU0ynPepzylFwLo+TD2lHlFL9NTPNTindVwF7E8rfFgoSA8GhMcodq/RMH5uQOS2HtqW40VbaeqkRqkhQQWNBB9KBi1e2J+z1bWP8Uf6JUUuXoTfylhhxv0al4j05wwrRWHLTcueEfTdOQj8MVE1RhSAzNQ0K4fFEFlkQNw7W34rsobCGg3nMGYZU0QKyWnlLj1cxwUvKTo2zlCMtYqSyHgEc5kZIMyyikXZ3YtOn+3A9NU67QqEXuMn4TE0DWs6QbUGNjYI/6pyYRjJd0DNCwmoySeynrWeZOIY2ybTsTxMSX6tO6NO0"
`endif