// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nBst0MtygoAlYpv+mrQ/Nm3k4pNlpNWqVD/bz8vURVeTkdS0lImhBSya9VYa
OMXF3yU0erfoc31SeqG0knzCyH3NLN+HhlA273qHZL3uH2tWBnWhVpE7Kwhn
z7ENJNwpOb1k9BXk+E5k8xU28Ueo7sT4VEelQjcrL6Y95aMLv16xAOHGUxZW
058A3b/vT/dnEAYkCglhzLgYTZNiUnwT6R09e4k8r3XgrMWXXz+FIcuBsyzE
cTQBJ5VQcPvK8MRjg724PtcbDvy9/HHjQRHiidhKzcIOD3Ex4I4yhOQb3/Y1
DSuOAdhpvgwb+/2WVjhbUyvcBUM01G4xq2Ef1CIR2A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
TD4KNNhNu4aATIpIk8HuGwIc/WEvfN61t6BVzK4Hhu5+qV8bTCDWAqmBAk7E
IBK6vc0HJAPvLBJKHNwpwQ7hT8c+pMPK9i60DGK4zTV24RyizigyNxjnNDo7
vfw2MfBSdU+IongrdK0cACGhAZRPHXjYfvHfaBARbvFxqwV8zJHfFn3OBQ1j
eGI2x+66fg8iTHeKg5kaMFmYn8Ycm88jE8kiQFqd0nZL3beFqBwM6E3b1acy
sS7VxZx8FtSPsLknyMykrWdabkQSa5JBRLZd6zNLOFnTv+cQiASvWx24Uf+d
w5qBeTEwUyMFrnQTtD5APgz1EKAOXKTwuSy3eqTL/w==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
A3X2Wf2hFld7WDGqAZkqeUTaGtMqjD13TaWKaTIPkVTdirwz79koItZaCY/+
EXKgfP4RQi1G2jqzUlQQrITY7q6vMmjEAxJ/S6Ma2Wyk7nyrtUz32qv/PELU
yCXtL3Yku8j+M4hc2GGHDSB1EYZ9/nbkL8FSnWDpwo01+thU2NLkFfU/0n7W
pJhswnCf5LL2JPBve6+BFPv9gutPeouKgyBkYk0OCYl2N8hb7JO/QZy2G+j8
WM/RfqFLzlFIHhAI4rkAxz5K2vjicJX14KBvB28uyB9D7CzsHHaDGvzXTR+m
5AKlB3ZawSJBJvggPIfE8VINy73wIVBGT2u/iyBdRg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
alwtSC2CsWBPd8QkgSkwyjGTpV7i+GZuaBlsHDohjjlXqVT8mYnW9JZOK1xd
4AGY+53QZ0O4i7VhSOMwCO9WYfGutJEPImSxmzrRwEMZVDdOHuUHU/v7q4P3
IgnU1pD736c7oJRg7OPaad7P3+hkqYWr3Nqv1xkm+IbesM8prs8=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
syxnFzgQTGsAntsJJBj1vL1DXuosg4XV45mMNcXa/00o+8uBfMqoH3SWWcbX
T2uXHPZwufX+bnehFJ0T8nus11FOWJC1uaW4TQvrJEWLiBYDPxf33zCAuyne
himXrRdxYUkirywuewKf0eVwotEL4fyqEm9jWTgcae2msAKoGHoXso50xPmO
kxiNlWDyzKxRXlHUEMfRSUcP6uoN3zuu4fgqCBeBbB6ZLRy0S+ESEDowqdBH
iBiFcUu60InM7YUMIUuL1dlp9zuK7wMb87Ye4u1kTlC656jjqtWs+qgxm2R+
dzPvBMfGqMuyHjrxHtGRMIyPr/XexCO7xbQ0pZf4+tYtK84igI8oFslCQ0aT
+vWrbHnNCZjzc0sndQZBunncdYS1X/g90UiJKT+yKEY6XfCBiXZLw5dfkUrI
MDUE/nPjmuIxH3uvi8139dYwIW1Av8NLPjdjBN288zHrXWJWv7HI1fvvNw3F
qOc+rNSGxfdwV2WoyN3FWIG1v7yy1P3M


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
BirqyK6Si/FvBocTtgKAPz1CK7AJg1SLD9HH4dqC7B7o3valt8FPwuRMgnwO
R1wEzdcydDxWPtSeFqwDBlb389g329lH3RHVwHHuHhzewLY7h4nKNWSI2irW
LzW/pjyvS1XhSIGqw7vIJCvJfEfozfD+FTJM05eqiw7MAlvm7t0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VlmhyJ0c5/1bpKAwsZJJ4dZOwrDs9rMhaFPL68mqLe7rM7/WOZDQhO7PjWoO
a3z2MK0IAYinnnw6N+EvIE6JRZZ4+mdwqlmfjMwuF/oTnnA5Aj7hD3CVKKiB
Tq/FWjTRjU58Afnwt5OlhwlXKbG+svgiYCmbyPmZpNV9jZ/jjwc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 100816)
`pragma protect data_block
o98XRJaAbe/2n+18/mqEKBda5ZduqaipEfHELJDNW6etZb9YCHqe0T0CdEi6
iEEx+twwDZUNWcJ1s1Axa/7oWktaT2P7EnMZi/dqNtKxiotizxAyXEXj/9hd
+nK6YdYti5UmTewtWW3Hb8nkn4gX2IguSB3oa9fgqVO4HnK+dkR1w7uWMGmJ
23jySvRf/yf8Hl8HQ5/yvXkGFqJL2sTHQczTSqEM4j2cRvd/DLeYcy4nBXii
ldgvLuxezlO6R3EqlEZs5RtdZmGWJ+x1HqdxC5ziLnBVJR7YgKnepq9OlX6w
kXuT4nCcduuVMX2rSsxpu12pdhXZqcQ/Lu1XxONSMAL3jVPCOt3aVfHhHxpv
Ocs0wYdhIoXx9R8/qTrIr0DqupPfk6ebYV1+an38pdIIvLwkVkK/aPSq2Ghh
pmNbkK90LvrxIohlOKveaPZqRpiGzf4swjV3cFzYe5mk/4y3fBoqnukRuVGx
0/m6NvCuzdVlnsSrBbhbBOMM3e441OTpVlCoj2LWeFzj8zcIgDEOVhn6q/kR
ff2lmYcTjd0Lliq81G83xB5YRHcPS4MN2/cJosCazQq7nZt/RRoon7+wgPlM
4htpyFl37Nk/rzSrpn0j+37GyfIRvpbZ7DwkH1TMnedTZGTqVTq+bdLC/VkV
q9OvCbXAmjJisYLpCM6RAHrlXYvcZkohH+Bmd7nxAOWw1vaHpOxLXsJnxX/J
4Bg3mC/PB6YoSi8MZszyBCvO5eudIycRxoujUOoe2XhI2ye2XDlp5a6wjEnz
g+LejqFMsq1QvjUmMh3mksS7szC0zvViyuWmUMl0hZGrn9biedA4zZsHnhhg
JC48O/IpEBj+Czdsnsl2mA+uA1sbBq7dut1XchFCQaOJlLlwesp5QoBuUNIQ
/3NyfIwdJ3/kqIkr3fnAEcOCYFFsMspWLqKGC5tCRawjZdzE4Yh0uN4vagKb
uoggXiAofQGF4vKP71wwh0mZfzlFMa9cgUmH5IzwEW58AqqShVidQnvSkHwc
6TG4nCM1QfGDwOv/gqg33WeM3w4R+kGyLqP2Q0vm4xF4ozm8YYLrldyJcdlY
BtTIXTtnSgp0AfFHdjin+gP1bA4UJxsXx5mrEY1pDp5dFb7UOZ9lB5ZFYTyH
NOcdheTLVqs5my9dpmWcWeOW/tWCutNGrYPm5hNjLDQd5a8IB+PNXv1Ya6JY
JqA8pevN2YitRWIbzogJTmE+9RJ9xz0zB9W3D3YpgBcNkkZKfXxKbKRUl7G3
EeJVzRU8oQUV2PpPXL3be76CajxgZwUjMjs8R89CHYiIp+InKdRkBZnwI1uS
TiV3NsMMe4zcqvIe0e/5djviRLzmqpQnwKBDteaYyHshfjo2XprujzYJhZyW
PLjska/Oc1HUx5Lw4+NINfDKs3PzuhmlGroxmH3Wx8xHDwbvxtAi1Mzn427X
7NaYI+LIoWm7RhQsFx+73eNgMLlJEDWpszyoxsfXTT/fkXcq6fnxJLBxyI4c
c0iaIS9kL5hhkjEyzrryQyj0mVzX+Yyn84fLiCCXxpoG9qFKHYz7iATBOtU7
WqUoG3N8K/l1T2BpvQZscaVU32oYltk/IF48ajIgBSFfHwVNIoYc5KJFPbu+
eZEgavbL/oGGR1jkpb1Uw3aaKFI4Wry8NLW+lKrMoPEtJSkqZ+BoKsWFb7Lu
qf7+7nfzK5qXsY+bJM96x7IO/zAZyzzv1UZYPl6LyFXUR04USp+P555uAjkq
ySFq7tRmj6NtirjYRdqRFxUyV9+DXfN6GCULlBGnHq6DCBU+qF9HSGeeaYzz
Qp1c/NIxiJl6FAGqhYVcRKAIw0NjzmsXx7pUq0oWVKHQmvp30KadToDIzrDT
Ipvrt3kCoO/LOEhlasMg2Uxv4d4uf2ApAgpUTLliKzrprB1plmyirUM7Lhez
jRMnCwYDC3DsmDaQZbefAsDyFen4MZ8AleYZRw0LHNB0Kx9kyb1Ua1JzFFrN
7KqX4MME3gODakZX9LXy5ucKFc5WUuCnBHXPbxWTtolgq+KWZDPSJX8gS9FT
ZeaRhM53wmFSWCS5QOYSWPLF32EKgGPeXmvd8EZN1272JhMPDBucdEMump+o
4eTI0E5M79YaFH9I7ZRDnD+U8rJXUq0TYyL4yXvEmRp9s8VOt2+mRWLXtECe
APushh0GPCxE/SN1qQm6In/aTcnC+nPsR7aT6bPtz0TlhSAkhRLIYgAK1C3L
tabuvWycmsJhOU8h70OgKI32RfMC5nsDB0W9nBGHHMyL8mXD5ZqxzypyH/hL
4bb0L/sbPenuFhsveXdHM+SpkSDX0tO+xCZPXJIwC1X6F8MWdhZh8ab4H43q
6Y7pdl3225xXOSH3xGAI73Xj1RxyOJV70tkLntQpJbrduRI52T7pAYnsApoc
LXTrA+5NPNjQnysObHATWFVYBNpThBa2PfxCwE6uuNmyu2PlGaDVq/Zw0Gcj
+0lrqD9D6TglRrWiYhsWQAaP030aJXhQ2fwQ3oU5B4kNMjYG8WkndWWediRL
BgkdFxctCdjSMQzTpcOMnqf+37teLpeHWd0+jN7mQTLaTq6k344rtS6QU2Qr
GZrVWskJVungPEwy4/6/668ussPR6S35CpxuHZd1jElZ3B0V6AS8ebCIJxSd
UwCosCfkIfQEmzrNDFu1WyYbB9LF5cu5nUGFkg7g3brSDh9jRXF3B0Ix8sM4
oXUFiqk0qCSejs2Kn7yYHVMk7xf8W0eXNgccQA4xWVdHuGxhrdJtp5GLBalV
pB38ZxO5bhXbmdGCay+s5VcpW5kOl2XxgiyrFc8tKZ6GR9/3eaKayJH5J5br
9m/OYF1OqkXbK23RNDIkNt/HCS4KF+1ip1h1DX5GdSAuD3dmFmU6xHIt/TLH
sXWQYSRNhZMUS/2oUY0GALebzdGqch7lOdRgVX3yDxQ+/8XSKJknDZMRHnuz
tcEiL6F/k5FYqx+ua2Fyz+QyqcZHtxD3lHQn6r/6pHWBLKo9Sd4iCbLFL3iE
WQKKgxQaThY6ZLUyKPaH1OUkaZNzq9DI+EfOuxu3XZdc++YmTbrUb4X/bmt9
dD+/5rvE5E5BYtAqjxjLEWGJKZYHJK/qgH5575QAdivt1U9ZY5lmiVLggtac
B7w9vpXGHeiqvVEx1ZZdBFlHeBiNheEqwu/+BKj7XdfwQ/qQNZOFrOSXN9oE
exrOH/xQj708U5r6cWVRER85q5j7xuY/UfS2nNfsIL6qMqoA521bdYBTj2Zc
a/rcl/drpyfIL84sp3h8uHtxJnqgKEtbNMBdIwxdmrSlvL5NFsaJyOk8d3UQ
OcuUDqFb1sw7RoVWHQ4JTcWiwV/U4Pg99COnjIalYp9DiMRFTBA/KLW6g/lg
HcaMhmn90rQjMgH40jmTfTQswcT/emZbynRqEwt5DIMCHhV5nqe8GBdO2IHI
1jHm1njNPWLoSMYj9u3d0II3T/lg5OEms9Kg5lGO2X3szgjjLLrig0Yw429w
7WGB2ZgcqTPjBQUuglLhpt7bDq0Pa7VOiXJZWxayniUEg8WafqDaa6GSR+6O
2vvu/8l0kMyHdlpH1tQf6borj8S3PJWtQk3nc3o66N0dXTPr8zOwsVBpzd70
JFUsTeDq2s/5Aby0XBIQTb+xxuKdm9Y8ybynn1TiGL6oKd/d7Fe2ileZ5K5O
gaYw6t/7Ox2vdqAOIanjYaa6EM92bgzQroUP37f6G6qmgXKTyrGiE/kX6Wne
jSHleZJ/dPaUnwIR4SvLo4hRceQsJqnlAmITppE9XGTnwWzSlinsn7zS204G
0mYjJzoFjxdL/Ub7nvC0AyS2wzACG/SHrt/Xd9K1ArgbaRWigHRHDpY8BAaI
+VIpfzgl5c5u9e4sPNgvB1IO6VmBbhw1bJoANOix3KMkKShGGT1XxDXBPhki
sCCGCG2DB0jGqVghgcs/dn7kiC2VU/FDsG8tJqSjno0T7fDXqx+eQyKjgt7t
q/EUJgliEQWiNqRef1+a9xOe7gQRZg0VjktReCCSMey+8LYJfQD/YUJ5g0fi
2CPJz3eLrGM0B6ObBXpeelE6KO1XO1emxPXNcchjP9iJBNp/NBbpeI42mmDS
p1suxA41ul9ee0zIhBXc71K9pEFdYB/rWaL1r1oWv+a/ZR4IROEAT/pUTua9
afHSjvj27khZjfkTyjbur1+hhosXzKiX+/QTvt5yAY/Hh79IkMV1nggCt7b9
Y6erzrFdqsrFRlrLB8WNOHKkZzpBroFGESpXcd11ixDm9ZUhEw6+r497a4+H
R/JDwjbdc+NyBw8risJnyUwiKN4kmTTsh1lyUtBJAnpRLrfwrrD2jIRJe7Vw
4G0z+jfuTnIoj02tySgxJDmxAScFrogjm6DfRF3GylyVgwkMU3ThtCs4v7cr
SeKWkqmAZDnjZJERp01clYn4n0Y7dObq7Yq3HWlPl5IpxQgpKFM3UjYgk6qm
dC5UFyw0Z39FvqpzUhsptDU39fq0qNIYOl9s1CkJTH8uHzvc65M5v1J2jTsL
NfsU8rwSIbqljBvVqzM3ATkVLEaC/COFEHdLw8z91HKGqb4pCFEWVP7jbn+3
T3sTeRQPZz1RS7FygbXfb9bg9LSJm06kGLDVBFPXC8mHVUeGjB0qhz6W0iqf
z2lbUBTGZKDyHaE5AuQ3+/o4dcZKMD6kXW5TT4yd6A5SxtZQP0ZRDJriYCCf
DLkaGnSaqIRJrL/l2MuQ2dUPLA6LgDtm+2D2c3tW/gsdVdC2kK5bm+QFDsf/
vQcVN8ehiq2xIhDi4QNR40NFG70Xcrcglglaf+mA92Sc0LkBAKYZCC49DYTE
305ZK17tqdM6JDYviZmZ+a72+dGbS4FmbyaoV7uwc8mGig4OrICPNXOVMdMd
RemmT1OBcT6vAlwMeYJB9CURXs4rRDvuALfm4BmHJa6yd8qBB317//p6ZiJT
WGujZjAXeLQOXJefUL442RWjLUDRYye9UdWWkp8Z+Jfz0QTy9YDvRuPN0AXw
ZxramsiaJXlxk2FomUEzyqvWCleIyJ2lWdAhqYloxZk2PvAIYEyYOwawzSx2
mDj0dahYI8y5s95+c588UhxodhsHqnZqeecGa4MnGKIYViXYeE+AHrzTra+i
aGLKhKRanjkJGsstRwaFOvJ8hUw+Zti+wQSpSKiVEG5JraOKKB5kMXdT93kx
BgGZFxSAB4Fx/Q1yBWzuHkV/Lq5VIXiFcYwG096McwpDpBLdw9oOLjJUK+Ow
ujPZgRrJ6t/acz9wHGpnkAv4Yj/8uYsnIwXX1yM6Vhf6zHZ7hCauv4XYFTvA
UCat/rO5HVry/PWzLB8aQsHiATdQHRWeH6SFEkoCVyvq8gMhmbOdKN9cEjaB
JEsfO2sB6vTb4Rd94zMBV6LVW1XHqyzLLpRRdRFT1Kn1aPP4N6HakZC0/BQK
UArOyWna4quJHe3fGCAecGn2LAaQ9dglRak0CYwHxzCPpAw3zmdvq630ldqj
nwnror9mX/9D9yucTHrwojuZ7FlKpoNhgbUoweOEwwRxhW8P1dhfphie5VGC
a9UUdIy+GkgucwX8r3FShVLmwRmZyCYCO2XqvbWTbd6GBNe6vR+lZSqvHikZ
1LQCQkYkaKmmzqbSI4doJZLCKO1v2Xi8bwVyIJN5QA5411VPy3guczjbW73f
em6MY2N3E0ooQ7HeChmNOdzYUIRD9z07W19NvBdsumA3R4YXQK91uZpFNqpI
b9UgZltCApOhknCOMIuZzeHmzZ+CmRuiqWrF3DtbLLHsY1gPB9B2eZ6z82t3
wXqClMo/xuspgPsUSxWLCXWn5AJyRkuzRg7CuLmr6cCWUIkmSO6L+Vvq8d4l
q+4mhQmojSexw5v5vwVM+bRH1GbnYHtpLyp3So1KR4Yi/n1qYlQ1FNcAReTV
msI7zEurI13XgesD9o5547npbglGMiGZnFWAtcRFJ4kqfNp3ALmmBpr/AXQj
ZyWhPLohWfjGokxxfXcbzDN7/W0xIxXeieLRwrXzXNmLuqMavaAiwqFZVo40
RuSjsLmf222K9SLqZWAQgw9JzGhC+or3weRCEnRTwOnREnwxOxu0mOlRI5Y6
lOA5sx7p2bbGZDnElVnJ01tc5OsZAMDqWFUYXGlUtGQhf3nOBHvyUC5CgSbw
NvVtKluXg3dCGQh+0r15/QMDoI/YJ6U3TXw5fVLLimeStdSxDCcsOcW0yNyi
tOK3nXUX1oLHMqW14ZuMH7JN2j2jpOMWhRZpQRbkf10xHeL8w3Ir3Drr/d06
9KOSKjaaIl4DgBx5Fv+DYluZhl6yiuRg656evFczJhkk+neznvsqybOsVtO8
/EXhjvs70r6Ct9F3PSA+hUzpkL/VIIYXXJZvZZcTEzamWTvI7esKx14Cmu9I
eXfS4311sAOnrm0if7QOnsv2UEEG3E6d0g6ww8TbDHzd5LrpHG3PRWSpziTO
WEVAx47d4CwSMXo4qieLvHqP30Jpo4dgJG0qh6FLTvb3xwDIsTGfv2eSwgBZ
ylmQyf/a6vcVDNR8Xb9Uvmv/JObKNs+M82N71x9QbjX6Y1lDbPJi9QuL+ngC
5GoGQ+VVoVveIPpArWw7k44lqHhGEMVU+e1S1iFWOyp9mk9qyZDhU8UpRe//
veCwPoSiUdpT8EFhut6jfq6hOU2xHTMM3GWMU3gZ/YWOoV2LQBgMV8StjHBW
s0+oEqq96uHAUjvoSf1ApQYNX1TFMUM5tQD5JQdYqaKdR9LWjpEffqBumk5d
hLUhpasyby9XQCslsG1aWbZaTZmWBY9KisKy8Ie3ovyUcfUjPt0EW0WXiPYC
yut+9ceWuIYpML4ECyLJelNSZ+MLaXWlDtp23ywtLNzT5MMRqWbgKIA7lbDk
/GLTnmg5oni9SE/cwHqQVeI57ZwDvpQx0A0hYZVKqhp0EyYp3RL4s5BQ9HWT
WSdUXBOFasV8AJHxq7J0lSXtmZfc8oNdKMJ95M//l7l9yETp6y6TdwkxdBPH
u9+qRZbO+oo13owwQw5aHsdSms3WwtmyfNcP6mAKwea7qeFnRhOOp4y6qdSv
2oRSn0sF123VXvtcjc7b5UsHtvngXQWyydI88qypN3b0wda6D5aRcEvQ1nEE
y5wz0XxYq3XqLsffu3ey8aaLOAb0XVqgMQKGFVJhcO6ceN3OdMAXyg0aL/VO
jzTvH9HVPkCIoXemIs5t3qvzlNyiQh5yzBOUFyF6xeBsytQf0ad7q/aO6dm6
AAssug8q9xwysl84dk8A58NioryxtPL6qWXqlVaXnh2d3SvXqNQQUO10Csot
ZRTL57VeORAe3ikVPZ1jGmRyC7e2yPY/SpV6+O/cL1rljPE9i2r8o4ZMW8ON
jVxZGPvKIph2CgP9Ik4xhgV49TxMvBnPKfIm2WYmMfZp24Pj3N1aiyRboYJY
WDVc1bFdr6bdYXJEO4hgeThI/JIiwvanU830h4aFJkfOiXxT1v4rq45hgeW0
3yfxaBJvGWqF+h4qZAzsVWrFccoAhrVQz7dE8k/pCWPWwKv6aH5audWpRuRL
dRXq1ZO4E2PTDvFFRlN3pPb3wzi63arCvtQfM9mANF78PqTZdUQEkbDVMENf
nR07QSVq3Pvs3eip9gln+cEWdxoeygSZV10ea2GyfkkDmZOPP7kLeOSccg9n
CwRyZn45yYKzGO4Et/kiBXbFivz57ArfDyEENqLz2QsXuUDGGKc+TSRHvBRM
7CjslUXxLc5X/cSgaB1WiuA2l38qad1iYHrVfHkKr+VbzI4JIeRuR+GJLaLr
OKeGhVg7I15bScn9HHNImX/YbNlxVdNTykcHZy5MxGASrTuOCCH28CHKrIYn
76WaqYTnj0YPkhvkUXY3XyCZGG9dCZrQyT//UGJacTK0e/ItpDtndyItprUY
aa6/5VjHelhx54qQkIV+ocE7HVWjJYnizwW2ThXPiYsQutsKoOgMVzOJPOO3
xktFnIkwDa7r7d6G+rMCGqo301zF5e8UsQ5RuTSWWyWC+9KDsyfeVnea8Gcw
BEXbQz2FY1hIly0LGeRebLBJRunqEhqh1v8c27eZ3JqE6liF4Zlodv/AAB50
Fe6dHmV0P1qrBiXcHw2oCxzZxcUkYlpfZyRILVfuR9rt06Tqr98UFmq/muZV
bsw/Km8XOpvF+mnuYP3vK8C6djBDyonlUpEGIC6zMAuZR6IpyzskYaiJ4sWl
Nv9H55gj0Hm7ehK8DTVmRyxLl504HUxVVcoJEI3huIMMGSb4hfBEDCFKYkux
RiHTLW8E1PPlogPUVNT3Wyuti+5t2jNRHtxDtOFPGahypnngvN/k/NYs9R7k
BB+iPPZRsANcms8SfAYVnD/owjOTaRY3WnYnlsGQ4scBXlVftdpMvvgz3Jxr
E+Zj7PSVt3zhBbujIVt8p1u7FjHvf0AWFlz8uneuALpm0XOYqPpiL7Zx8zt0
G7pnfYHlsbP1zI7Au2sppJtgqaV/LUqBlpNYyOwQ3/CD2jbmClDgP6Fn7zKs
MmJt+LFb1u5kX/DQFBNZuweE8Gjvnt5WcFefVmm+3llQ8QGRl20ywqBCF1FS
yq9EHrFeZtg26Db9aVU1L+zkJSh2szop2MW/uJGHKlhwF4jBBT4ZZ3GdcRBA
gg0Lro3MmtLgV4BNHsHUXGC5V7BD7doalMI/tBgnuRSolzxIMjOUDgbBRRdF
M16IAgcVSTd0n0zpwPxjlmvZtVnxYhStjV+W3DFHNka2FCb6Zea/DFYhaXrP
CAM5WWUU5z7oTeso+VpCQv4UJry5Hxd4YGv9vPdBQki0nP246O88dsoyVvA6
kUAq+Ewte42Md6TlplhlFRqfo+mRPIgUIrKvqTlVxDgfshErpnmFnz8nmb2J
cy+YKIhsPFgTU8esFhs+1F6m2d+SUj6gHbWX98iBF4PV+0axPN3HJlv0TNSl
pX4pIzQM4JKztOO88lmsEaiij6gORjy7PCTcde7BX5Z57u4ZsoUgRQajhpl9
L/cUgUYqio1L0AYRkM596rZZPMJiDlX2RQ3QHpqPjVBAHD+zfuY9IVPNN9w1
+fENqXHPCH/FnT1gvFEdOxdqJ26Ul5TNgKtLGLpKvd7bCrV+5BM+6DGeP4LU
wlCS/ODUWUqzlUQS98ClxMjLsln3PitYQ7R0EmdPXKbwZmkKHcXSYXXVNiFh
NrggEdxrzcFobh/3abQ26zw/pXpCmNg4UD0pSkh9ieL5xdJOFe0OJZKsnEI/
9EwPHqWm+RMe8wPRGjx7PCi0EBp501duHCvBYkTT10Op+b7veo3abak5gWqb
ObABJGZatnzXTHSEEsvj0FkQ0umq0NHwZI5Ip5q/qYYt+7ondqKluhIK7zm7
+N4o+mILNFsQaS4uRZ1bVij538TG0W7r2gjg347SaEVRyT84XxFW13GB/cPe
Ej25fe+0FpjAhsJv46F9E1ay8Qz6I+9bZOJZ9XEWtA8otfigLTzARUQWTdhT
7jXuviNtsC6jdAg7UVMux5SQmweRB3GvhtGXUpQjPA8z1IxK8HmzPOXsKque
e8kv52NGjI38I3TS1n9KUALtU0PCPorqgKKfR63H0PZ6XPVCVkiINrnBwUAE
sTK1CLFom1yPpk6Q4IbIxpQlU8aP617U3MtcSROrit4Dx2vxnAIAk0SikSvb
qVGfbzAXeS2FbcXpuWPAGGoluA2Y+C7ILQiozT1kiXhZ9NlguhZuCvMHt2/V
Ij8CuSRcQTtd3BNbwUIFKlAOZBBtlyCdwYEcrRdzwFn39ApBqqfk0h3HYnDF
r7KnvLwf7b0HWFRIEljPCQaGCV83d2ULLZGeXpYRpOJ4NPq7yRB1/JO2eeFA
OPdE87pSVzGoePGG461kn/5wClmn0pIZs/JOU6nBftZ4bB9n3Q1a4Br419KD
SntQ6W8OulZbAxiPKlWubzvBMMWcIjb+hmR7+IhoFODo9Av8gsVoBNUSVAsD
qx/2ajKsl+J8FqJJ53RLjJfs3bL8WLo7i95jC929pEjBfZ22NbXQxcHYoqiU
7hIlf4me62EKbJzlKWrtpCDbejG9xnBhdGETOi3T1xIES2bSPbLQv4PO6ZsY
jEoqU57rQ8RSa9mcJMQwskQroIrZ4bB0Je9Y4DFqaQIaSPVe82NcO3+ro+VY
Xpg5A6i5Vd4fXq/d/Qic2Aojk8UZ7Uq7527VPryztVT/l+4kFYsI6XYsI6pI
Hi+3dA+j56LzDYeDmpcGE/EGqrYDbJIblhuqpjiKn3n7yI2nap6lmrdf29vM
l8sOhsCYAW8cml0+BNcKzoTCH4Vj8e2FL5e6kiMMgWPkVMrbgINDLqLlpYnF
9K01E5ufbETbPHVP6LZYQMjx2XemYchLKMmRJLJ15OAc22ysFHl+wNTPlql1
Xra7Y9QwxBJzd/Ey8hMj+bX/KRCVWK6NqLAnyOcMsRmZQvsZ6+MQSfJDZnUm
yJ6yT1GmpfFiRNPKbEqaEuAiiI7Du6SDgks1JpcQZDySn3aCMAQ3f9C3Lpnr
jzP+Mkr8i3QjBBExm4fgM9bYfTbo2F7TQaQ7y3VhAAPssG3QgNQYWJQPCLau
csA2FXxYHz4F+tt9nozpJgrqC8WZOvVV03eW3AOM5m87H8vkw8p6N1v5i5yD
aOpy6VTtWyO/jpH+qVe7P9kA1ICX2I1TbKp9lVx+YcJII5L+PR1PGuAqKt1C
1Uq2Likw9teW4nVjTHAlW2m4Q8mStWyuZ/nvC5xrfWu6+iQFqHW5JS9+dZ18
kfRpsDPTNMUIWgSZUcPJ1HZsE3SRmjesi9sD4Lq10J/a0pWkbUuXJ5FxkYvz
CSLKJ/DB/siF4RyHZeVF5CNc3qnNVchCt8QBnzGR0skCcvb6x3dDPBs3tqM/
sk4AxjXbWCsTdLw9xjMuKftSFlq6MuqCDuD+HeDwsNL/jTVCTFHhRT+JM/gX
8bOs7xAVOWFfajWr0cbyhrgybwVMFGCIeoFJ2CsSX87HIvpRNvEe/m6iZw6Y
7osvUAtP153lQBF3NOx9Fj+07VqYYhFz9ACZ7fXKkYRGSC5vM9K0MSbq29vt
yyee0vVhS1UiovqJ+wQDzMF8uZD1qk8ywVcTaknprFvUOgUvL/O2dWiqFwov
eiO8gF4Ipv3/xEu1u2EnIirOLXHy/6mZ6GEo7mCeJv8wC+EdXkgvpTAhu1Hx
pJjAjqUkzgGu+06SYketrhF4fhBMI0/52enblTlg9linMApC8tep8QvUX37I
X1iqS2j/baQtVj3OS94wpYXuTYo7OBf6BtKbM2R37JgungGotUOgy1Xbs1jD
keZ/wn0owKzEBZaaMVKK6cf8yh2nq6F+W+bWde9YhyjMG+UnGFAl1pvf6D2k
XN7gsIw7RCZaPuGLBgRC7iSV4B8pMbTESVJX19fKp3eg1TBzZygEyAIa1FBn
qRd95IdUVsppt7FYfnblQrHuMX/4sUrYnNaHgLB5SDS4ZleK8l3cWz3oi9jS
PkyfAW3LM5rq2Lz5z+qwa2I2BGRmZM1AJ+/ZfJwCHafEG1rZU+28YjuzyMEH
QMoZ9V61ACWZc05VmU7ozeeUSxHUncwsTlqcyEp7jVHOg+cr9h5chR3FbTi5
weVieFvllKFqorQ3Clc2/wCLPeTURy0rpw+sJBBRiByxzoNzDZS1tOd/D31/
tLqs84H02PCcgMfUFi3tnHjA6UcIFv1CEZFE5hwLCLW5x4xUOzCXKPHlaB8j
VetKl8Z188uIYw+ehub/PX5sNotdesuu0+Amuq2ofYhewvb4bf0Tib0qfVfQ
m4/kf4ebMfgX5wZhnXylkzht7Hr+pRzzGE/2aDj4nKzE6s1xRTqrIWTOh+aB
2DOwVsQQ5w5Z2qqQwd5uA88iYKMYD/NWsP12ygNafTKjwJoBeaNKqkwgbyim
J3EMOasPrFHBW+Ar75BSEJ8VKKR6R/BRAaGV5GMej/7fp/cxDPSVdmtBn3jl
CkqULdTjPOmQW/4ELggeg2zHgocwE/qbMiotOPVmHyIfkaSC0Pt8PFNd5PjD
KepwGLfwyya6mkxHgIjcTbRNCGzGUGOFJRDM5Fjwie+vgrL/vv6o4IKgU57y
r+VjTMg5AviOYDAZ2ikn/qehgXpHIo5Q60pkFUJCMiwwxGFmiLN0zj4R1cl+
GBICJBVl8eiLTbZ5P6NJIm+9qM2miK55cxwkX/grN9xoLw5Kp2p/s7p4/XVY
dCDFjukGZSQU5hfn9PRMTSsLC7WD5KInBNx5pM1jZMR0NObPakBim6g3Rsll
9SDMr6GQdU6b798KmNljMFdyh42YpFUq0W7WY4HbUeSTFE/OBm+5QzFotqKT
9Dj1ru6ixZz1X0hMibIblHnHfyCel6NMai6mnfCyviMKL8gaWuLnaLxIMT7T
/K1DB+w0JFY42YCZYRdVE4MQTiltuosAmca6OPSDsa8qtl9T8b/M7aLc+WjA
c9NeTPNlhicdhARfD4L9Gz/aEObpdIRCT1rgEnbWWUkEGeXBF8MOxYKqy1xz
bMpW01UzT6Z9ybr81crUKelM+bXe1zy9vnhCHMrml6x74BGlnniQF1V3jbVz
0iTLCf/dZ4fAOeRMxaNC7N06ElbtBIITBZJbIPy4MX53N1r3zXrqb3CSUNXT
PWLNoZ3ViWCSDCDSi20IhVH1HAWxkY7W434HLdV62Tu4wnbL64GHWVDjuaNH
rfZQCXF9h7zsHeLgy/+uW1PQeSKprIYWQXdgCUYk6LRvUu1ZeQNZCJt8SKRZ
RB8lLm9bFdwynLpxWK39qK1J0J7aeyru6OA5nB3t38AkoF8nBNy/5C1XrVJy
CvUb01e7cakVSWiO+EkeNmM7IaVYDSwMpDQCQOmnk1x/sGwgKY34Id3Ofmoh
I+9AH+Xxtb/SZa7C7C40/3TBL3W3Kl91taky9XOhLSwYSnT+yDO6bDJhiYNV
Ky4Uy4KL1EJfW731fWKrFhH/Hoq9Sd6oqa63WAIX0axZ1X6ARCs9c/yRABX+
/B0Aifo5fRqDq12Q1Q0ida/0Wvp0XBFjJV7E6vIbyyxTZxCJNqvKjE0rmEDd
8Aecw+AcoQbABb4rTRJDYiSZS8+ojdoQDg9uM3NBNHWCZA/iEg7SrcrNqLIQ
3IfR+ozYLMEvF7DLxm5emQN8kueZjg0AIUrIPylm1SsJ3UhJgHM1y5YoSb6+
NIoZ8LXcXho9EeRP5inEbz3TQuh4h9/w48kZ/TuFsWEl+GJ1Rqs0wXOnyX6v
lHFzjHx29KPFp+HprRm66dV7oYklIE4OasmfQ3M7ySeZs+B6pup0/T8mtfAY
CFSwbybYLaVBiNDXDAvacYs92c2FVzC/QWQCTzwlu2uDWopz8suDydaucOCt
T9BIGxnIEyrEXWe2Jmn0q1BRS0006B29aRt1BqfmgWIL0XMtQa5Dc1QT/VUK
k29PQLce4l7K2Hxg0xYOwLSNBMwvz3zN9TWErGf6BDXqKfokKmk6ia7jsrx1
ikSGn6ZZkVEnKAgKk3Iiy5CXAWhoEiOnUc1VAmcpI33Cummvnp0y8re0DQtP
Txy+B3W9gsLbpTy6rkmmwi/b9WCKh0/JQLpCNTvEYAWz9RJv5Lz6GVNr0v9j
uWh/MNBPZWbKLyjRGdzGWnCd+WFeD8d4p5UF2CoPlnMRyQdZwTo+qYlBbfNO
X2N4Ih9f4zj3eKRJwLCi9njZ0hEklnuQFaHKHR6IJiiWagke2kO9RAki7I7v
o+uta/3m0UocTFKjs3GMWvQl+KPS7spWTd63ATySIT2hhmBJrKZaKF8aN08p
cXBhDnI3RDs3R6TevMmOIiyl8HLMsBmb5BQtqf8C5CHiUfonAtllrXYfmv98
hTAzUPInmL1p6Tt+KYwYjLwnShYY75SnkyrHOfDxapxm3qaHmd5IHcb4En6k
EsieEXyGQgJ/gy1orQmAUmd4LWUWsdMzke0I+NJifnVM1r5BtCfHBwRhDOBZ
98IQHp/lmaJOkoiTPaU7aHBZ/TARaQa+XRUp/EBvXaSLaw+yW1uxA0E+WaoP
zY5VGTW8OHX+RHy0fBjrLHyJvgSHPYBUKzW6x9do18RLaLW8n4Dxu48uMaRy
sMM1XW7xkyFiSQAD3uW+yk3fhn+rgr4TKYBshcPMGeWkBuI09qY0EDBTSgCH
53I7pyd1IJP7vyp2e3QnnamUZl0AHxTzjehsjRKCGDqskFIi2tCOCjWxNZYw
/vafj+df7jSc5akOqwW6ssnyUPR1Ae3CwA0nNGuEOb475knkw+7qjfUG4NVU
V/MAqsKYXKhqG5T0Jh3H30B92TTucHTKg/2C13ABbKUMSkvD5zoadcivVqDz
es63mFCQpvgsJWfqQ2jqa5zcMLjFjmjwqR1/Tmh/XX4KGlOBJA+PKcqJf+kE
Qxor6oerbK02/Mcq/euZKXp3L40LEnrNcXVQO74q8+r/cYL7mjLwzwPXZc//
dPL4ZZjA22x25iKJ/NpA6oRECjTFFQ2wt9MfbMvfbN/N0hdz9bfQEe+X6YRr
xAsy7qYiiybaB2Rj7XVDTqFVhKZjkZ7hWz0gacNP3j91qBkKGP73ehfOw8Ak
Eh3lEFpS2F0CJ8rDHJo2XOfJEZSe4JYuoDlT9YH8yFh6o6XqQ4XO+MUTCv3K
7oNGEMjgst9X5EAaVfznOJcX3O/iZiw1G3QkQkg/rAOjS3LU5boLovXom+i9
OQHK4ZA8tj4ucMsed8EP1hiXVBLhklEe2aGP7pm8vLM+UYkQKcfOEK1N9pL+
sLVNhzOl7LGLTg+3NWnl1I2K0BANdzh4yZKIf4bb230WRLYMsv1ZKIHXucLb
Tt14/xAVstOBF78gnp5SQhtAvcRtjlUwDUBYslXgFWIkcHFDvtlekja4BAJL
GyXHD/o2e6tytryu0w+yLimHnrz0QoEmwc6cDASnhzTX41F7pc0OGVFv11jT
s4f9feVfGBFaPYqcpINTtgBDIvxBGiy6eoDmG9hyqh7cXNPTa0Ek0qZNitAt
+MwzAGa8BVMnvj+hcVchHb2XRZgNL0uZN0MR1RS8ozm3nDM3DGo9HC+MiQ/T
xg9CInwdGx2VI9I719r9bYhq2FWvQhQtT82SYsP4fJFuFhrwJbjMUJ4pfcv0
CBBdQdw8OrpoDYpvIbCSDryhwFLztVzJIZP4VZ7cDRQs7GIR8Ng/A4SWckhg
yLs8kpePg+8Qx2eCOuTUFUTIz+FDbGxBzgpTiZD76aabvVNGlRcY2rAeMOtw
dVNpa7zGlfLKmGVZFi1w49sbZ1FLKrJjRi4MwF5ogRigg6sWrztZ2Xl5V1uu
GxCDhUXYLArwH2cFfH/JEOQTtmldQbtYRiaWR1vORaYvKRbL9dr3OHbDF1Jl
6OOqli6K30w+dFy2NqUJFATAqmbmdIGGy0Pp/3TYeVWdzq4HhYN7pNuQ7kfb
gHWWTQcqy5vqMXdxGhQXys6GeqTlTAObPZGq9Axd/nWGTlEG0o71VX7VWnhf
x6ndTWsPm6YT43PgBa6B3vNWgN+sq4/yCdIC2MajM6FhnEt1YazpICNJWTh/
UPA+g7NrUfd5L1fmhBE/mZ3bthrC/TIeWqCTC4TuEASuiNrVbpV3hP/hCktQ
SFXAdLjqg5laRWOZurxIIo0gFyWrGjIp9ksMFNXJOHNKqxADVTxU/lcv+xl3
x/gFHKuptBcGn2kZI1xd1eT+nzlxpqIs66aPB2OpXZ2z44k3HG0fNtgDK/Lu
2k0L5ibpixUI0kro+pL2DLymGMZiPxe5ktTjLpOM8XZZVuPvx/VEOTt0T0g/
AN8ae9lM55dUpvuaNtDrpda+K5X+fCAsbRXXNr7lFOf5UV9bB4Gz4KVSmINn
/YPJOouLS+TpO2Mvw3CKJ0qVRuNLjMnjcA7S1D17CFljv5ydCaT4eMOVbeJS
46gjd0XMyjSQxnUXZjD8C6BzJQRyM564YqRxatEPE2B2KjefrVnJCOq6MDI7
vmtypscPufmUwbtchpPn00cd+oKBB5N7Z/IuP/Q9oZOTDwmHO5LMiE80WCVg
EDpQ9R5SHsWrRq3gYBK531cvS5byBlC97s4Cge+CtfOoglLimZo2S5TgKkK0
H8vg5BrkDweiTz517U+ToGPFkQ+Obyvz0yLa3u9NEwnk7M8H9mi53h6ag5S9
g5FsgpkHuw0uaFuiu8rjiyIhIawV0TxGVm/5SyB0lwJh/J36TALqZ0PV4vt/
sTOUaMkSjGqQO9t5satKAZycslh/39WftodfMOg0JNKGngOvu2xAwFCJdd3x
mDhMoESvlrrrC4qzqLO2bB+HFHOSCDIrKwS5CPhNE0pvbMLPp9MCwN/4DhP9
ZAc6nnAAnfBJhIbNs4e4rKMhLn2DEORhm0/8q3nZq37SMtCy6PR9Ub2i+e+n
Nx29Ocke0dz/6GZkaiwaNHTp9QqUTu+ltpd0AvO/9CGVia1HUQbi/aPh8oHy
5cCj6os+Yhtaecp1DxbykaL9NEVdRbCf5xT/JfanedkmuYuHhAvAzCxzWoU8
IGUhDWttIi0jMQJz3YKX+V/ttv6sHkPCaUziPfNv9AMUgvKauzh0IMqzJd4g
0p5mo2J6xcw97velpiQ814B72YxY3R3N/0kkmG98K7SuPCmZF28DMh9AHwoe
uBAGZ0BMn115nsuDiS80lgGj0iZGJbOn6R5siPugb2EtKl+ILusCojC07LfV
0yC4SJkSojTP+5qkSZgwSwyclxgC6SL5ZvnAtujKHbpQ6ELoVSCw+24SO63M
oKAldv+cxxZBY7di0z99ipWQKMxqbVzut8mTDyOB1tSySqX7x/AfBtCfi6qY
OcpHW/Hw5EOdWdxUWhRWlastgqC7KTByqRZ9RzqsOYig3RttjcLSaAk+lhzW
IRSWzRB19kWuMliP+voEPgpbDuv01FXjddHn3P5aeeW0svbraFc1+8amu6if
n2WnZmcFxSMFOQ7wIII2Pu/9456oOSJQXgzkr4tCrHcewZuZWNeOapvlJYJl
1UKAi5+PiB6NBTW+dbc38W7a1gaNXHZeHoZQ2HdQVJl04Ej15a5e3BAjCt5X
WD0PJa/6shtItngmO4pnVrv9YAcrTiCsUaBMBfIqPD/6KJjpRaHz2bNyN7GO
fSNAHp0PHXCaicUAEY9eQOULceQptKb3gjJoPr5Fd2PGKEvx1IaztbJy2B+h
epprmiJvnv7GYATkd1VnSh912NrXxaoeXErZzSZNJo37n4yUeG6GXiaRyCU+
QDDWjqCFIA412nf89lNsykrttnUvlJBMS/prVvu6kfTA3q/IlQVdYtuNL3Ft
oOFizCUgVESRUjN0CVwwriNDZAs0ooxELs2PKhIyklzLgLtZ5bd6OgCjXtrW
ChN6onZbTNzsOaP1UVynJlrBBRIktkq+2Q5CztMXV1knghyAfWAuLXJx2w/V
IkdVuK09xSNWuK6UZgNkBWbeThkcvUo09FI861RnVNU2/5aq3QUIn9tbzvdM
jeDJpbr6g/wFSMHzWEhJEvCpY0eM6WJoPhVjUYLk68cF8mfaItV6x5i64h1H
GuLCyjCDejgrUV6kyKArGBuha5oWha8z8Uc8bR5FbjtsNu0s0vy48i1f+h2A
8N3vtRu+q/Yn7cL/56QVXsBVm7G9vwKjmvI9zv3xYmvDqDbtKUahlmmKgcFN
PHGfAw8G63gZb2hhZiOpnr23C7zz7rWRWp9OkC8Sg0Txh2pHczsgv812r4NG
eRqcddwZq/uxoTTxR7I5oE0GE9C8z5QtcQbDQ2vGLcZchhE0az3mcE8glrGp
yhgKm993BD2cRF9XeQyXdqC9jTuoNpeeF0GwQD7PXa7rt+7YK9h1ifGQQJaa
+7yf/bgNnPDfcLq2oFwj3/QbMXiTMS3/bPQB0FEQInyjIe3yCmL5VxoaKGWU
zfzrE9F+of1eb1sI8Rx+7v9j03+zW6K0G9DQ/MBXqJvlM0UzQjKJQl1ceTZs
e39eK8agRXWr26ON5qqCb6SipS1X6H3qW+FEwbv3Ww55rBAG+7kBMBbs3FyA
PEr0vKvRPVD4Ww1zOA8th51vym05WSx1+jwzMMVqXlty7OWXSGEWo64/1RPa
98OnV8SA+c8J1UGLQjDpXM6fPAenbEZICXaG/PrDbcvBdj9/nSmllMPOp2aO
wDlazzCLVLA8h9S+5sovm90TLwjj+kHv5HKbo3gDxnIFmiBZ908t2R/pAJQl
tTabn65lUDe0F8G32yHk/iN4K9I5xjlPpXVw0GiqsbJ+8WU0hykmeKwIE5Fw
kqz7KoA2z1DCZnIvayx7X96xAjRjsTOTDio0Imz2qcbldzokgfmNP3dDvbY0
o9g0+0cnZaDgtAu6+sRiQrSPKyIhMRS4WtkyOf2Y8juqQ7ot2nk0vZ6atn8T
iFFfrcKj1CPx4zPFrz57TGpm+wdFG1s9prrn5xtBvzGDc8fPfRrf4tjvzIVH
m1eUcLnrtzH3YA5ufR/IvpkXtcRTLZ7Y42KTM4TVquzm++iT60fzzXWDSLRY
nfrSijVW6+dzK7kuOoaeJjJOcR0YTfbmjlVetJS7o+evZah8NWl7HK8ZaFqo
lt5N8vPrgkHxC7bFIiKuS8J+W7Jk0Rxmz8Y9Hbz2Qbxgx9XRUGs26ZqN+geA
WrfDgvxGlvRRkMglJ772U+YR4RmaWyHPeZCEGljTpA0oKBTkD6L9wcUlOeJR
h8+gWsh/AA16AahfDSl0oMiv4GqRk/sxJLyb77NCcLaCDb6cxHK3XDCe0ZXp
wJhTYWwU6U7AkNj1b4TcIslqVFCpFpWxWlJNEGlvXS0m0s36UBAAzzyJXH60
kwo0ghmeh9dPMMTS/pxtq2ZxvHQhh1vIaCVZaZkKluXYyvqQZ6+amNv5X9DE
PG05pm9RLx50Q/Po/WwQuEGXpAP5JmBYqXT24pPfKoE1vlURSY+/PhGrUEXH
NxM/2EmNbUFV9U8BxMexwppIJn1Ugfj+Unog6QGgZi5eGgtG03PlNx9asAg/
/ISleHd5pqEiMiTqmv2/7kuX4rlFJz0lA7PvLDi3+GEOfakbuBrpMxuVPcA0
BVNEP0Ee+nIKuQugWShQD/in5UXgzrTRc2KJu8cd20MHosJ7f2XulOvkE0Wf
01QuP2M1ZwD1iJigAsq2n6YtLLpCza5TwYYTCGd4H20Uucz4QxmNZLT09Bt0
OH+hoP5mErlbkVbm3swHs/eUgVu/U9O+hBjlzyLw/YgdXUCtrHO9vh9xaJow
CRdSF0wP7UjF1a2hXcHdBza31RbdnTdHzoP6J09T65bfaVVypdJf9h522b0B
5KA6gPbmOVCZnwMZ48huWdNi8OL6k2TvlciJ41TqFCXijN0TKTToAdf3SdY9
Ck9WQ+s2VJpfxZLn9D82ICiKjxsUfveErb4EWQdcbGKK9V1ta6XjwK7ABCmm
5acVLGqzAwO+j2+DxhgvvK7QD26kTHjEyBDmfIEhEGXLns6/H6YTG3TRBysO
eVxSpOdqHrjgj2qQc+N6yzWcEIP1YWyWnv+eK82zot37e4aI+TwXcZUmhCGH
KSdZaKCughsmlPCs4Xt296Sntbjc5XBNjafc3QF4coeYbFWFR2v+6SF/CUt5
RrJ+NSxytJYtwXPeFP5GS4+JsltIl1XFbVIX3S+kraam8guG8udOr3p941ut
xlh4vApGCAzW7gDVIXqA0LPQN5PV+IKpMxNCgp5ATm9sqo8+LlZJ7/paCaa5
UHr52R7bo0Zf7l6Ebd6MmYyUiZrGJUIxW7xJa3a5bfBEEYBcurgqZdZcnMcA
MbYPW5nMKfgBVWb4PGwK99dETdAeAIOf6++rExeTS1sQSWWUssiZsK69P84C
PTkPHxyY0GTFPH/KZNgJPh4lROunEgbqzKwAUYY6N0H+XgOGq1D7CGw5rl4H
C93DyxwdTqGyQRU04DFLAdm/9KoJ0JEZ5aGacZ0tnG6wSlnE/PC/Lo9QJ6Gp
kd2FbBCowxz+bB9NBF7EV9T155LtkBltraSTeek385yW9be5U0IOtcaZ3Eb3
9ASokTmoiPyE/g2o6a/okunzaBQ/hMkpWNp23SNisCBGhl6G9I+AKSOhQP8z
rp9XjZnwRz2u64/sPvrNVHlSvOCLaUstzT5F2ibT993NQZq3vyJsEdSzwhC2
evvbMApAF3fFLAueVfVqCeUyZnDaFV+T75MSETjxuJCNSwQhyHhX/YFUlxWx
G/t4EKH5xvaNcMmC8U72xdYvFDd+Dd0UUHzOPZzdteNWQRhPqDkj7FhyAFir
IW448Zhzs1zCfVOPB/U2B/A7wNETtwlMKsI2oRQk9ZfU2hfX9+JCD1wSW//j
CbNvW/23zDKCdyx4Bq42Ns3rhDlJP5Jz73U6Sf88aaVYeIxCTyKlVDkQzpue
We7RnzdlY2FyoSxlETCbVS9ccbicRqwtniw/Gqgw3x1Qq4HJ/mCVWL0IM7Pu
50Xv653fyqi1WAO4Z6dyA+Xozr2hBfdibCdwTe2aJwYI0ZfBAMfkxGbxbzG9
yD6gH+bBda9ioqcUOA0rb0gDJ0t/UNsde97ntOU1VocAhPlJ58Jlb6zydQMt
gBl4RB1a8RGo5ScZLnWCo0emEsj7z49Wg3FBEVU/ShRMswoB/YRhFp4saxzd
ljia85z0xDrakVsnqJQQjRilaerVl9KZds9cEtFoUj+ClGGJ70qJFZrOnORO
Uc7FlXIkcRghc7vKjXArpm45aHKfUdfu5vT7dfZNsZreHHC+2ROM5pZOmo9J
TvyRB0d2UKAIXljjGg8lKbwegog+2toSl85GilblVnIUsScFqTtJD43tTJNg
ZF8W318vRSB+b6ohjL5+qrwiNlcm4C41l3KmTnph2jnIVulNcaNXG9NDlZ9e
wZQUi9gF5tVAIWqS8SDlD1jh5cJL2cGfT1pt0ryvEUWG1w3ae0WlK/piYJcI
cBHTVu0UQj1GhLXsVvkO6MBUYmTwKTI/pfmN1Lux3enZH2CqxAMrXzVz1E0l
cUHUHMx2aQdLtX9huK+Xx/eS75OGUjpFdcvJCx8u9M+OFdK7xwuNUXFpTWKw
5Od/q/TU3IV/FRkVpVwfpY688FqSFGmgyEFrf8PBi3Y5LpJtmni9mCCR7N1v
+vvqezaIk9imY/71PfgknE5RbJkJI19ZFvpO71+fyVvtMtT7AL5VGnhiVn1w
XEjjmomXgB4bMbfpQ2McGX8hKopp0ENIMwUyL96ZdZwS03KsD+u3fx568HWU
N5JKNJe9rPN4xnlcHyYjLYFHmlQHYjmkARDYWZZBp7ZbO9WBUC1Xtyw3fvSd
rnJ0OdAUrHPHc6Bse0m3bnXRZGQPTBO2miQJRZnSceCKpHcwjTuiti188K1G
mrOnz2/fTYDY5ZSrbxt4GxU5NWmlkKDCqBsYYqYmcxaYl+WH3U7LHEeeNLMh
jgeUOGsCkXGZuwraJByjD/pd1I4LNcJy56djG8jddslpL01KGmDbeZ6/CulH
AVs6r0c4tuQf1MTjX+cYrEOKkRbH7Oj95qzvJWcMXmes7aQyqZEZd+P6eXvS
KUrINnf3zeiwkr04r10KShwdHj07fEbFHXEnJFi1+vI8Fgx8NGmYUH5ybBBw
S9VsYbePFsf96GXqOLzhzsm4i5/2vASewl4DzryoOc1pBslxejyR929oWWD8
d7ZZzZLVPnMB/FCRY8TLrsbNhktleTEjkvxKSuTKtNPBHWv3rd30Og2FofyI
BcJOWX1O5ClmNu1ZlgiK6nGxrmcW7/5/Tw2ibIetFLL82jX1VpYHhZHYQRY5
cmXBYuOAoPuo3ptJZcZQaOf4FacA9yOHMC/hHN0WgZ65q2SIDJGjX4Cd4l5x
dLMCgDpd22Y7ttasPMQ65Oy+CT2JzmzCaupNOiaNAcgqDAqC9ixrbYipA5SI
WQFg4Itl37u0i8ZuyUVmyGAmGcDeGGMs3SqNMLZBthyC+zrGTJSNiSD0yDEg
qGK8tyWR1u1Mai5+iZx6BzD8VhqdyJPVyEnYU6eV4eezyN7RFB66Q82I5gGk
7AL1DssGSL4vQnCZcpmfalzlMd8//3xkj+t9UZQ4Y6gb78mWYuhgl9OLAsi5
fDN/gvcmbqXYK/SOPO7VOjjJbd/IZFOcMYGHsqwjNohsFJzVrlDjNnm8YgO6
WX2Eu4xhxlKxuiBzkMw7gi8Hnl1+6d2bd4ZyLGlGCHRdxN763d8l46sUV47J
Ny9K0bZL3iMJHA2HU1cOM3JbISwy8kh9JjzUnyiRREP5i94rpQ8qqP/AUbY4
1XXw0he7XTYvSjXYJJxz3OxWByJyq3aOWgkrk2AWd92rPI70OWP/6Mazj4UJ
tMAsTyaM87Hs4Yr+IYF5PC+fZcKwIaleEpuSY77ASGI4hz+iF/VTWs0YFJf7
eyZaqiLaiF814Fv/uAY1J4MIXlx8yJshQFMRn0XOkCWtiOD2ARcb6QANMFM9
0V7H8quv5nNKL+irfo+tcS6nuKIwTvhFKUVoS23k/d2kTYxtyZY85SgPK7JQ
pvfR7wPPwf9ypNh+Ccz5mbV+ypcbABwub1BeOWnVT9WzrrTmMZggmXhudjIl
mlRy6PDBdP5f0Mc5Ryk/pFCFhkMVL9gvcvuL/a5gy8lXAps6vXML0l+0voEe
zlnhNrwPmAZukxuE2zA2bLLrcOAADo3TN71Jh3Mrs63PrCYJpPNSbNddV+iK
KDcAEzHQCa4tM8GF7Dsdssb6Ocp8ME4sMeCSbsAVL3Xkog9WKLTEfCfr6ebE
gb5r25W/LVqBA/YRCTandgxNsPfs+r/6jtqjQO0Zc6uvtkWJD2pyeY+u3pU9
YSROtwcUmst68c8zK/KDDATzbm/ln4YrTsV+e5GSSoxw3yFElJmOlShoSdoB
gqi991oMI1JG+pcsnTgb5nJCgOcW1rCfgOcy1hJnZe9nnvqErXaLlPt3im1Z
09Amw+OrlXgHa2D3uatFprNI4YGfWBRS5avMRU7v/PJWPk9EoV0NA6vcusVM
RwZXSXgaiy7scKCgThEy6xClIbzkCBKl4YJ9KLAQM/LXwr9CXCLFRJSafCAA
IiV/mTwC6QVfd4aQ9K9UbMVpl0MZqwQFtqL/q+ps455zzHSsgJaQYfElyZOP
yH28Swh8UISGQe9PtuTmFS9aPbzzKfPRmnuWbU2rLKMtYRxBDMpUdEK48iT/
FPk75xRvDg+4r439Y72MgZcTVUpkg7iSZJD3CLm4uifO7m/tLB3773thSSfg
YHXlkJFnmkaKmdbYxw3B+zdZrmTOH9w/sjp/Ue2BZIXjbaL+DzBMtjz0P/RM
mMFWCtN8rPGkD5m6ndHMsn8SI5Is2vEDLgxoJj5LByaQaKKcqLBDk6he/RKp
6J3gE/tpHd4fFcIHoFmYgmHUGUERb8toUR4uiSzU76JL6DnLc9GXjz+2kS8j
rWTepwOclaXFo0FQnbFp9P6c8wt3q0fHb9TrNLlwAOOCNlX3U9yQliOIEj1T
5TLD0fTXDgD5ogfgBKV2bD92cbROXiyHQ00j7ubwkl9+LHMJMZfed+x3dAiX
5ZF7XCBIQBOLWb7x5EhoEuUpVu7qkCXxrAI1mn+JrHNnjQWpmsPU8P4i96Lr
ySP57eFPtN8uZxx42VWcnpSlr/e9FFQk33KXSgUDcto7dAzEW8y0Ye+QpD/7
7PeW8WtUGIpnSP6795fZWnaW59Y/pAMAn1wUkMHbhySD2a+jh39eIhfC+Vb1
1nZ7Ig1eLdzkCdbb87WSzTaY0QrVYR/N3pCKygFTdo2x9tvBFZ9kX1PrF2Lc
hbXcUaNQ+T8p34pOhxCUvf/ZUng6TG+6J7h3sJ09UzezLk95rSFojlzm6ips
JgtqZ/g4TyvMigFvYtk3JLN370oryVMxWiEEIyXzeA6/2EVrmOADxdv0Wfws
kKZyVVzYaONfA6BgavjMb9273jEulw1Az3zODvFYK9dMppCLL+s6tMjR+rlP
2hJXMDysEzK3IsXwfwj199QtZrOnuifQOj5CdXBp0UzMYgyY8D+trm5vlzGD
tV+DRjGSpqI4F44LGjlyLlfZW9MfBfAXaHFAFXtF5S0fYZgroJrwuHRZIcxP
VwyTCBAh0PDt3/jTf0CK02NeWMR10XJNxUtIEUPOT4XLPBT2rDqiXGobR/98
KZ9SQiH3AmabMaib2jKOoNZgsedffcwWELyEZcX7/S5FEz0KTk/npkLvdoR6
zpuS0D8Pd22/hEsEc0OgAW2PGt8fkhJG/pvxesnQRAwEKExjejTG+lrRR7IT
xVPJ8vT39mLBWEoOW6AXYWR160xe1NVNL3chKiVLefDAn/xU7f1HsZwGaf0v
qf9ICsJaHC+8FhTpgTB+f1W2cfXq2KQGWegs08YEncBc+0/AK17Sa4/4sgP7
+uD/5hBh6GrbzOB4H7VUtp3p2jpW5VmbY6TlCyJssTw6rkXw2F8uJXz36z2K
92kso+WxLB2C23/rl7vbbDhs1qNGipvBVn59eD7ANqdeXmg0b98WViFKgnvp
pHa5soGwowxT39pFY37IeF7pWxrsYqab2cTwq0DJiTQ0V5fL6V89ENczWBaW
Ls0g1iZsKX91CDqWzoF+XB8PrEIc2fcox65tz3F1UHuJTnRA/Jzw9udCSJZ7
iLX0x/2FEg20n9dGabDa6CaSxXGa943tpzy+wbNEwh5bpZpPQ7RJXbdMWlmj
ZyfkiM+Z7hQAglyhkHBnIdBMMoFwQOjN+OpTHipuQfXnGE2wh2LX8tIxSTzy
j2IszlL/Sr0RxCFJDHNN0itSmoipHOTVs09xmvguPKvL+5p9KWX3igzbPTD8
lIUePSkgYOGwbnxuTTxOx2NQsw/7+FsN8o/FyNo8fEl6WqhZNmbWF4GULzj9
/C3J4SuANgHDwvZahf4t6jYE+FBX+gx5pgas6jBI2RCMSk/vLzsuTKGu1X0q
IwKYFesh7+4U/V0PH7Gm41sVecBzowFe6FVT6u+R/W44sYYirRmyLtrvrHXT
Xg1lCRgrP1PHG2ubzjt9isGYp2BdhQT19HiDs6d3z9vai2v6VjZGpcaxtQ5e
Ebu5wp1p6bIejctvGoAj7S5T5pPVuIqfNtoiB/PmG+SvH8siNZv8LIlj/0yy
m21k30FiexJFZi7Y0SjcW2wpCtXbrci1vNZPtLunmMH8l+sp+8WUXUzmGiXK
SA1nmFIHSPUMWfBhvzdwj4OgVPCLQOJzXSJ21YdVupwBEcWMo37Zymzv98UP
m9hPwbLuKlWCVsvQyG+OwN97QoRzChDfCd/kNfvh1/bVzx26SSYt/diTyrRq
EtCNTXUJ6AaSnMaT7P3H12I4JajdPhomuDWoIrvzT01dsEuyo9w8SxH+8pcz
w7iZg62sFrYH819aEVYIn/RreXDUEQS6bi8K5LXT1ioLKDEkg/OXhatsPJE8
SWqoUxH+9TB4Bgz81LBcg5ygNNNDXDu8iYQX3OrkaJuo9R0eVnfD+RoBCGdZ
sZ+AI8dkTRtHByXYU0Nsl01L+9iAZx/fg4alj3mOHpLp6giP5FWJT9EbXN36
Xteue38EKYLOMKpMKb7KWr1WUmLKh8WbURvq3BswKjukePbcyP6m9w5N2LpL
Mct36XOMCThdVjpTOj8/fOGxDCOBq9ZTsNvAFkHy/qR2mdo3xd6rUgrQWib9
3L3wlHP0aOjXUUswXnYsZd0wdR+wwLoWHojPqtAQPEnjJQeItPW8hAxfVZgh
MBoHX2c1BAt8rzyxV00a0eWz2BgsBZFnigOV1VHeNJzjg1mqA8GgN1qNyRV/
OkdBOJjNFndWnWv206qAPfkVXrCKGvonUSCSggKiRa7H759AOH/xvPXcndYR
W3dkWQraTHksiLg4UaFgfR8B6FJkTnqHnBDPlsXB59WIy+ovb9xO9i+b81yv
2Oy5SZ1JHovZBlaMIOSyjz4rClvV8T3jImMfZKLFKl6kVNkFEaZvKx5I8ck2
mBy5y1vjOsC/bb+dRHCZUM8XK6ANPS/WNGJAz9dbGM4+rbLaSk48ZJ/wBVEO
+ZTjQGLEB5xQl5mzyZD/Z0xyZvP/2zmlVFt9XIB2l9hqejkA72WjzAzil50b
O6EwVQMqYrCNqPZf1mGoppWfAze3HKRcMrUZ9IkyNPozm9ImUR74yF1sXiTI
hMRimkwerLWqG0E++soLr3SgvkYd7qqxT4s7hsXe6Dpu4tnXssLAPmdI3vgR
aHHBRjeidynptZYzpKZvzBKyVdL25Cz4wn1oC8XA1TOf51OcEUlEjZEgJ/Nq
9vVnr0JAuE6WioXAmWr2kYuYWLRZFmZFPb/Ed45Rml39VSFhZYIcmkkYpm5g
BZZcNmDAavIWgIcZkDaPrVYlWOXprnOw66eMLNDTzSj/b12mQM9QmOdvIw3+
/EMLZGWUBatPvS/dmmXWGBYMEoory2BLoxoTcS/7qHv6yPdJtnUy7rHwblRG
iWQ0AgtbM7YixW/H3ywOF+/ZasxqowB6nM2ur+uqiTL9kT/eyZ3hvqINX/HZ
In6J20ph8dyUWyzhQe0q2kWlYyafoWwGIOs1AmFrFCsbyp62/34wQdCaEXlJ
AJkUnaojKxV5gd9Lsmr48haUpzlrWUZcDvq53NZzKtgKdzlFnt7oj1kfRj/0
1B6/6foV0fzGmOwb6u2b/hAQ8JAzZv5uo3FRkdTSWviwLATfg7/qWkhytHwa
jOKSo8PlQaHSFX6ENDnsXXheue+a/g6EO08u7PQyzC5xJUG178ygs+BaGa1k
MYMwH5pPwhs89gbjgsniWj6RjX8j0VroaAHMqhVQYP9dnqyaA2mxWP81+OOt
nEeWhugeZhRS/7yTI1/a9+J7c8nPnVJ/Mx08hLn9aWNp1gfz2aM3libVs3cu
n0pyA1DiL6MQOJxuaI/pGNNAtD7q5XkiOrl6dBsk9m6WxmXPFs+HTi3VIqP4
PTSJrWeikUMpLGWT9G3DZOORKZR019d0jFp6hlHyc1+8b/eSnSe32dFkt1qJ
lM0fdFUKiNDNOyHOLOE/MTdI4n8SAClx2zY4Qq4/C8OflTWkqgprorD6nbE/
KxCLdp4kA5KddkRtfm9aAjCmDTToPR187DOzEH1CWxQ1+QtGf33ozYpw5Lxx
OFadQbflmIzsMws3jNLq1AuNVUSD3+4YN8uOvjAOegbjEoGD9/2Uox4rBomk
bRcGSJo/StPkZhEB1jK5c+ZAAYwhV9w0EW7U0CN1ZmFsuVsjkSxCVzm9Il47
rvQ+tRtwIreoUfkSGREsTAjpGWUZRMMsjkfyvGyAHv89hgKHqtNe08QPQhG0
nVX+nf8Se31Li9NkhOP/QAAO/PecUbaIz1PDIOGtPhf4yVty2zBZFFWYD86v
yMnIVMTnqUIF0yPET06fwLS4udzjEr4b0bW/UGrnHXHliwZ68m4c1dBamZXy
bXEt94Ly7V7fByPd8PieEfZ23UGtuy4btmYo9HJMANATC9ArgZp4g7UqIYNQ
vV3oq+l29HKiTsS3MuOAMasffwPbtHKztOcWseswAYOqb3zxKUAdFjue/3Yc
MhTyfdyRhNVE45eFWUz7DZVwWpcO6t9JxBpxEegGDMQYzaeibPjb13MhwDN4
wpnU3vdunfsqYWo+edOutoi0NIGTNrnXQxO+ED9vEtNlpsFoHIEWSaXkMjkZ
XCzCNPAGrhvg0RhcoWN7Y8y3DcoylLCeQB61LmyYZ9K779LnKWdCjiTIjb3y
3bQgcdmk9sXBrrkWcBkkiEAuCi6KPc0XLbnxnO2QJOen+t8iQOogp7o19308
7hMoXKUzaZj9eIAxhTG/IoOdGwYMApk4DH1Qnzx0aebchqV88rBZ+qCNvDwl
9OHihfTsBABymq9JaxPjk2UfS2dTzlZrqBQlBvalTsQd4SUdhy3sQLeu6u8l
6tYd0ziVgXqhtJ1Do1+pIbXjPr1sfVsAo3HBzVXGtKARRGP+Dbblg/UMUr31
XTBPNofWDdpX50VHLKRCfIDsN9ElV/UpMJvi/YAqNwH2SeOVDUdpg9TjF5qL
yw4r4JAP7RUR1MUX8M305dg9lpV5oqpeVAOXqSa9myOHCrcW0ecTTG4RffNs
9i+nVrHEN9sACM6kre2ugJOYc7cKWoyxDwyvYHSmR1Q8QWxFwqBZB/tezWOm
JvWS9FPVzwp91XgsoS+dGaU/DCeVSizBVLzYk33M0Z5tJLovAKUNTQRQsWBG
P8oUji1lUDEsVY3nxEAEsWxhFV4Mf4e6Xq+Nqhkm61dV6RzlrpUNBul1Aziq
TlKHbPbibMT9Fp2zNgcWZwggvTZwytc6uMnMSYJuaL6iGpN/kkv33BDIVjiC
6N4eISMygl+qWn+/WoZdJpaCW8sMZqmyrTz/TBDtim65Kjr79pbHxacuT+NA
4GqxBvFPvbpDum7ZNDYd3rZg1aIk5FX7j7DM/6ZykmqFoNYLxbWCYh3Xyc2B
64rPW9Qp1ziYyLgc5wcwWQTeSRMoMebnzayeF4OHloAPmqbNJsJ3PQnfR20k
4R6GPxCFBZfCX0Had17Thsgt2nQpsqxlMI7gF9xwtfE204pjwgaE3xkxfg8T
hDeHtRN7E6TEIAwsXuz/DQzDAl7e4W4FlS6WJB/L1BdceNpcqqqzZJVkfMIC
N/9mmNfa4T6OqXtbHLdgp4JaOnqNO31fxD+Ymjd5q1NeAxI2dlz0Qm3BvRkq
3E4eybfFZirDWvek2BARK3l5F6tPTH+4I/6fup7O1lCRpWP46dMyHQhbLfjW
Pbu696MizuTPMnAeU5euA2yZwQUR3mfIyaDcMAfG9Q4WFBMRzGttHks+jHXG
nZp4fRdLLz31kFie4ZQqxZjvzb9dN9CqQoWmO0+ahgWv8L06TYWwd9fqjkre
J2fJi7mH8miBA9zf8aQVfWZ8bioQ0ituKZCiIIdjIn8maGTyi+c1jz1BFOtT
pGbxiCZ7SMPtcKgPVpPISuaoxclfK64Qew2YjnlNc5+3DHUdiFptKHMTS+z1
BlXk6p16RpVzK2ua5sDnC+47aEd17Xh5+KF1boyvmHes7MzK73kR36OvR0Qm
VQMVCxMEo2daI386Z/oWXpj9xPVa0AYlsbb4hhRhUQnEfhMnxzoQZFA7M8oq
1Rtj7RrEhhRRcaEkQDfZAyHG0kQr75PiTaneoO7JVUAZAqn7yTM0Rl4ywJst
y/aJMiWV+HiuY3MJJ0b1KmNGQ5lDERzycBQrzrHIY6FlXUO5tTDifzwH9UxB
MAsIF/gHcgZAFxUVet7zHhuvCZ6oLWdB6shHpjyLf7tvbLH6FK3gh2tCdFiX
3WhJzxcERPRsoG9bMbKToyHEq7Xvn9GOqmuoq26syDemG23LqlkrHUAf49My
bLI5DmNAdz/pgP1nx263ZsajrYyc071qkf+691lQgEIyboyA+acRfQBXTfGi
UbtcHWvoyHp/klma6CK/IWlHOz3plC2DsHOt/wP6coZroeb2ctvq7ILiBNZ/
rgC1Fd7/+2BELlTwFpFnZaXm3zE8iAJcr5KgVbs+JKq41SENQWZsry8JoMVN
66PomBVf3OqgtEk693J4vqfZDZwT/IYpFroL/AbRiBhXgEGIl6YoVi6XKn1w
l1bsBD1FJ+1cyzPrwzduEMRRP9OC0AuTo+iieS8PGthJBHjXg3orfVIdRg3J
OiPmWnuP2ZDFItylbum8pZwMqrgMRxrRnmUos+N7hRMZExUthrrJ3tD28YFO
fxXyXAmPKJSJWJdXH7fzn9oLpQ9jEIdd3zOXsb+UJ87BCYuwShGeKS25X46D
G9obXXoNCBA+qXXBjj5MVVkxL6ykJZNmH05GXc6kKJNyGbOSdh9W3gu1CCP4
SV8DF3RN2qaOdyh2ke+EUExZWI+ek7vYJxLly5Fxx9AICL0rhSq5D4AcxZX+
lwuBkGPOEdRBKWUKyeEF8tnm19uzsXhkWx0D5F9QLbNOgzhBZYKxhPGAaT1U
/DljS1mpVm2PtPLjA91OyA0X4tAyBY8lRKeUM4IkWEHsfK4sP255fBejyZau
cZ3mmOre1gGTIutjFIL34Ur/+9ErhFgofZtAJCr9uHT4aDgRWrj0vfbp+D+m
Op+83N+U83iL1VH/L0K2D2XwWR3nt8j2g36dkvxYbh3wjO95UyVhNy9SC2x0
xlp8i5VXv7D4KVn45/7Gl6gMcSTY1M/T/R7HdBRP7OF+3X5n3iclQxtvHmxt
yOcv3nRQ2BG+enWHkFAFIc1TK0Qe6+VOVdMZ9n8pK0h//WKNYdFi3DBhNPQl
IOg3FtRNIVx5FE9ZZADuC8tjUkwki7pf/Qw3OzP8h4bXVZ+esRzMJDnY89KE
e5lnOzkkc41/MjEfUKhWoRRQT1cyFuao8JO4Sq/+qvjQf3Xj8jy6BGfQW9j5
cfVjRYVMMhVkuB1zTV/h/7C2GQTStAvnmV0qQVK5OQILjpdrsWQvf0pXnYpU
qTLdfh8IyRL8h802zL8JJv1H7y9tq6Ak276BrAREnZTy5nDiGqszj1r4/CiU
xwmXp43gci8RMfIPY3k4lS8N1O5OmxF1AQ5sg2+7XGQwzeUOU+Man48U/+C6
vR2CrnERCoVLOn2S2PuIqPgMCzLaVMkzOrOG/qKaHWXGqhJsCKRmeAfnqCXB
AW/RpfXfe1KKSktOJ5XM6wqGVQbRn8+Ohl/6uFA+HkGpKpM5nsnDtg5vmkrZ
VjalDPhauuw3cKzSJwZ8QMvA1OFU3XNNUuRstrjd+lgI0XySLI6vsLe61R81
p26bF5h+3+xvKNKyBzcxx91FECix8HIr4wSvXtODCLP1mQi9VCVCsDldWNFW
SaeyxcoPVcloep9JJDDliObPfN9S41uDcvGrbXf2xv6tV4wYlcJK3jd/Z5as
mFXK3HZjfHdNND4VQ/x5LlNWHjshdbgaCsPRnQiieDSBzJwzZeNfkzDauZB4
+j92z3dGeK20B+8v0CRvcE7InT4F5X8puiW5a4kM82X58sn5He1249T6ZsxH
n5G03wy33UXR9NgiX/Tvl5w44Kf6Z5AFH/fl9eC13ddW8hHSw/NzFn/xc7Dm
2duChGwsURL48P4G18xsfSJk9r7TMQ6Gbio3vA/eH5udN2+B5b/xq5uTMq8b
mVe1ERD2hQM+owuFrqbXh+YwHODYehlZ6NH0f17qNXvU3A71Y56Lkg+AxTv1
D2AVhxB3bx8seE6B2vtj8H9B8mcf1RT9TilGqBiDygbN+l1xpNJahFQCDF/a
AJTw+9enq87e1YUuBJmV+lEB5h6ddx+28aCCz/ROPPNbAj4GKrl0qfDgOKYC
fL0YAcem4xWpdbYNeQ6XqZF2jy7I0Rim8Mz5iw9/8zwMWlHQAnOMInddikr5
C8Y5FHM3IUYyl0C+tt40pD98teVA9wIxZa3yHEUDs59oPjC30pO+03GavXfD
O5T8EDwg2mQPEJp/ebWZm7f1afljiOzjYOZ3rAQXG27gpI/BYwX9DhD9IroI
mAQqRBDv+bca5BH/xfxzQDMPd/Y750bGpEsCNFcBg8Ny2lPaNvXD5PcE9Re/
1WETb3Ikr1/oB9BHYZWz8PosJh2BLCF6QRbDchBuET1+1AIYEAxoNKHSr2LE
+A+oY6Y3NcDIxUc/n3grbsMNf3Il79b1Ls5gvWcSpmiT1dPAF8g3qLedEcBR
2fG3MV6DSJYAWO0c6jDvHhTiJ2RvfcjJP7slEG4YGv6wOOtAcbS0a0gEVKtR
CUMSMiL1O47HSHGbwhBkRGe/JVqWohp9aOoOCfbOz1Ac0vdQ4a7u/YBVOUT7
EvTWw0PmRwGYp+6Fdtr4RP/7PqWRWoDtmrDQvPiXakeod++uE2fSgHZwyO2r
mtX7giAKh6hQxCgdT3K4SVXnQYbrUuN1bAdsCDapAuNyyc08/KZUTx6kV6BR
MvZdvtnau/OKpCaPPYwE3xQTqKFSGkr0fSW8iZOMcKOx79WXvM5kdKDBZ4Ox
gMZN6hOzjfk/tZojPMidgpU2C4qYwgRtA3XQR3jPLLU5dznuD8S8a4kF9g2U
0pDzROqoAN+de5sqUfSX5CeBArKq/LUzDtBJll7jC41CU3+7DqqwdQiupTKN
LZZalU6K9YPHS8FkTCxswj2QzZOPNkI7osbTavNzNE2c4Y8zDYbtHjx7oPsi
VNxbrLVNstoh+BhOoODeVY+Vfsk17aUnOy1yf+B+7d9CCsQmIw5t7c2HSHVY
MR5KTHujkGyJOuhOi9TtGDQerwijPIQl3jDvK9S1UZimfOYuyF/iLcBjnZ5C
dOVWo/hI4zKNnmIE+5UEmjHjYRKvVopu6wcEioPcB323mOl5a23EA+JiIXEe
TIUhvWgwY3oshf0L1mxBqlPhmX4W+sxLqj9BmAyUsK0ZlRm8uUSNV1/VMhsL
5s17MuLdNtJhzLm2+69NmKq5/y+c10URq39aca2Qt0D0RwycislPs5n6SOZw
pWYpDxRaQdHJVmoAkt0qzQMg/7qMmyPYSUeQ2xw13d4uRf0ra5ShnrisqRaz
OKpPnjd5BxzlZ4T4xR6OMgtkMfKnHbq+3tFvhdNols+xvPyQttaDWdAQkIro
TniF776broI/e/evOKY6se+sSasHfFc8kfbktm/TapjgIrRfmdNXvsATirZb
WIW6QtAdD1p342i2zwY/7z7/WSmAmB1Zg2i0XP64dwo7M/m847dB/XDhYcIC
HwNMTdtaOcio7oO+IpoaqkTFNSSgi88lx8CfzMjvOJ0vi0lpcSOSQGe/HJw3
eLkUtsqg4DGJpdzGRXz6oojcPmbk+DYTsPSZUwmxB11K5AOgzeU9lUe/6z3R
gmYjFGaAvE850df0KBp7yxpzlWbgcFl62qH6O0GZq+G7M1DlKdcnIm72Vcb2
aBVz4hAcy9dY9Y0w2wn5pji5nK6Ve7NjDowI4CUEXOh4z+oy901A9ehif6pn
MPookkKzVd3yH6z4YAzfNuBI7UfDL1cm9x8voqwNYXmO8gQCwq6bL2G+sK9j
gDggqb+tdFyTyGG4rRObsYoa8jo++WxV7de90s/S7iDm5uKwo+7KqpEvCA7k
Fs6WL+0c38xfZpT/PO91DEztuKAfLZER4yf3JpnUY6FZ7edVIu7nYSlD379J
oWybggYHhMynxHxyyKF+MLHPWKrlJbDXk8OXc8G0BS5Ruh2B3bc3US/GmS44
4OrOckaIUwG8ykF0Q1EgWr4l5eewu7VXvwSJESKRsM1ebZV85x3fn/Njz5XW
PkvcdjEPRgHwnaMiMhUNUW2SbukuOClO11aSC38LOdHAHVJN0ZVULE/LHk/C
o1mrvcEbi/3Zc5WsZ70132YsO+SV5hRbABos5UPKdjaDcanHHwaX263BcKCc
hZ8HSuY0yP5dqQCZWqGCi/Yjtu+9KeAKREtvoE6t2vOQOQ44Z9BW1ai6dZhp
BpzXJF6sWTRAFOwo3DOcT4t9CYmHiiPowro1sfVaBrq5JPTYi7gXpHN+3fqe
fadAN5a8/FYtTdziJWGgF5cV+ZSFFcTKVoLZU/Au0173TaCDJWGr62pNym+y
6Q5Dck6QCbyYQDO34T0xKzjWPyW9uG5LXXpYPbJHCJyphDYQOoOnuIJGtO8L
/1dbWIwg8AqJVJXMFD3CBABNqVZRaMbdubfa2T1ielkrte92/1vlOiCzMDUl
zbc9mgzX8UuUZ7lqooYnT+G3PPlbyiejRfPnLAxSYguEm3rm6CNFJR91MxqZ
ejVUXqcgS3G+79S2DmVtlijPldbzHTukUBxo6/9yt9yhGXxIh/cI90u7qfkn
hK+LSdvzrJTc59gRq+OnP6jKOvdvdUluoibccsqB6kneKwrrK+KSFKuAfDQp
z4URsAU5t1jpr6uyeJmboieGIAsUTz8F9iNjLiXvyBJysrrqfKGPsNERZh7S
5g82fXGJ26v86iHtd8IOHX5UfVqd3j6RK6a+r7/GjtXEM378T/+G6E1iOQAQ
0Qqyz+5OqxDplvUCRQ2qBdxbgepl2maYR8QRm1lgbpx6BQm4U3covJewENh4
v9dawlL17R+E/R0lLXygsS6TfG5KyLjHlr2tKF3OEI0tn34r24yc7uvyGQXs
3JHhrKfKbnygvnXRNhwZp6W4j58NOmMysUxaHTYjEIsMlNT2j0Pftenlig8R
zKASrFwTj+p1iOvjp2mRJdmyH5GdqxBX9ILRgojAQ/46EISYs+tmj+c/MgAg
yTk8We2heGX6xfAGniB28g4OKmvyPswCGpsuagR6uJFDA6/Ps8j/zg1WgK4E
8iU9OgNB457rOIgojoJCSOl109VHzGCivg0/kAtEg5rXOyqLj5p5WDsti7+e
p/7SkMz5fkLY64q8mUTZ213yXncRUO/Ri1vDsWCGz3yTLwy8XZ6DCb+D8lHz
N6QWmmoA4W9QNpE+BGZLHawnnxoCTNMEtVhpxiFsEEezOBsNjPW/CkfcOQvb
Dh5s0/ODJ4dAWeAJUeBlIHdEHHeWyp/5760PGzarn1d52AI4Q28O1YJcjiBq
6BmUtM89Wqmb9I4Weo1MFds7q+0ee3myh1vCaln4mF6M9zQOLT+uIRl7fa42
JXvajzP3BJtwtpEc0H6cnfzUuQ4LOyfLoD6ZJQfXUFr2n9m5hEB90IufQnG6
gx5uEtJ/d1rid8ivEzIptj/nyLPd48P9O4Sf0ljbjpFVYBTzj2bXGyHzPP3i
Q1rz9DYqx32cPoMiV21tDErg082CzmQa8d7wkKLRcx0fOt9GhYleMoVzY6w0
IKH1J+5F1fbmWYM12yNsMEo2t+bZWRa+CPPS7oE+sZzshMBLwLs8e4oRzPql
PxByfAQPbyHstLsK6SRe/KZKoZmiMl+4DFP2iY2wYvxXkvoO5ZBxt0RYbGY3
e90lC7vVTseQDYkRFfLHIcK7PBXgjaQS4Nuom903UDY60MSGymyxXF/PgseD
C2HMn9FREVXYG9GyPrU2jhzNBFaSMEacICKXFUNpYxTLv0SVIcjOWYsORI/Z
YTuStdhiB0IWv9eNvovCm1K4B0egr3uab5laY5BiWWKSW7/F/fWICmXRrHDC
Nwv1+vToCElxH9RXIHRBd1FUe9vHKWlKl+ZmMPKaGuXSOg5hgeQSJRBoeLFZ
4a4rWyVLa38STzmzGJpjzNbWU8G6mop3yGpLNkooRUlcP/3jK4uComdICUPh
X4Xj3qHjUCJxC/LjZl+GCm5qwxVtpWauHOjh57kZ6+1gATBTAGefbayEfDb2
WuvW4MOkyhCVlkNfclG6fmRrBiTjEsWP0HQmRv+89XSQfKoQ/OpjODuIN/Qr
sjpUumPJOdxIU7KJdJrWc//dnZzdMK7KczR+ik5OHAEgE4fhZhj9UAUGeUZ+
+9/r9Rak15bN47gxv8g2oFe+uS5p9M8j8dYj87f4mu6QfdA8qE+eQNmPP48k
44tRm194aqs3Bd5dFhQubf/PG3WQP7GSNEGkKywj8CWyRcDwpDpVq4Pv1EUJ
EQyyGy3Poop72xzdC+6KInneZukgfpYBmPIKbT8HuTFcUaPatbGSkl9OrhAD
A18Bv+trM0uUNwE1ZyBwY9nyQv8IrghKVrf6sFPMM869i4w6v7WSgVsk7dum
5I7Q2sVOi+ufIKQ4bbqz4sWlFJobw1D7t2+645OH2AdqcwWq/hA8T5SUgmaJ
tx4XGspRq23HFhXfvvX7rjut984lx3U7P3T7BwnXiApdltSzBD/ozQSdsqjH
nGp3G7uHN2lPbb3AdMANoOO9evPnlsCFijkxPHnX5B97jPVzPXmD4hQmjkbK
u9kPqk4mSkjewMI/CeVSoq++v7pAk5WagkGgZQ1AcT1NGQYPqouI7GfjjwP/
CI4cXSYQsMA9BEQCjI5vHH81I4wMXLEd6nuMmJsOk6qFRX516jk11K9OlLR+
BTQ/bB7NtRyXaRZzLukcg9fBrXkhEJHyDLJN9pXY6Z/n45MjANGshfRf0jsb
Cbe6RdbLiG3iFCGP0ZI7hJnoPXymlF1Az1GAhaCIyii4tf23WoEnLrQ3v24X
WHISaVohPfGKKe1qpiFtek87u32GE0lzTkPFe97j4GP3VA1KBNE0Sr6lktbj
27FHqhttRwLWj1yMonbUvZlDRg9U54QJm5dmUEm6XvnE14v38Ed9bjKhfEAk
GI3yB+Ud3NOvkaUKBrnkQ8FzwnnkwyC3vBe8lR1EaY07WIyNmAvZ/EBnxqQn
j8LVS8tNGyoc1CA4Wy8y6qQ4Sf+2izaSrIMsQtru5YDml1p24KmzDbmH3P6y
ar5lyPF0pqPlcNpA6JBDvkhhAXUvzB3jxOhm3PqVJVvD/YBJ/IomCKZ5ScyC
t/CU17sx2DSa1LX+Qvmt5iyNI6B8T572w5+yj5O+pUKay0doeuzVuQGQ2Mh9
GLU81oJaEJUFgdjWZzuRl2td0Gm5Z3yFF1U+boVc9RBYcU8mKOknqyrxPL01
V07MOoB4dUf0R8q3/Ve1ry3s4OpFqAMMRtRwVwbJoCiom2ztRCX/QY6HNrVS
OdfgZktXRKXxQ55qjOiOjJvlR3lAnyD0AilcxkvJa/yjFxVYVpGpTqDmWajA
FKEhUh0e89KHemsAeKmQxTetpc56RPynYjayO7+yueBhQOwboT/INomBYWSK
Obr7GoyXxSGJ9xy2u5paRGf+K5qbulAIgO48Mp2DF/HMXV9bl8H8noh7ozc3
bgjSMM1PY/3Q6p1iP1SYRiEhqrJ9YGyB24dWlp4N59WBnN1pWiMUDqK145vR
EfbcrwRg6E2YW6jG2jH/EUgXnPcvnkSNNG5oVOwgfg9UlWEk7q2/qeiDPx2Z
2U/hiqU5QwJTq1EgLxD6bLZRTGn+WU5hBmDmiXfjU2vn077LwOembd8/fg/m
9IQgn9iVbKJRToEqIis895bML5ae72x4j6VYlC+mjBcCNY/oV/v6bbYw95Nx
4TwMQJ2Cx/oQHAdKqgldR2TG40S89Oo4dDF17odH0+zrYnu+FWzGzde5AgNv
GgptucuyOpXSTTgKyEIguvCpuapsMgJzVNGaV0oWCEyZ3aBRF2H5Y3LawPpe
tw0mkrynhS/V0WUcfBZvogJa8iI0IDsdXH02EXsVlDO/SKi0ecElgqYeu50X
OkfvvIow7746qLRFxg/yCPEm2KnfnExgwMec4Ke/zPZMZrb+xZc8g0mYCDhs
z0qvwomGX3aOGsXL9S07BL0qdEQiEBj0ekfm5nfXCi7oNwldl+4EKu9R4EdG
AAhIMhXMRLZXgg4niPpA2Mbr9VneRglz+uHK4KyINDXlMLlBeaRXVs4bo4y7
qXs69r9bvWlyTKyOja17ZqqMzczi9wwJwm0PIb9rxBWH1sZLaFOonv22IVFj
+VKZEwBgDkw7KgfTKqmsfrDrTsgUpdF8eNcL+CpUUztfPExxWIvcqc3pP0T4
JzwYtTqM60Da9vyfFSRFfWR832MeyeR/5p13bx9ypAht60Q2qx0PB3GRn7k/
6Qc9rsI16lrKr0DVXZR02hO7duekES/2uLy59SpYaQSsubcvuFaVyoG18oeu
69/z53F/J1WmbSqfHg9DO6kD8nIY/MESGGpGcuu2v8sLKwJL6yDZIPgHVztn
r9uE5BC7bXhb1GMlbOQk3+1Xrxl0AuqVa7X86D+Zq8kkDGL2T7vmwTSHNk5f
AtDFuIWf1sfCv4ZuL2fiSj17DUH48nmdY0JCm1mFt8pmcTUW9p3JYCPYK513
QRcoQBgWu80pIj2zjz0xrQyeWYzcJjz0DkLWsmNAfnBdUH3xqEltP6/TLGLy
0wHwRBrO0L1li54gtx/n8N5QJO1iQgzblctTz69rUd1p8Dlm1sCYqy/Dd1Aw
8K5cBOAG0Yx/KqOWY1VNlP65VGof9Bx4rzNaXxdpd+mC/m2acXoQZ0GSunSh
saVotxtsLou8khBNUOguGWrJp8/l1wuFGOeGlfNUMOGexGksPOnIkTPdJDKZ
S2a12+3Q63tCrB3CrvOKDMRqlXQfrkBUFBOdfU9l4wCqnaO4uShLmzHXhL4R
V8SuXAjr+kadKk1mqDpEh01Rx2zc5ydPemk9TBXfH927tZyFfPTWjJq5dVu+
g1/bW2RA1/EzUkwE2pVlSgiUEANBIRUVpZW362G0sGbx+W4MWaq3Jk20Ga9Q
+Hhpem4DZKt5RdPfNg3oFbs4y+UYdgbuU+jJUayeF393MiRTQmO7PY7isKYv
G3Y88dRcc/3ehlr+uMLHJ/cqGcacdYcCfbgdV+cWZQq1zcQ0LbIh+F3xmCy7
MMSRtY5/7onMr8u6dxMTcIf3VoGOBqbzGFDyncNSoFN92+JqzsfYwO+QGv8n
9DzoulZcybCYVcNsyYZwi+vgF1WbREoUDu0MaAvqmA6fksOdCwLfSShbJ5Uq
WWUuyyX97jfEUr2oSguwnNMTKUCcR/6MWrgM6CnlrfTAI77UOpVNKavI4jA1
HsmfVj8+8P7FqC1uawi6ErwfTZiNJVzV17d+kspUl05DKjgG2jILKC430zP9
tRZkKZ7gYGq4nnvT2sbUxM18NHSP6Tiok2UIzveeK1OF/jtUHwjxHOTfHNFk
uf5j00Aljfwbm/x37nQP79KmasIyD2FRvwy97U6mS5h9txhZ6H4av4b+fJiN
1dvj1/yEfJZN8mK/P/AAgWIxSSeeBrI/m41uMyC3LYks7Sf0bxN5j4Ft+tN+
1NE8GVIsr11bpjRPkR1ap09c55WrFnE0t1a3RrN39snJmlWNs8ohYRZ+naoe
/JohQvRBgSzgmIpowbQcSkvgGGdxkVu8xBsaaaYsVOyKs2g1hEEnzgLUqGnA
ksHL4a47+ZD15FO6y2ApTcXBQlwQMY+yzrrcEch/+2YLfT7SAqAwOllplMnl
tb89o41iDxhyi5ktHnfbx/qVtVg7JgYXgYsZ3jmsTdWkQOAkyMka8Zr6FKtE
WbUF2Ef03SYVWkFIQ3JOC8Rjz3zWG3Od1YJp/3eLpSHbitYIa+IlI5L0omhw
OnXdhygj5rm6TtFuaQ16kZq+VyM3jENnZsejdI2/8YTstXM4cb2mRwvTdUKz
L9gSLnu5zsjzTzJj4+WAUiGvT4Gniht7wtl+5B89dOKsrHk6pOqQlpVeNgt6
NWC5mNfFv+OXBQhpZ3RZVSu/PvAlNDZf6XYyC7EmopzktmtptLksDpp8o5HL
dg9848VRFyzNxmfhVkljK5PDr6vHv5gtC/sqDPdyUu80XiGeB/ekVBJhfV8D
DGNI3aJ64DK6fcmHD0AagPmA/4cEHq0zNsIFN7ojASu1KVO/6baP286SPfdu
+0yDTquVpEnaRRUbtYlplN+NI/lK7xLidzsA4/E63oSgMVerg1yUeS1MF6Uz
C/JBakmziOTsChuQhStN797bjkOd5rWbNk06Q+GL6tiQYOJmtC4y+AQcSUsa
jYDw2uUIQLyt/2431WHxNbhy0uFY08cmwrSbAOIc1YpQnDenpbpYpeZeU6Kr
gzymlInu6t9NlKvdLvi/oX+Eyqi50rDQzZ2kzkb7a9UWK+skFqBX8UaT5uBx
/Y5Lv+/JwZl2NK2MgJr9Z+UIG7h3+P2MLJ+odGvghAYHqygBYxOBN5OlFWo+
+IvmPHZhDjh0dJY9X4eXGJ+len9BOEP29MqLAJLeQ3ScG1CUMe2PuYJH6sqY
uvMXeA31eW0v9+cNist6xLj/yIGV2IwxaNuOONsfv8zD6lym4GRnRALVKRp4
KUikywr1QLESJqsIUa6jOeg+/vgBiBcuL2L8eiJ8XpnPYhm++ieUUQuIaZbk
7dGc4QviHBkARi7zOS+D0yE7k2lVevRgZLcmYdNqVthGSQpnAwpGcia1PSMV
2D0zTiPjv1LfVdx1eu2mBGp5Gmb8KqxXjI5QHi0oFZTWSRiuM7kKJ8uyBmKC
xTnMb+ySmQjBDSDg1Ndk8F1A5BDN/Wsq6PBGOIFd9VUKYd81BYfLU5KVdWUm
nv7w9mD9zF9UPKpK46QXHPHCdgSUImQE5K9eS7z6ZeK6cthZy4QpU8yxFg79
QsdHyi///Zzq2AKXo9u7breqicHLTrYwr5c6D8XhD/YCyglx8O+l/9jpxjLL
KlKC9g/d94HI2qSBIH3GP7w6FChIVOjSXSlmzXfMiOBANkYcU6TjeTWMhCr0
g0LWxQHHV3Ba0mgOLTk77EDm0+5/Ur3wnAxP+UKZlKL9XN5nFwap6kUQ7SYC
XJX58NhSPLBMRXjhEN86yLiHCJ0UTE6QIEPUj8rd86EHaJhVBhNRt0qTTz8h
YPK3Bkv9WHvI6ZzMCHKozw4CwjlR8kMnovM7jM7AR3aecCen30onnoXHxUWn
YrclZ4J4j6a2pzpbSdnUfni7uy4f1bLs5e6sRsqiRvhIz8Jx6H7UhQ0Q/PFl
ddM1/EDwOUJ7D1nZirmDZT/heMr6X8yTYNmMjiD7E8YvIcAl3ZiMGpaLa5UU
9Xlcc2vHwY9kkyis9aEOu744rVSHl18enWfN+ck5aarfiNqyDxUaEqPq5qev
aMy+oXpZA288wbpEt/tSoVRKuCVoestTpn2VapE6e0FJAxdADcUBZJs1tbpB
wlUlYzhVYwtVhNQD4HSZmy4v4+nJyq7rs8MXgTq54ZymRLF9NRHaJI8gHzmK
BWBV/CfuAGgysPRShTlVz01F3GWhKWboFR7vaXBm33CEi8XwP9+HumuZtlPu
UeztOpi8yntcZxP57GO5kLNDLNnTOakxAI0M8hl/4I40YtuRb+1a0MBwhsSA
ck9/Uh8ZuJvX2Zvd/s30xvldNyomnTTPmvF5AMQRpaQQnHvOGKkbVoPPDD6D
Jy/GVaSFC+pbtnz46vNxu2Km4ikdqFv4zQbtfnYKVq0waweYxYepTXyuQEmD
u2Wd2TkJO/p8YhDKycka4809PMwxZJhmXo5kOv6hn+L+UH6t9/wtj7xiyjPb
36hI6SRqGCEMMxBE+lBRcOnboWS4Svx5+v46apNvJEjGNuX1b0lugbFGLRf1
/skNWjs5+P0Wsggkbgvnp9SPg/9c2Or/wkNxqSVKUEn+gKQ1QUmMR+AjZrFG
nl8XnCx012jXHXDA/PQao3VTHxvIebkgIgttYBop7ja5gWirDsRFYFmCO+2h
G5YpXWXPvVoW842AQRAskDSfoBVau3EsXkeQBmReczi+TMHzVybPjCI15qUe
PDHOzJGlczizGuVyVkprw4jY7N2YbuZEgGidgmh6c5uF58qQ0ejU9aSvhMi2
UxJ9eZvXKvlo3CecdR7j8FiDPG336sapEe/1hoOvHIm659KG3J//ZBFNDpEu
3IKlkqJlxoZ3g9KU/1Lo0yYyvIyiLASixwMeDc/hsJttP3F3O5ALA5UQRmca
1HtRgSAm00BftI424X/gQhUbklZZhnud+2NWl5TrxHIfDd2k/oLTi3Av1qKr
pkiyEUNg5MWMjO6OX8ZoWqg6r1jGuPY3IREgEvqTLGW0lEefGaVYmi1V8eyL
resx2FtiWFbndq4pNQ4WXYAa0JwwwtqETSqBjeGBk1pgId5H8kHLsT/6G7cS
ttpe68xLf1sG/CvEnZEl76aCKpchSFZgGVerjQMFX8a4/ahsTg89irDLL3sR
cPmykZoghv8oxFq8RO8uzmwnBh36z0r5oiucfLoU5BgxDEvFEnXqkqnuVILM
HO/4us3qYRlflJCbLGiYgs/FzVrm53WskyHmOyVZ6bQxose7STLyqLPvSJTT
E7ej7X+Ok7P+niDFmyUWBE+Nb4ANzpnSDAIPqkjq5mJX9OIQn5EriLGa9Zfl
LIK04OYzOYI0EMRWqkehfCLc+8N3FpbQns33xUPQp21mNWs8/0UH8gpc0duM
glKG6WVPx6zVFhX+QIS7DIPwmu+9AfPruMX1x5nMB2P0WkLQYiZIMXKPub1p
9LH5b3hwAOctOXGfhkaLKTxUv7rpeT+l9ON+VfPs4CQ/dFMRVT0UIDcgJSJv
qL7wxO3XjKTi5EgfrVWBqQT4ELU5EaAtYZiDF+7UWPK0y0xZ8ClUFhnibczc
1rdEzZIi6t8tqc098LBXl5lRHnuyhuG9LIQVbCjknievEfjwKTFKyQEgez/U
e/MQ5hEjmxoaNfwH7aQFB/xkN26NOV2Rkj9wpJ7SkOMK4cvb4/TDs4F0hQC7
TB37N4AoDfhLN5dSP87NlWqWypMHiiuRI3pzJjKJCv2fyS1AQ91uixltu+b9
xGLOWk4DhqwdsPkVUbM2nUQ7EXq5NaSkbsXpCiE0jbLfbhcb4O6EfHJXu7To
4uJT5P1MrLgCsGUlUUdVr+paxCQISuB02jTVZZHJXUU50ih8J5MFVuW7BmUk
0ZegtY+w+QbZ610xLdMyh6EvfyfxqiSJa21fSLdMDqFjfUT95MGkQ0eFHpJs
2VJBwiMVXuCrdGcuGysFJvY/yUvfqIADKd1mDkv2hMrVXBgTN/9fKZ9lx7ZJ
lZEGWrGOZvlChNZ7KjPKLiDIwZ/6t/4Z2dN2N+UsPsbUDPaNRlY1afMyNf25
JfF47bXlPNG/x66qXAyvy5Lu4ICFKoHMVnQaHZ2UoCXI2nHLCGXKsoCwz3Mb
XvcEgzLTdiuewMSKH2Ro/n0jlAGRD3Vipul92vJ0Pc2LGVZ+UbpH0CJaP+2V
osoNw/MY3J6YQXgNNuppKNeKOrvlxZW+/JCLJcX020OGXCldhwe/lYq8qKjR
/nRKlampLbLCdkSWM8d6caFLJeYW4at3smRwjJU+9dn5/nL5u6ljEPeNnntv
9oIIxhHsXhgOpthhxDaHDpIHfneA+zHr9kUk3r/+mOdrdb6Yoc2JSEhzr7Cd
hrFpEFw9iXT5LOqvjUZyVSWhm1VHD3f//Jv0mO0M7KSUCU7m057HFH0zgjix
4Ej0Fk6KytTulCIPa0k4easft+Ox4FpVk4WufX5CUh3+qpAyvpmYr79ulKEi
onLVg6pOdGke9Fnf8Jf4mFy28QrqdaqYudf60ilQXoirJb7gxptdheVmm8wa
vm+S7/18GISxrVD5l6poeUe5umePOqjqpt9y68/k8R+sardq9WKbtXvP/jkJ
z6D4zI4ZrEoK3NolMw1vgZK4d2iC3V8CH2NySHzAZ67iT0KI75WyIqXGc7UD
6iKfiIWIk3J9sH+MvTFWKFAqBe/+N4IQ7ioKlRC/TvBCAJYPQN3Y3J018i2L
RKKdh3aGUKevYaZghqGkGVgQlhM8dWAo/Hp0YMXMYEq8Rf42deGZhowNHRud
MVKCJn6UBqBmXK4X5Lb7Oaey9uRkHv9xfyFQAgGIsX2gSKE/BHDsznin10LP
KbfCkS5bnak/b/rb6ViM4Rv0u1wqaZIzoho9nch8ur5Tqr3bbSp+8rqbIJob
V5BYfjRrookSKoUQx+OZcqIdAkPO60Xby1Eizv5lwFNSkgyY8pZ+OaYHLANY
wU9/h5HsHMh67664MpmVuEVe7Ba0QRaKC5qdWLQw+zAO24JVxJKtkicX8C2j
Y8cDJFAiAQV+/wPbWUFLH0sTYde5tM1bQD9/nx4HA1Sp2dfsjgfpeh3YLXL1
UOrfVDltLmv3aBe9x6sqIeGQTcH5L7jUuHuA1v9cQFLd2DUCq3oNVhMBmSJ4
hag7/4uaIY7AABWvNqRZTF6U9cbg8IgdXmRtKnmGyO/zaTBls8i2mbMNut7o
BhK14Ea1l4lyuWAWKldVMSAExlC1/3I8iJ28S38Bnc3pDphfP2zk10LW2vqp
70pcCYviqKU9Vd142aslKRzG0w4XpBS5VYnnzKNDc0gsAFnq9C+UYbAHvYyE
v/DsacH4MK2lQtj0hf2kIUx25c8TzmOANrNSADY5Oi+qAhZ7NcWadWXZ4TZB
pY9VN8s8oNl+RgsEZ870GyYtJyATQLrl+B+u/LTdUY7Ccg+N/vrnZnQdkBTA
BFkBboBUyxEkbVrFARYtCr+vN8LTxJYXa3MEcMLq2xlyTPMWa+iq+ZG1mv3j
Mu7IzrSEJd2HPAcD048e7JPpdYcdD00klcY0rvutLNCW8vCSChTqDrw1ElFF
S6yyxIRmb9clc/hEo/R4kFqtIMJBmmPkS+8I+bZQ0i0mfgEMgrHWcc3DgQ/a
V66sSMQUobKXc2rTdiIp1R8GE67VptRlEOqhkh/7WmqxTmOwqdCQ3W2diWQ0
GJW9I4a95oGAHD1nfucEF8yfu2rj+G19aep8JQCSybrA+5j0wND6N/zFa5vq
fJck6GCadXb/+rgDhUE6Xidj1/k9BYvEqI4KSOgGOdsMVNDD6gzSEbnUimcD
LfVZMQHtbY4EZicQUv5MN/lZaWMT6qPpaLrqHNU+NmHMMVYv1OPNmAlG7EFi
YIlsw6p7LUR7ZOfFICf/48L1zJ+GAtOBTAeDjzOwmyC1zPYLTmyV2xcExR70
tqNZu+aO9h06DJfF7Fc8ezqBh/0Rx5+Ne7O/GFszjiHErhnSBN629WnEEwlf
5EXPrhX56fm0ynjX7/yKNEiOdDAOVVZwVRf3DSAfaA2bBsSqL+fv7Zaa1CnT
JjLd66t+xciZNFZTtZ6OuagT/IiNtEgcLmMQPlzDUFkJNf8+CHOeoLg+QQd3
oi6/arFrOVdNmmTmE0J3qSmW2LyElJpIKKDJDltcP+mnBBG+BbiG6OxCpK5O
l4utEDEgoiZ32Ss6LZPdNkZSeyY0o8y8n6AxSW9Da1h4vwBUErs4atp5lS6S
yqVrnNTeJBsuIp6WrzxBslmnlIg99y1SOOS/B464ZNX6LU23wP9dHU1KVZqJ
cHAkAIcfZFleFjGik75ayLi6DfCK+3TisLgep7qE9WG5bam1YMl1ADoD4ZLD
v1hwJVbyu8jOjwFnSyPWH4w7hSa5nKVetYKg2oig/n3y9HfLyxHbxLEPSJf2
ovUiKy9w8VyhwKrBHpYecvSWBKUS6+Sg/yc2gYgz29JHitRrbaQHW2xDpNaM
+8Aj/BkzROFDaboihd4AMEzJzwemcFEjkUDhQJKrD6BOa1UZqq7HlpwMhSmK
3apXeR/2E5F6MPOHdLk5R0JONIPeGyPIGjspxOgiopUne4KdUqsWNvYvAR0f
B/mN+ptTtBw2/pxUVDIsjiOSzryct1ptis/VKPkp0ui5mxoRsZr7XxjpjZ3T
lzI603qPiuIwYnphhF3/qA/rtBw7YzoL0rT8CCP7ZodYglemCXqJgAVS0Xf5
ZMLq0/uvsXwXKOKEZiYOuoz3K/7b6aiCABk3XdCQsbZQTlEc569MmC2N3nwz
kSTqO25CF6+pUDJUujNltrGBi5kzID4qi/KdJX7yoKdW5JYitKq0N8JExeoT
FonbtXGTxdvhNqcime2dJEe4lzXB9WMxKjxCJEtGX8+Ms6up5HvAZMwAIXiy
hq/K5A1fCXP7cAQTeck7xIL0FUejdHPHjH3YNDtz58Krl8xdLPFEhRMDPqMq
8fyyKB+UFg23F9z2pB3hU6k9I4E1eb1YWD49wl6SluQc8j5bWCOPI9GeAERR
RK6gsDe1xKnnT2TCEMiGgvkubGZlBFFJoi+iOW9G8duCCFj+BzUohgKrp3QM
OBxTyn84r0Z0W3pS5pBLPx/5JgONeYJSCk0qvFv5Z9X0m5bQGpp9UFDZ9Ybj
16z4OY+1apcPefwc5LFWzVSgoZemSETURBRlo7egcEyR9G0Ku07Xc3bdzNSn
J12T4KiLGJ8SNE8svSnXNwgrdvwI4dQnH8B6yCTE1IYpLndr63PB7IWZKOhg
LdJAh91JzdZXgr1y8ZdxQoqkQIQ0uCNTIfVEAPz4LBHZOHCCBUwBgKvXwmdc
xJvf16mEZ8iBYAckXZvHCVeWtQwJVOhR9LS+yg3avyZT2D8nN3oW7lPsBhau
RAHiE2j1bCRqn0+lwnj5TGpYWUn+9VNm0geyC1B0YtIx0WGQQrp0I7nfEOwH
D5lQ7EduEoppBelOSXEsMTfdX76zbtf/fka9rWcuOJ9cnFdgIerdwnE7h9FJ
8oVJgYrvnzlJAneJMN15JgOMIFUm6yNkniYSrBCVkbtjRS8PXtTJwVcBVxd7
DR0rb/4/P+VtZTvSBjLy78qgbAxIr7V2C2sJegHelqfoZPIPk6o8w7g72r9Z
ou0d2ikRvvCbw58ZP+tsYQkSoHUXSXswwxork2RbhPkgL/7PuSZoLpkRmici
M63BJz1wJ662MWAfzXDYXsQIi+ciq+i8Ab/BJ566S6cU73o1Bku5xZGoJ+Sg
3C6PTPnyzitKG6M4tB55QV+nGa2jETAAt0Rv/YuJJK4iEcO95ZhFhwtbLlrb
bwvx9vxza5oVtmUmHzYZkZ/nYJp5MFx9Fkdy8EVZUgb9BbAgS11dJUCXLG/m
1n3Oc2e1PXqdlVr6w60N57bo+HfthRfc7D5PITa7MgCZB+86thWF71HGiqHT
n2Ru6eU/om/HVkVGynkRQJbUYivV9QfuXHaBG0MIb/TchY7kTPm/IyZusnV/
wLXEutpeg2sX3mVlil76R6ff0g4XMv/OZbPIGciWTcK5hAWNyfIixBVwwI6s
9CNrbVrvIOf7bndzK8zzDnqymnH+SSVM3h121VGJsaMNOoLIfuRcSHWTj4Yp
1OoWC5f/iYhI/74UDxRg11Y2N1WiNyF0OhMGZpMdhiFGmIHtjsSQ7G6if/B7
m7ulD/LUQc7LpLlRd+sjGOh2j9UnrFZ6GbEprXDs4cTrTy9i0bLbHgGW5KeZ
oGLjgn2a4D8YWYq6ue3sarK5URnaxWO4QePjhcsFiHMQT0xFXmNitnAjmVPF
9iPwf+HwvHkXD5t4gFFxFXDQ6N48T9w5jp86vzXKlfUa2iI59bsuHfCm3RGU
ksMPjrfmFbgPyVC/egXJu2iTG3Wj2JWkTep4On51hGMd9wEcSCsijLch/6li
gvMiHEt6B9/Xize0xhXPEhmUO6D7m7qoBbhqWrydyGUxuwGF7AKf84VayYbg
mGjDwewges7l0WwNOIRk9xX+Qxxx89uwv4hi+5B34+AYt84MI83O9IAaR3Xm
+P0Zyv/aCbLuFfIiCiuAVO+jGamujM4Ca22XiM3zrEW/WZcvflMVWBxtkeSG
ALVR0hImJJafC/+a0BIbm7mN1ZDuAFs0otW8n3liRdNBdHn/9jUGmzXhs/BP
icHLOlFHcZax8Zhgfybu8B6qlxw/FyJoMr1zvZMS7Q8iJfEsDG+DMxpJTMPS
lA+RP5ZE6ZVHVWvSUcKD0IpobQ3t/cqHrO6Vxw9YAWAUZ8R3lwuo+Ky96AKb
MO7xbNT8HJ4pb6BspLaNxzRMwkqgoqML3Rf7rhngnhDl11NWWqiauO7ymp/D
QDyBQuA1eLb584b41K2u6bXoJU2sFeEJimaI6OpW13fOIU4Ocwk0/RYtSpMa
EJGqJQH1FtZCoUoRa4WFnbx5P+zBPKa+Toh1ZQYo8z4kzqMQf+rniKosZXTO
vculNczYP6qZ3hT8MJJC5HeTE90SFlkYpj+0z3otU6tvRsz3CyPB0Ek62B8/
jj4uglFB2QWOj/px3dA8QDXqpFhy6eOTr8RpCGQ/xFYW21FaGxcmPaQ6N9WD
8XfGzE9vucav25WiylWWNxsEeP66O5aOrZHBdun5aIpIXupKz2icmoCcoO5c
8jQMZahIOgyalcjCK+lgH9sxDeA7jJg/EfeH+v5ZZoZ2/Nv85zXxkZPg7acs
9twoTTnbAFHW67+FszWwxbOp8VU/yOFtsK6/ww/BkhIvyK7Tc3xexrovuWmW
9pnwbspGrjGPYQOeh1hl98+RFY4MV0We4RFjp6PCbWSU3/qy+8UUt+5kC7y1
+HmtFgwtREHe+fUXvVhFGUh8259OoCB35666t3c7mrUbNQlJ6jk8IL/oaE+1
w/dS67mxakTDus4THfF+AlI3xkARN0O8eNu9V8w24Sm38RfQ3ivEE673FbMc
8YlbhpnF/DdRQo43J0ukhPC99rkK/wu6tGKWX3cRWameJXHBc4nNW144cp6H
dBkNpfYI6fYP0Fr8xTV6cePQHjwZKPb1wKlVo6qhPlf2L/LZXIRmvRvMpmEF
h4Wq2OGOUMo0vGHcsEy0Cy+HnmedCnSy+ku3KnFLi0x2LFQhSiYrwvaGbcNp
eACPGrQbQqJ+1GQCqrx4pJH3pyhP3//mmMuZlNH/IBd0kYK9MJ10wMMT6TdU
lQjhCbxv8HDnPaoZFjii5zD+cOLHWpfJUeGEX/BEGJahSZlFMMz6W45nwSI0
bbrrLzy0w9RBWlJFEULn+Jh3dJ55IjajJHyFZpQnSVEgufXfFnM7nPdd9woc
1LdlpYE4dd3QzRBdK16WtQ8yKlzhOfXW9j/2jyy1bv90KYCt6z9a02NANdK1
fbMEnsG1CTqrcfft8/y7J/SEuTZyDop/kZ2LI+1d0R1zRD9IcWPmFHxMSt7e
ZExngmiuBvNkUGNVcRDDvw0NCJxajQiH1FzRUDl2guCeBfB9JC7GeqZXb91v
T9AUNEWHP5DEfelntrnVXpFjW9aYcfoQ1FIf/tpSQ+g2Gyr126WMWoswpE6Z
Tm7dXe4jeL7wHHYumZMYA7nUk1zLWFeHKCNpm2ASR/EJb2aEmPr/IuxUcNk5
1DiJYQ8KPhWpFZM9VSsVxhqjjgW2bJRkDl/z7sF3JsDLfffL2O9bfWafuGtp
9iFcZ7upGr1SL+kEkmKGa1su9Q5M+xtRg4zg9JE2Nxh6jS5bS0BAga9mIW+j
uulsszuCOTxtXEhW2BeOQzlgtOTnHUVOMbn/BE8TOWnwum6ccART2SX9BZxG
aCb8vCIJ5/6GWhjdi+A7ECpSBrzBkJDa/rgZTgxvU5Fv94w3kZZTU0h+kN6L
6YlBLdsPoNNCyoNKolLz/NBySkLRd057+suUibTzbL7jsUn5oYL3cospwFV0
z5kpk1Sh8uWqf9OpgCfNv5EhXQ/TTe/q1YkWSKfubpzBDFxVe7o/XqlnmdzY
zn3Y2cTV2UFwskoJk7kKBKn8SrasiQEnAXuu7OvfbD0du+wpeDBokgMfZvKW
OkTYHljilOOgf6PV7fbPoPWkttvfeX12eVxZn8zIWIbvPmYGw8MZdgb3um6j
8OY/xtS/cgCNP9tCvmVHCOM8W85Om5Yg3SXkY7veLwQ9ZUi9WCX/rGTeuMls
JhsxZBUEw7+0RdaDELnHGRUycmcTxuO581u15eMIQNgsp+n8NKnqVQkMYZ38
cyR5t+43+rWbEVqXJHDBEQN9Q4eGW+fUO3J4cvvEZ9XmnYxsWx6SryYLNle/
AYQcrbMcuEiss4AwnmVN63O15r8sDj+ypqA7Nr4zbiDaPp5BVCo18IEA0Xi8
VG49IOiPnFF77GdPnaOtRWQtRlB5rSOCha8BB/ntVo4YIc5AU8zU3LZIK8dk
tuQh09KJ1xq0Eel8khq/zZwieLU8aXPR9nu7T0MhwwljpSRfnDTgAY4/+wBn
s9KuW7UGjmx2yIWCNbFJ1bxTuKKm8jYqPRgXua7F/W8CWqF2wDN4cAmHDlH5
CSPjUvC2f1xBsd8Aw/ZeAFbei6H/LfL1B4ZD6v1xuUw8INDAk5WrIlZ39a89
gpc1tcDeYVb7BII0neJ0CyqWHRvBBsj0d8hbxfSy98NBvGdjPteutkuMDrK5
wcFzoSq0hP6MmNq2VmdwvZGfXdhZ6Efsb81DXvsausXtQRe4y8PH0WY4//NG
pgxSbbo3+Eoz0e2Sr1OHweiXGVEIcFovj/2d0g+F4Orr5KM5Yfrs8nsEolZR
po2uu4tAmD92lnLuv6q+9vPTEAazVniuV1aFcZeYj08bbYfFj/Ad5Fvck1ro
S4jzUwVO7fUG9hbBKqC47UYXtmNBYKUY82hLMrOes4Z1yS96KY+TEkSZGpQB
o3FgMmpxY5bIw52GaS7PHKWIV+PBN+jg0Muiy2VaU2uZpbO6O0XXsMdqLSl0
N544a1FZz56vy3any1C2c3bineybX2++7XlX7kYgPP9GQurAn0Nr3qp+O3St
KAyBdojKEIn4y4Q/5Cz4CKPOc3CzrWBJlCNgf6CfG/2cKxmuY/ivQKhGiHD+
UZ6ZGFyeyM83NQyBdbfzJGVMuYk5S+YYaF4sMdG/TkD0OI2J3OaLSEzIC8DU
djc/5udI9kXAzvU6w+VNKTBpNheGYkNJoMdqUMFjszbgPMrLNgDmXjR4NKZe
Ds0SLkf32XxXgkyuyVUuXWR4CeTWFdpXPp3cmY2L7SbyCWkkn5JDawk8QOgR
UeTheA/hrTJTUwikGekHEHc9MxqjQhfduwQsSAh/GSHbldqN6voZLJqycQVO
eDAQUrsMmGTUuTTt0rFByQV5dPJ0gbnMCH2vMmYVavCSr0HUbmtFvET+KI/U
2HwJNEfUlxMu9AcsCwGSmjj8sQn/9H3haNZ6DFxmbP8xo+1OPd8NVzOcchJT
AetPTbI7/s0y38jNzqxfOMIfbFyo+ocFwxWutHZpLi+jJ1qhJ8txlkjOU0y5
DcPA/ZnKBwTCqGFzXWsCOflfAPv/Qol7mh1fIj8+K5iaomtd3VqXBqLaBtqd
vXl3HdzmiKlmsI+nOo//67HKy7+5oP4lO+ywM707ybHw3UM8we62uAAC/GHy
YGB9aW2gAb2FiEYUqPTwqa2E+Hj2v9uc/CUKsc9+HceoIDMoqQwCVOSjqlVv
z0DmOXQvc7cfLv+ge72UJS4kU9Q3gN/Ll8oIO7pRKfEW9nyihS7r6MBWciSb
2XGzvnlkTDJD5X8yJumxt80DyFFhY1csMiNiDUvYq7MI6bRwU01ALc/Ufh97
6dimgawLEra7wPJ2LXU09pD4s14ZFVrLpAIRnFLSL22RLXoaHftfFVt8b9WK
FuDmf8+Lc4pZ2spdi9dHQZWwPPry5Bavud4hb0BlZcOwwm476BIMQn45QcSW
lT36jk353y8eqltszyll4zsYlqi5KMd9m23aNtIPe2m7zwOEX6SM2TN4I6d2
Ru8HRal3ZDE4JuY2fkns6Ag/RHs1mQRF6ujCJQyyo4XkLfRhmvjp1oak7pDP
tEfD6UvD8MpbfGLEZQgr0YuwzqMxR/dKvF3VvF8W1aYTH/x3P5k82Cs7QZhB
dC6VA1lbzbvWGaD8+icIV4GPanYnELLs+rm90Kvg23tlUjLL5Wr5lAlitkPp
zARctztwh55PXzSG60RKm0YyLsUcNXRTFv9+OCu2ceZhDvMLN91mE0aGsYr1
Hgc5diwmr79DnZVNk1xOC2SA2ZBVwnMk5xZNh/sIC7e2mpxGX0STIOD7knGN
OlySyuBDjAb0itiRe0YMXmprRLFCwjWPDUJv9HnfVzOXeUFYXfcWitTGhZNS
5XEzvCWIYPwdlaBtuouvryrTGLFd4I8YAHPrJaKkNp+ty2UJSOglNMNMs7Gc
QGWjxopwz064tz45vy5poBXKGnL/FBbIm5lvzAYHb3UiAX4109rltW4Y/NB7
u1qTs8JvICL6ROVdzZhGdV762sa5o2TX3cT18WDAvSCOfLAEtahyBt/JoWQ4
ygNoBvDRa+l5HZ4RKcWUF2Czu+Izi1mQzd4X9qypWrjuJ50xpZHp8X+eZE2J
5kUDIAavsd9rPT/Zop28vFnb5Gjj63WDRJ4CNOHCb3j0CXqiTW5hbi7B2xN/
UHZlp4Imlib4wqleshGBFRuLntHPbWZQvLJnyyu9Dh9OM+NkG5BsToofCQJO
JtXZieXotMtSBt7KL4QRaPK0q5EDm9rbdlxHJahcQAXhUWpYkYHH6m+2sDFS
X3ZMYgng7SRC2UXG1mBsmWXpftBwovXuz+9pGij1GdZoY0v6C4w7TSZ+Pr5G
JGzi+i0z1R/1BVonVo9JWzi7fFSxhxuh9t5BmMYphJW+rKVCMqS6JXY1TMZ7
E+QWrtUh2qlsfcP29X64B1AEBCtxlfbYSumFnPiq/Lua6z8DWxQour6wjBEb
FyTUwKJFbzOAIC9xwzm+wvCYn4BuSjbFIljX+aqSru2Fh92+QcE/7yAOJ3D4
d1Ovg2O1e+Tr+Y5Oc9yl+uo1yf1863QwX00C0I8k7A/ugwDLAUYyUs2juf/c
V18o+D46XcS8isxe2GOXh3njT+5kR1CB3jTYyveGdhBlP69JmTQc96yz8Glk
MGfPUzroAauRmgkDOZ2pwCQVvsQgKRwye/Q4O0EYXCi5mzUE/uPqGAlzaWNx
cI7WkpK9kbxw0gFchgC57vgkB/UXzYDS37qgYeHg0kQcV7Xubb7s8YL1DjG+
boNKejmDeFx9nMYNPto0nKEQmmBwkHs++l2xSgAt5Wzcq3bI+X6P6jxYyE3o
ML9WKDsjMsxej8BieLHNNO6ov1MlgtAetMuxlr29vfh2k8c90EsYf4MVD0OD
Cyok1odZPqhbRqkSgDOZ2mQWLa6K4hbXBhNPyS9Q3CHr9fsfBCQeJcyE3JOs
i+m1+Yeon9eGUtaaRStv8piPPG0mLsfhfcqmGMI4QlyK8HDXbs8t6AgwWmCB
4pzi+kj+BRvQTgkHTtojW+6j01+BaxvO727W9B1HsQxq8hF5lJDlH9ko8jVn
QgY2/NxMcZzWL9BJNm4D0adj/AEDE/nPvKR9fC1GL/LIicsHtu9QeK+j49eP
XBUse3w+oALkEQ6aDB47MSVJrLLFvw7qW24bOJ58+QcIzmgFiSVy3MSyIa2i
tdOFhkmXQbqpJPFuD6xuUmZrgU0G2o3rC2bzjRKZieRWPUBxlv/Gn8YVlqB7
u4Hx7BRM2lIOKoiSnhxv9x77X73mqvYsoJFRPj3wMzNif4MY+PU7q91ZujRf
ZZb2idfpHaRVrJk2/sVzvDDq82am/OWK34/GB0iJwt1m+211nc6L05LVmS3p
lomDoIgr99bZzkw41BDmJNOUsdIriFMcDfpL/HP8ohXsPWPMbEpp5POisolx
TQ2FGRq0SlP85ZjQoO/f40bshJdphPyubYv4mrxIr5UYCd8PUOY77Oq9uid+
hlFZk8jlbzaYcydQLCYe8tcznY+xZ8RjJxEHjO1kAlp6Zjwntb8/mpC8JXw4
IvCQJbpca5gxgWA5Ldv41wWuUldC3J51AdYeocvC3NtWUt1wVo6mD1+kfN2D
kLqvK83duN94yK7pxBtNYQBKv260iO2l1Auolxr23Bguhy0Yo4boEra4XIzc
i7iPUZRTxCy5ufyih+Iu5HAYGPGJrZ9IK/ycN+EunPeTje/z42a5wzyeY67p
KpqOOuDCl7mJ8HHPK9Bm+eVshrcuPOm+NFQomrErU50geBQ23PZqGviSIKyx
itk7PcVlVVXt04OJPfkdfrXbhmbSABE5gMF2SiA35bua11I00CunL4ULwiwc
3iLOc917wP1ptCAFSnEZCEL/V4pbT1+GBV1XVgskgrehsw/A1HgcMtOwYWAl
aHEn1nZsRhPEyqlfpCT7Vd8KLy7+rbaxPyW/P35IcYn3PjktvhfCBPCPeBME
kca5qY/CcAKWPkjMaWtnpOKg2kldT8zuD7X46oO270kHRsyZivGzdf1pG5M1
MAZbIznAisS+pWFm7TzVFLDaDeaNL4CazEDIN9y7w9hG1FNCvFow1jOAsjD/
8pyuHwsn/NedUz0cPCoDX4dJrf3DJQxPHUpYemDUf1sHvITGFcvpIsO1fG25
AwVie/2vLLTSXpdQMsAp0q377ioUr2tovRcnPzA3hoinOR6Vg6KNp5x4Mkx1
mjYLfOL7bQkk83sS2ldjZ7Df1upYI9udoI7FMTtPJyvHfHW3eN4XhZvVw1ck
27w3ICm+Tci63cqaEFAzMkHl2iQbq2XaZt1PB5klKP15sN/22OW0mKpHbDLU
klK1h1u9dBWfkxg8U3vNBjVNo1Rm3Isa0oim8VL/1dKRHV0AmF9yBPXSfZXP
7EZsC4V/6whPltN6JMij1TQLcFaHObhVFvzrySso3y761S/tNggJjtGvH2oN
kypAplEizkxlaAJZJqmPN7+aIofYNZFdnQbjzEZL0T/cONQYbrL+C7BVazLd
Ef3n0BMFPMpDCYi61JnHbS7rDUrVJBjPASLKoYYoeilXdci/vKEllVVZJm71
bRIqGRokQOUtjmFxNy6Fs1zzTCGuOJpzDOsgNrE9xVbe5BAu5mF0Vh1LF/cp
9OFfaSfSps0G6CH5jWvgh7crArjJ7JsWlhiCvUkvXL4w/0gOAtJPOVmnlFGq
60AFVdpJ+yZ+9K/wgl6vVMLHbpAPezU7+M4mAvv40Cx2RqLLKT9h9wWqoD+n
kawgXSce+BhvwtowhQ4NOnKEnaKKiE63j8eLubaUtgkw+hLRrO5tH5JsuBln
wVtTXLG4ppVDRFziVzHMrjLi8uIQDEVl+6wTrpVLGK9CkuWmZYC8nlsQQMmd
0DmHmFun0FTSkq3x8iX8DG0wHVUqkQS55dR2AYjQNOKKXGbU9vjyBvhYGbwO
NlS7tMl/mli3nmCUN2kTOe20zoXqTgCdtID2mhrEV2XMvJXQJMEzDbHwu2tK
bFtgMXR7fLCp2iMSMWFnYv0/x5lzyBvlEr/qakHu9prkUBTgwWDHtEK0RsqW
w1t+lXy5R9do5Hkgc6ra+09X6SYlVwvhIsvWyIXA2DwNOdDmGmeiYh0tvdzn
pYjnjOaPgurz7iyf3R7OgpnZ1ow0W4NrgblDCFR+2Ylj0HMyuuSlXj+P8c3W
1/PojFQMx42S1tdyURTHTTuqFb0jSeDrJ56CQ22EDqy3YPKxtWsxuQ3p5Fkh
vlex0R9qHzRcZo1ZJQm3tLfa2oxBHXr2dqIyGlo2LULK0bMjKU8VzPjoTSBq
0LL8LDFNyJhoT6uWPNYiM/tTQZFKrRSh53iqKTjyaSQE3hiW4Adc5KZOYW2B
DoTxDIlQ1xbRdE+bcfG99/MSDl0DNHNpG/V0XKYG6me5ajpgDEXyi03PfWO+
iSbznVB6OTKBGkiL50LhZ/yZXYgCkHJlCZEHDD/lOPUyUaFDe5k5YyxpITp9
3yRxXFI8XMW3CW1loj6VHNW4ysp1iy5N6rZvBXqXIMKAk04v9iAK97Fx3xg5
mHDKHbrqPXm0qHGUQC+eqDzFTulornp4VzKHvNXfPaHn7HICv3PVuf7TDcEq
APP+Ao3MIXtJqlJ7P+Zgt7r1LFVbYq2cO9Nvlcc6QHPtkgNfREXV3RFd6n/L
QoepQu39986gDU38LXKrZSDxkzKWNiecwFNoT6NlREWZs7TyrZFG5wcJRPK9
11X7CeOjm4nUCSVM5Z8EWepGEF2uR5roejNDwahjk8T7Q5r5xM3Nfhr8g9zZ
62Rqf5ILovtz3Cke+luHOWbmlbLhFNqRF4jYq2NPEyPm0H7/0ygUSsMrQMmA
hitWYyQhEzRVbTVzQ4ly7UPCzFRNMS3qlSXIOGPDVx1kOk6Jd0ve0r4pbjan
1JVp3ZXUVZkOYUbACEnmpn41oD8m/Sfu0IuKKHDfYXRlHBVgzptbstQphiv6
dSRsWUFmlz9mhsLNijTs/kOnrFkEFe9L1DG67TqHA1j8wQU+n/lsI8dl5Gaj
fcWCrCms/M9vQB7b+lmkWTXnjkj9Gf21w9ipMe2O4Awj2i51LGFy2y1+mHHa
NkTGdxq7QvuFvchApy6DGAZAMjIsRpC/B/eoIq8HnIXtbnDJ8UK+MewT1qR7
iqYTPRO0h4Tf643xFQagpDv3SytQPaPVmvq3IDkFCMQ0rhxGb/Vywm/NeMP+
4AxAbRiwUaZtK2SA/QT++OBMXVGrm1pFysX0ilrfZOwrR7K3AgUzllz9D5It
IRqINEU90iP1IbmgJd1z3QHFVZRXiIUQy4VTwp61xWHfuaazGIfUgZ+LNWq0
j3WO6MkyqPGBqa3Jo9GYJqSIM6yHWDVhLvz7bm2nv+oVfceWrrm8wKDfR8k5
FJSuTDKftbNlGuwrfQi9VDlqSzVbkrnjKVX9YNcRRWxMgRdwNde5KTKk6Nft
RVFPR+GFKpJkNb0Jh4irvukNFB0lvYqr5bCpXq7b9YCRI/LmQxOlf2nuC7J8
m6j+7UW49IkNLUbKogFjOmY4H8aP2jYDWqCTvLH3NDEzPy6TlSppyJTgnbLv
GouWx5ivhXf3Zhdzxbt3Zkc2wz7CXYBOZGex5u/CAiiR5iiyW1pfpM0lpdt1
Jvs/hXa9ORWWSje3DT8rwBhy1FHrhEAJjHNnc/6LrkETzmNIjSyLx8wv+klE
Lx8zWLTKS506TNYBbLdiBDwhfqAZ1K8kxJj9/kCxs3WyrHLOIizW8EHQzN8B
ypn6rzeN8meJyNccY6n3TII4DiCIuSY1rYWMykcQvqdosur3VYMt24Rtv/Wt
Tw97bMOOMUu15NbZDHBjqeHt0ffjNoSM6fPjRg+e3bnr7f6QI4UzKy6QhcH/
SnsxPN4wrSiUyFNArOTe8AmsfF/wU5O4W1zKiq9GeXEV26mND9WJNfzJ97j6
fu2oyfCwVdr8aLuME/ubjHhE/0F7vGi5ij4HinV0c3VrTuMiL+Qo1oe92PgW
CxvGRCTSr40gouxYYDyDvFST8m8jwyzYS3pcEDsGGySTaJNFtkj546sEhTjv
psKR0YGwVCJHOiiMQJp7E1VMHdrOzc2wo/SNpcMT8rYS9akmrkdH6yr8tLIf
7bOGvdtRsoq0+b4i9+zNO0xT0J3XDPFdQ3pS42V7uPXTebijAf0NY18DUhND
SQ1tBAzmKpuaH9sC1n0gr2XV3pLUtj13A0Dyy4/AW9jD0In7y3Ddvp6KPxt9
VtchIVpjimLLBO+/yr6UNzmaLEyyv42YsAVhpKI0YPcoQB7Xn88tmiWeSYJh
xEQH6yWxSMCoj6ZzzAh/j/o7cCLSl11lq7tEOR9AJAkXqiEFUEb1+FFxbtsV
i9t0jXnol6IN7t/ePsKGmt5w1yiVFSjJ0Cg8bEHqZ3CfSJ435qum3jXRMHbg
mLG5aRWML9+6kTLus2BRKC8nCjQZbCop0qO/ZO374bgo1X7EKPUPVcCCvuv8
kKfFy3WP4d5XSG1ZTxIYCOo6CQAsnv9BqyR5kyugwIx63OSABxvlzCvj/801
NW07xsSEal6aOrBabh6WJmGTsbJTKPf+ryiX8UYiXgxJXVqdgCcLwf5EoUHw
gZvRWz0k1JRJ8G24+ek8CBuwL8p9UrhHVpd/x0K9wnuiVt0LkYnICXKjzhvS
B9U9IB+Gm7hnVnYB4kZ7ztC3d0t5TitkkFBepAPtXPjgLQG8ylPaMUlzJH0M
PlqC3CoRtI9dbXG8R/qUU2+5x3dzGY/WFKVcXxT+VWcBjoZYRjk6Ve0xCffS
hEAEufmTeYIdS3ZmslPtQbPgBRHtnQtEwmDA+A5/sJTjLVDhBp2HtjqdJ/W1
7gsfF7pT4Ecm5UzHPAI427nRfzvmSFUetxLdaSQ0Z2e9mbiTCBtlPMdX4GWJ
fsF0TOybIPCmOHFu3DDaNOcauNcthyeI2O+qcT+5+iLbASKZbpmMuBgGfbjE
IQff0oPww8xMvJaOhDkPESbh8k8nTlzutEzQj4mm/WxVnSCgUBQ29372KcAV
oXafmYlpJUwxi3MLZZ4gsNNf1M14CXiNySubsoXg5Fk7JryiOwjfCdQyDvj4
J3zjrQ1VJbOUU2MkZ546ho6L1dcBNrsdPl2YJcooegZQO5pFthg/d9lOZ0HL
Y7JL3rNmzf7GsVAL2oKOfdYOUx0cOXbizCIgs4RVuUX7JGl+4bSD0nf0abb+
EQov6+QT+cgt73oTf+bqHA1FNwxPN9Ed1wGHfeN8WEDcDlC53QaWM+qSHtJZ
pOIUVXN0Oekd56cRoIcCIiLtDgpx1xoPugkLPP5QscVLZAR3E+OjkyFjzD8E
HMg7Oe81xHm2eYT6lmNMVeQYViF0rjit9GR23YhE7aUm3kVmkYWsdo6GcdDi
smsJ49ogxzeY9qhpZgcaMdaO/IUWEhehc4JCOdtHI/j9xKHsZ33Tn/VYv90j
fvDPEJoDoX6qDfQFQ/Y/dkiaE49iPncxe4VyTAK67TuMJwaHpHvMxCWqJet8
gV+peLvXfPGMrAE5z6abNppdzRWmBgAQ7KiFuIUmpWzwAT1BOT09gNFuNhZU
pR1qIfXepB+4BQ7JgclaoyHWJ0RNYjm3zNH62gerckHWbyLa5GQsUtWwkQlL
4NZx/7LtGdacxtEiwBDR+GvUbjfvU9pEP+1Hm2Qndm4zxWPPTz4jLbOdrFQS
2muYgFq4IJDQtr6kwn+oUK2rxVCfoNr3lAs/urotBlIghB/DIN3AuSdtNw/+
ebeRh7f4EqJbleR4opLhrNafrkg1wGgCQrojkb+sY1Va11nrL7TlVWutIRGx
ydhR6N8b+EFJWFPx/YaDpntLn/czQIuWlbTZwJBrNiS9gYp6ZBRoBiPpP6aY
6NfayKSMwrwt/XoSBOrMMAIO4SW5nGyDuYInng6flX/5df7nI4HOJKiiTJjS
vz3XNDKp/HCPnvJrB9Ik0zvE5YNFPUmqhGJHXC0dwIR0n9oBXfU/VkJmlVW2
Uonc/Kf2ILy6OQddZKYT6jbLts3hX8+J6U8iSDeeeYJ1pVYUnQqHcmWfMThk
XcVxSUzmRHrSN/gse39REU79RIlBL4FwiS5/bUsOraDRA7noj7RJHZwN08eF
Ih9+QL60c/ONfEAZxUgeimhqffTu1LToomlCaR7YxDzUHH1uBVnaWysHecmT
Cn24Ra1JZ5kFYEQCv1brm9Q3IGxR9GzUHjMC/ytPlLSVO4z/+mufIcFP4NNr
q1baf7GJHJRaTFpW9ZGHC+KiAv4vyqTv+7m/q1NrdlsmevUPhDwpxOqz2NFB
FVgx5sIds6MO3XgymSoTw1K6Krk9hwtR4xKFwMcN8DZ8S8EnQRGIXNoTj5x1
dWOq3/MbG+cPqqTpe++T5MwhS0wgUFUyZJLBb7Of7OjyoEuLq8K5BGQRS+Un
D4gAKyWno5j6SrkXR7+kZfTnp75AoP68AzZrIxR+yOqXXpLZtGLTCi53WQKR
q5SA0YKrTxWuMNlCR2SjNUgVlNqUBzf2LEMbA3UNdPVQvvLEOb5/e7oWz4qB
3EEAZSdQPeD9+s2G1pxSrO7AF5MWHIhk4c/IzIfgVsbddeEwdLSimTmG22+q
XAHaJLjDpxgUGgCCsf3/52w0ko4keDHnhI2UiHWiBGJdCvxjR/uvYybEh97+
TW1cHtq4wPAJmAcDQA2kAk5YKHbPfS9Q16rAWvwlno9F8DfcJ/jAW9+ETkJi
XqIcmSpbNGS1hCHwaGbADdVOO9v9DkDdurIhLigAriyAHeDZY7Cd/Md9a72/
VRlAYf55NhU2cJzBBk/Cp2P9UI0YfPlhEci57f2nTHYRoPn+AU0WcgO5e4gP
ojUPzNspiQNj0AwkJjCcKYcm8Mb/OarpP0iEMAmynzIZHISpCrZ328C2IB3f
yRUljlNe3QDCi+Jh4lt3u6nnTfz2veIXbqzRLbdvmmoFsqtuhHMnfBowaprP
0dB9Vq7/vSszA9ltEXhKThDXPINZ7CGki5GIjXaI9uJGJ4Aji7qSXpNH3MQ4
yPz4cuHhYx3mRSceBIy+5vrPre1ljVugTEuqiwiFSV70y/gsQh5MRX+eGJf0
L+JIFjuaSNpljoYxbxKft+0mzdrbd7KquNkMOYjlR5djgIHjiDqQl03wfVIv
B0p691RkVpsqcmlXefEmoLdez78DZb0eyRJfqv0hdZSs41T8bqfRDzZmB71c
E97LArykDxSCszRD4UBuWCqP6nC0YHekROLMkVUKK8orrIbD2iJIO946JJDD
ilqpmEMLmQG+4/TTM21e4kZNXoMc61tKXLqdAMhcnFiU83Mn1snFJGcqZdou
uVtnISSZeVR/OHpiP64Wh7jZx76//cecSMxu1yyfHCzZ8vX1YnIlXbrcejhP
izj4RxiqMnX0RJ8kbCxawZeOMVM1iCscOR1IFiO03oY1V22fir2Fksx8wTdp
JQOJN3LdOt0Gl0LcWSF1bme0gWNsGVCUCCYmBkYz9GJvKRmTERF6foQi1Vwy
Z0liS1S2ipeBC0xiulKypZJus3rBd4/fvDa9XmIYmM5hnsbIfa60GBoarfLk
FE7mY6xsMortWkLQyfDK/r0U6+grMdKKbIlqnX6rY+nShAt1YJCu19fnCexl
NyO8BaE7JqzBiEHBDl8Trw6Hk2hVK+LITeF7agvQyGvtuJ9Lgb9Q3vphiiX6
rZ5QJDAjvKnovQMAIZk5aInUC2GnVRgIWhDCPS61NI/YsPTYckek1oMMbmiz
867aRgyeE1KQnjPvvP/G+bMXsNIAzNktg4ZatedZk9jshkzvs4yqUmcUbq4H
ht1y1avAQOW2G9O4Yjnk9ZOyuPOAFWgVuk2aI0NDId9A3clB4Fa0lYDgXEHA
EbWInBbm1j7ZDEetHYU7Co2al5uVg1leFoPHZX7Iv6maqK1n6SufJAV8/01n
FDVFbPV118lskD4zM5V7YQzlrEnWZfWmZWLAyKI9srj4+eGvIWboV833O210
tpYOfxKySwUUug3xv0YgCznPExk+WkG096i9xD5XD/jytxLIKR8v5UEl8ucz
Z4X+Q1lEAN4mMxpx3YDgPFC0tTL8cVckT3GM7Jw6X2eypNsmXJAamGwR3kHD
u/Y6M+/VezPx0h0WiH73bxnSeYnFZ7cVQcSiXrq/1SxWo7QAootI96Ah7k9v
1izACHLKBCeYs5QfqaaTrjKnRP2wiUmMmbMOsjsPyOAMU6toFJgss0GDqNlo
b8b7ZT+RiJWlwBq1Avy4u0x4/yAMmi1omqsGrbCcbFbjWyoTEantr7aaZzJU
XMFvqc9dokSG1qG/vpDSH+BrnL7kaSiu4GkS4E6j1Mylx4zltMZr2C7Z7A2m
7Dcf2KA+4ErPSmD429dxswY3UdTmHoe7N/ETNJFzKqMI3LDzcut6Mi2mg7DC
jUo4ZIZZ12uP4rd8CbYtFzMsQva77Q2s33bjNuQKuXH91gYplX1bGczK4n7b
LxNVNf77e/K8H4BdOVyRvxi3cJ4MtJolWjBxqRB8Wa7WsdvAI45iZG/RDstB
VZlmo5FOSq747jcBVLvG0yLDvUJtK7CkXdmuibgcr/ynh/YI3y7lIESL3nU+
GC3h1vZuf+Saev8oonrTLxX2CL+ZJhtOLYVrdKQFfd9Fxfjt421yxUuZY1Ow
2E+V/oZtbGeRAz6GsDbjXYEL+PU94/C+QM1WRD+8/vIEdYb3suBp4SODeXKw
LmVWxPtRxERIOtV5mDQ0+HbG2RnLDJZHB17yKWCuWkpiU9rHXe98opOYJ3p6
dduJQvixDQNgwbVbvKNHpYcmxkx/ztlj2smQ06x5IoyS+hbstJN2XSHjQWGV
MHDrp+9sxjgaKYsvrcHOSsG46XoM2P2eKD+1Rh4YrvxqBZNwGnUUdTN4JF6q
NaGobuI+2jdGvHItj7DMvOj6TMM6+YhphNJJPuAgKyt2JeN6Ne82D3a/v1s5
Kd9Dq9eec/2XdQ9mj6JWETQl3MUAo3XCRXxWTxkV5dxOxNTZBAYHYADC0Ou3
0XeXovf2x/yGbDEEcaUFDavEZVCZ7HhIbWbGk6bHqDqBN0ZRzZmLc+uW+o+q
fAKWzDAfOjOCA6QgJH5f6eEe+e+e7NGvGVM2mL4+7BmoeS9J79w+KMaJpzvY
eh/7VjnLe9p1Pd1HNS6pmiNnQcSGgMQhnksP3XCKeBxfDD2H0YpzG6g+4njT
tpcE/4czcsHsJcFtTYKxTr5vZn/XhdVTqYFdrWgTY1C75i8pE6TV5YpNfMoB
1gUtwTPoQROgdbVu34MNu+nvY9Xyv5yo8Lw08/+z3GfTQc8Z4eBmGNNir2tj
CXTrBijFJMXfGD94AufzCHd1VQdjQbEgSqULNYrERy6sSxPCBCsNbir0aIsl
IcUbimfe7CPaKn6J4DTDufsDIPoaj4WJVbKaIMPmRZwGJp/D95P7pg2eX+In
xLJ8awbL0sKT2A/Jerz/Yx5oSR6WMLB34Nypf30iJvQXRS0doUgYLZByHcC7
TsHj0sKYok2/fgWefYyTDz4xFAiulZsHOmuTuQZatKTON/+MxKsDTWj0RCny
kBKJHmWe1wcHbVR5OrN1//joa//VS4wL67KimsgOYozle0UKG6Mf98ijVSLv
4CQHR+A3hBMb8hTrpJm0yOS0536B/0DJfybDVNnY3SPEzA4nHR7fg7BATyGp
oLl1rXT9+sTr6AWSEDo2CyPDi4AmMfjbH8we995KLZjk9+vWQrDBvMnTjSwE
/SPTXWzYDD/zeH3i+8J8NSHDmnthEsxQuLgekLX2xDhQxRr4oX/H7iqG/asc
7xULYejCuMgqykyw2wb0+gGY17QLKQ73IkHPFpsLHtPeqjL3CobfCHo0HES3
T/hL9EBSZzdP9n0uH5auiGOCvBbc7KXtT8QF8KUWGxnfqbt8hotKZlns0eLH
bK/xHckVFLIIkIOu240MSbvCK6bKASujdAdJ+GNFy/M3AUfnhkDHtxeDcS5V
kWZhI/ayBBJUsgY0xcmmtUme76mZwLZNFLV0MY7PbshbT3Pw9HWnNw9tx86X
yY2kQ7IFkHy6DLgxLLBD5t7opwSA3B63JkJaG5WTv8VCvYampjr2m38w8Buj
/8yMz5n5rXnKfq5SNohBnw2CP8fCylrp9BnFwOaN5sJS4ZjuZ/z4EEmeBPyY
QOqZs75zQwFVNK0OgZ0O+AIqj3l92G2HP3AWStqjhScPt2efEbbcnXs17xyq
3bVZUTPxF06O1yjZN6W1VppbarP3PsLjzICkab2j4geB8N0x+VmdPZgQsp0n
HWQWZncSJVFZaBh5gc1T+Y/wYSOEYYoBrSo5fqAQRySca/tiFJvXmkWPa1iH
o7yyRebgZ9CT2T4FEpM8nu+vqeF/1n5d5YKQgAXzDGwm0Ke7um4rbsTQITWd
PydhpyuYf7o8ylaAcEzIhlWDnIOx4VBY0BDLwPgyXItiFGJ2oPu4QqP3YEx3
klsSWRcwatMfvak89ZUGChhvi0IK+S3UOr0vuxHDCb3sfwLndbeFiDWEeYV1
D89D6foFv/4zo4Ka600DAhAovU2VMRmhDtrhZq1zNS7PWHnKvWiBRorCy89+
rs0WjyMOiAUKfBZs5hw56nNATY/p2ZJXww2ghfSW6ihjPIBOTf89EcNAL98m
ovS306UPru3QwV+psHp6+PYvg6vCkTgToo+0tWciLqNJM7TsWYw8f6q8beye
ZMzR4vBkONWTLlUHK20/w2xA+VGvU4xROPMmmMsM8ZBRgUz7RRZSde9vDQK8
GayIJPhArFN3y+1mmp7BpVKV7tI8fX7VkZLenvWgl6IvTHqm6/jfcHWrB5Hg
WI99qeWNZ3rdftUIUJDxJNASttkQpQJTD1pYTelVPYp1Pn/rIo51sFQow6kj
C4xBCRVxb7yo5PcpUFLlNwyCk9onbO/eJGaFyAOQ2I+HgF2iLnOWOtW/8d2Q
eOrRZXfcNsu+StWZBEimFpS0+rrLJEcXhZIPjIBnktFYxn3/u8pigdf4tK+F
fXIwgvAa1xdrqtZdi9pXlPq6RJ5J1BCgRZaTfoirg2ZkdsXBIw8sri9CyOFF
jDiSGnMpd+t7r53l/DHuhSVcOMxBbI3szRyB8butPiipj2nI8eRs5tL4WmMp
2Cd26ZgckMOHT8T+hEKiPsKVj6vXJ3WZaTKj/bGTLNQKM+p1x3WXV/hrKyME
qvNX9EpHfhdGSdqJBlzQxmM8FnIlyZp4aVdRu2/a73Mo8frdkku4AG0fgWtu
DwCCGOPIK572qDrwABa3nxdn2UqNBvlU9A/4RqBQ2EZP2TJS9kWoaNlD2Q0f
rx8aixPUxq8m+3H9AymBXlV/QMRCd38X7frZpGDKgwatN13aylKiD39opHk1
1cE1KNhBydzGT/Jkm0/REVzUkz3l+/Pjn+DVepI0EBA+lvbiIzHAYn0jkCQv
3yJ6lRLOJ/quaAx2g8lPLb0heiCfpc0gy2MWULcq4zAG4TT/1FFFlWZvDhvv
MXnkiQmtVS6MYSSizrWg4mZM6GhQRDndPWtxqVrmiWskt0duS0QfxBuatsar
qhR/NZKtqkoJyz85KEPg5fRiGSstglwpfjG/4wTHJtSh8cgMGjEGcvtXOYEZ
2VuSzIvJOkRuO5bYNkpAd/pXXWwGfmyueo8jCa0hwaBNgT4R/EZXgoNW+iDM
5B0LewbO9W2VI4i/OPrmASJGKNGPQv7FOK/lZqPJg+jqP0wFdSfoatfEucnG
5XiDQeqv524i/5z+c0dRBMoPs8r9YqMNC4ne8ajlA70D8mxq16RtTIgDiYo1
SEbqvFSzqul8a9ny1B+sEraG+OxtoOkdgdwAxvoRPpO37gL9DBzLWqXyz/RT
7ubOc0xTIyywbFr2dEdXVSK/gZLVyxOSN1pmQ9lCmDk4oBXMRQqnG+hQ4CGP
CF+WayvuP2xhg7pI7fKuxVNiJqnJomt+RrxKFN0yyLFvqO47QYVkNwq2M51y
k6mur+5sp0Vy2o9cxrVv5ASoCyXN4GAaumEF9QygTmjy82qzkwGI9wA4OMre
0B/FkeMUK7HmyI/k9OU7oXcQ6amaGKzGzfjOCIIuGKczUwujbNWJKv9/Wjo7
67QT1zJiQgGP6ATsVOnLBtYxlZ8JlnCwlfal9EbVbFNhIrIM5mAW+sRSfG3y
cnwA2CO6YrPZh7XoNaZ856aKIJheaxvWuPbeN12cMbgBNljRrH6Op4xBw7p5
o+1IoTJhfw9iruX1dL/T5jyhWpMuHI7eJkCcAZ1AoSP+Bri6aZafXShmvShU
NR5qGkaaN5vFvgvseFVHoN3OGOSTOWWmyW5FaFphVUYTL6k8y5+lEQMfVAXV
3TgDXie/Uh3urtCn0NUeUyKM1DBlSEJxlg5fgupz42gPDkh2pzCOlEB26Q2Q
EaoS/ONN0BtmMEgxTOZIjAknQD5xVkJHOtqV/xAyhG0AczqlCaRKVY9w/6wB
vtb3oKlYwolZmfD5tr3vNc8XJBFfH16/YSb5pm7h+VOVwHbsnxGGeYhl/FcB
UmNHL/kb3qvUiAop4UMMHGTuHr++4yPcqZaDq/VZa6jYlyYyq2N5yLGFbkT3
2sYEzSvWOUGq0UxBybxMg4rGd2EhiUoCVEgmLvbG1bF46pdkAfToNJXMNQFJ
asruXtIDAPCnweker1lqs6va27aZcWTcnuSDK46iaB3AEf9OsoCI1hzafTEC
Iw/Yg3LS/AJMpwz38h3sfYYipIA9hXNkuU7CntyCET916Hns/DrNx4c/zq+r
60s/ReZchlgUOaYxZNfO9lhQV6lqBPmGhrfkewE8+tRMOXYrwIysrOh4h6CT
L9G3KcVuJtPCNToDxw4JwDW/HBuw/ajbzewIAjvXYicEnD+62EzvP8treNDs
CzwzsW3jexEolkStsnDeko5/r5HDrZBNzhtQK8ishc1IANmL/8j99Ht/KfGO
36SqO5tvUM/YGJsEdQEbMnZr/QHAKyTS5Yr0diiYfxeMYfB1nmgLhuv4BmcD
B0em79EKE8QgKRDmOnvJUyPr+KNGaCVCOkBY05HzLXhPQSUuqSU9++NHOcsK
xP12rl/IXgZh6yd5+KfQf0IZnufy4S7Mql7u942I8UsPodm4V/u+PFmM6HRS
QZ86oaLc1YjxOUKjr8Bwg9xe+uPm88xrxQUlBBbbdXpMaEEFoJgIXtjUPWYO
bSYzV74AZ09JMbmAphOW/A19hCU37yy1Gs+rn41T79kQO5+uxgMJjc9zjLMz
wKVHWV3fFTUFa7QV7ofQbN1lVx8G1x3pnB8SI5CRCDANvjKWwLtUi0RV7/yq
wvSkLM8g7caEFusS/XEehgsIj2PAXmhOckRbGbpFZ57+jJerMrp13YYO+UM5
+SuUvwm+3Sw0EjkrIF/6xee4LPUdwKcanMptcpIFGnJoDka/wXf7nabt/1Dc
fytw02z4mWuKtYtC4yQPvrBy8vT5rbSa8+B8EmmREKPM32treBLAGyZPKtcm
su08bF44xrUzc/r7hTiRWnNCdggPEV0KFxNFSc0/wxgCvSNpXGnO8uWqtGrd
UrVI+jtUJ7PXF2cNqwakyo6BuofahKb7BeMmiZMu5V739/pgiWo0T8IqXOLz
zhwQyEgNVJz6YR19PE0J7bEjUcYCu+XWstA8iI/lWoDG3O/MfvHlg2bhMV70
nMMZhfHYLe8m3DOl/j0f6gs+86eXSqWBVa+QbxwmiAsW6ChLI9jQR0qzqEcm
31A340wGOVxJGDF3P9sEkWxis519VJ96sjs5XzANfQZaF5LYinzTxH9HU3gs
IinikYrk5svS/bqxLV6mW4Aavad8A7cBXvGqJ7aRjfmQy7CD5ixuZtd0xRI3
nAgrfEhSqltwg/TmjGwami986esIbhMpi2ERb5izZUzZYDqYgLSJvio0q5cP
R9/sgZbiD/CASENpgrlhmE9t4/5iL2KNRrVfcETr6rp1u3ow8qM4cVHSAAZO
NyGG7BiHl7/gDFveBZ+h32mQVu3ddv9HoCpQcNz7mdEWCDsUPFg6IeNB4M2u
R+ZK4o/tijZ3szkXw9LfzABuNKOEGKFQ1/5MAILVBd9swuoJB2iBqt5NKPjk
T3FqL3my8ylFsDGIU3hR8C7/w8Ow2WiRj8n/FIlV5VpbJBxOjvOaIpYn7Upf
no+8NBXqmXfueIi1FccVmMIpBFFmZ/f7sEO/n4i8vnoOGRYjf3S7bNX7ODHW
ed4oF14ox8ACE8NnjianpdgEUYjtOIQRklE2m49iTe8QX6Tq8Y+F+ZnlzFs0
gHVQYq5QmgdFu+iNua9vFaJZoXxuoB9hTGObF0ucXucaGt8VI8bvPmPSGUEZ
r/HYOKXhZ+Y98r0SVIvFVRjeHs0+NMDmxxfajWiyf8lo+I5AlALb8lTizGa7
nKIa1iDyOEVN+zCUyvT5FudqRoq7AT/LGB48iPTK3mP+TkjeJBixobhRFZL8
5bQD4MgufqhSfJkrHu+3UBhf+D+0goRx+gES6t+6I/3x8RRX3eddawPjwUN2
es8Td+pUoMBM1QWK2WgZhR3mFybLz+HE29St5fEIJw6XyjlCxB1lUm3P2zNZ
kViodJ0LyjSKhT1uLg97sTMsVUhHJUitWOpDFVCSDPO0zgGn0MZLK4011Ptx
gjafxFL4xXBpwEgn0Sm0LZwUL/wuM27/nRMabOOEzm51cCaKbsVgd/sk49Cv
ZIZPsTAlPe+liAgD0yOIegQyzNgwx6zuB6cNpWi3dVdATMYUb+WKhemzazA0
IGdC+5QWbfsIyc4Lw6kp6oAaD0DHWQsyfApxJRdmQRqK54wJiM54ulXpKPPm
CsiW57+FzLrAYSGIVaRDgm9ZWGoLhG9eyoMdnyshbXjMbydk+6GsHqtlhVEi
6zkWEwP47s0AhgIdnNjoFJhJsHetNtvRgTbfQ0ltayink2AWJdKc77I0D878
fCYW13tBAhS4fFY51nx5d8B+6u3bdc6y5aEFF8xhZCMEyfZ390Z/Tb1cNdrc
ZjbNjAAED33wz4AvJZsCw2PSfOOGcw1vJ2JqrmertSgN1+jJDKbMFuJna+BD
dNwMg4apHTWLqU/KX/tymPZ3NlErYOQ6F+QJZFdLTd2QDQzQRFWfDDDS2+zt
PA8khcsXONzrp3XhmHOEcMkL9WF5z3awzDVSlmimvoEkppGQl4Kxx3hb6xrs
4Yn4PAMj6Fy6JObFCWQu1WGc4gCiZmBafR6xwrcQCXeocn3rmJcI8IRIl/Qr
0jGvrL45ckUGXQ4YAF13bk1GoERnXxbPNiZn3yES/ZnjuRxoS+KbieP8iu5w
shEDrfzhKNh0/Wg/6vk7MgyQ/KSh3QV/XaZdst8gH4pvbDVfKud2vThgBnmH
ymKuMK0LFIX5xOV/9u9I0BU/lqkT0AYn+w5IchsQJzF9q6YlLNCVsCK6exxd
hckrycPxXTSnxXLUGn+uZUDmCVP+SKA1QlQfPJe4bNlJmjcsJ+3c33syyf1J
4eoacqPDxwaaFbnEFTjFRe+9iG3rm38tfEDiNt/y+23vsEvwjB9v4bIUuFvq
f0irwmeG5feC5CCq1cKQbMzoUqMEeqBaj1vA6273IMUli48fPrxq0z/9zcyP
bi9qqRqMSAv2nEl/Dua01tLlsaPpBmOQoGKBp1qXYb4YLdMttMQbfMxYjdDX
QJquZ6Dz0fPBz0riYfsrHP2nWVwpS1kQ2WMfPDuxMrxIRLmyP9ejWcClWNOD
6ImOgkc4bw9doK9UC+FPxm6/v5G3D/7DIfjVflH3WxMNu9K7tMADsXqRyP6Y
Ity/9doxZfYAKVoi2Yr5wy6Y3CYSVV2sxees7XLtkHFOUaTJKVmIy6xjodXF
avLTktcj+j+5n5zjq6+YCwK8V8m4irT7gEP4NXSwuy+CMCUUFnz/72hjo2C5
zH+XZHWyp5SmJG60V32EIIg+GgM0V08dbYIvp/4eoF5WvGifwCIJNEBDgKnc
VsHICRlJJOzsGcmFfjuSCFP/W0yU0AkoCjMGDUXSCLxqZccGNdfRB/RuA8H/
mkIpyT22Dq0XGJY+B7b7mgoXYbH5ojPMLmIqu0aBvmMKd+YpVjdhL7ixYLkg
pKleCse/3XzglJ8NEtBw+lnlmn7SxP64+a/dXMyEUpEEZ8kWiRvZMdm3uWdq
ryklbJEOwcvVpBAWoypPG1qtG2dS8kgk7If2IrAfjwfZA1/icuXEX+Yxc5Iy
apfaxobI8wrdNz7FsenRK8FIYyMKjYNDODRcfo6zHGwK26eVJfp1COp6n0Tc
4b3NmFR1VPKXCZadQFkLTaQn67tKn6sFV78ziz0Pyt0XZxGcZusr84Pzpc2j
9VpUfCPmmYyEeG2QMFQoFkaIHOrh1EHrVqxiEqrUzqqP5Tr2gewk6+3EQTJa
83thqgJb1TtBgrswaZptZJbq3ncwxZC8irKp19qsunORtE/4XvLcmOby5zVC
W0DJn1CSDvMuECGM0xAzUQj0DePJ6IBqRv4YPg1xUp6/71dvh9Orha8R9VpL
h6DCqO17iYM3yWTy7w15+OQZwDL7uOxgA6HZvm9pKODbJjh46RChgtBKA//5
KgOLmn2FG1bnK3mIJkZxB0v3ISFJzH7/Fcb2LEzFWHdSAdl8/cNyg/UsC06m
2tu5GC9dhXckz94Yl4FAwbwcu9+LnMjxVRTrp/B5iEkBAVfgvW4BtURnysnV
PMEaMgbvMau5KiaHIGQzpmGPed9FcudqAksFqw4D8uqBP7FRAIy/yFoCp07N
Bej9AgeUPtC7W0byjpllYM6m/+G0/+TJybrd2z2A3gnj32+FvJYC1AgFfcte
yuijPvV8ApHRpWukwC4oSfGVrdxGtBwI4JVLuSz0+iDVhDumAhNu+ha8lCss
VcIwcCn6u1mkYKMl1ebF1mARVNjCOUUMZqQtD/wlUc3N03T5KaH/BG+Y+K8W
+RypWfpBXJUsbu1SSgOm/fnSJECxko5nCOfVkeylglUbe2RnUyhrA8yweBBK
SEhXRxMGrg29d96yh/qIP3Byc6psRs6771I6wA7jAWictr2KUNvPA6W7w19V
Q89KMqpAx1iYG5EHuUZ3DFh0lOnqOFlAnjmdSXn22+WcDhdYyC9ja69LUDjV
b1KfzMgPtXIPog7dspiaeEC1KncL62i7CbElfTgo6olKHKNKsVmoQgbeAuBb
Afo9jARJATPKEEC/cuq51wYd7HadQ111DoBX0lGahp5xrHDZzVN/bKSS6t3S
GGXK7EFSdQSsCDythpecWMfYUaeBxLYl+BApqH7RuA80Yo3yzEN6/bgx+Se+
oNkO2oLBCcT7pcDfDZ3BUgHfRGomTxI9i1Rcico+zD/gfolDzzG20clckJ48
WyZrk3eHWrpMFCmnW7IKJN+7skWdR/UVhKnRF8v4Ovf0E8Igdu2kH2mbeI80
4B1bx1qHCEHKfOaEl4RM7pFmDEHd2lYEgUu06CblCxOx1D2z6zlb/HLkhxG+
kQqMru5uO4ZxUsWGY9WKagO7zet4oX0rUM06inBjVgWLKhZt4CIoSW4WlcTj
yvB0V/par4q7i/ayqDoLOsPjWP/MCvO1Yz5pxB/7na4XTwZu0LjXC6GJiPOn
gcmccRTLNor4+C/HEFjBnMftKppKMMxMDdCkk/oTKfOw/pxK9iRMPaAkACwo
wda2T1Lf3ot7Yu5iqCSNNGzE9aADZvmJKcfSGrJtiRTk3voTJxpPgfC2i33G
2Rz9siEDzID4W/vp8OzpU8ZiLeWg6W2944fyNp4WXkA4ea1eGThw4c1v8MGV
YHiaOMZbIB5ZjmNB2fhC2CofVutN1yoVmTXVFKntWvvgwdxtw+KfYFk2nat1
tDqXDTZyUwX4P1JBmF8mC+REmdkLibhyKw1weaIdZa61lnZau/MavPfC7Ui1
zPoEq7QURQJzb3vg9L5G/6STbaK0+meH5ELuAapdU6hFbxyShF3yF7CTPCZC
hVNPanIrE8oyNI1D4JBIA0to04SwjM5uSq/ZvPjzQd8yRg6WbgPQmrAZzKdS
mO9xKG6oDKE+8ZrTbGKfGatavkBbUT6NpbuEezovgBfBkE5QRJ9lav9mjr7T
rsXH3GMMXBUozVt4n5ufd8POXVxqCML2HWyHr8FgT+hAgi7gAjZI57Y7779p
fFWQTpm+8H6CYslSBiZi9UTFN1OyZPb9BIxd7AsP5zBseFFUGgFklIziguQI
MjTMVwN907SPAHbfniOh99mJM26x7OixMJzjwzjna6jm/zu5yFE8fRQBh/ad
4qSsQvL2iLyrI73ejSzZDBkRBQu0t/hNkCy6hIBolh88JMH+4etaCdTCWwJZ
NxDJ/FRlLgMNmgkYmGPVkUxy4REnfd8kHrmkx0wBXh5R/Y334kp9Fx5X3Bq/
CmFf6WTNtTf5KzHjIw9i5KskrkiiWsoqjbJE64LmAFOKAfO0MjskBsK47hFA
cNd/8gpTIhaP6VJ6KnmJTl8uPJtjqo5QXq1hmnREvv6t8uztCnznwN5JdNoR
hy7gs4PTdQpy1UPWp0Hs9HZcWHDxc8IWjp8U9RE8EhGSaBqjrj7nc6d+oRZx
+FpNksKOUwHuY2r8oLTXCJ1XAAdSqWTFN4gL8MRKjXNIxoBbH6Zo9cCQLwC/
xcTpC4IFE7dGtDphnf6UmdRFz+6l/8sgVbbwt255PwWIqy7XmFO9RMSI0CB3
49O8aN1y/jHbTjWC3jnjtKbtpqnaL2xzmcphJs8M34kWC7EgsE0ZWKcL1mG0
K382n99fOJ5YoUcIdsa5yr/Vzg0O3mp8ARYY0rD89AYZT7MSDn62UQnrxjiw
NqsxViH+Tij6hp6uTDfID8dP28e2aLEgOegEzUyRIY2gQKNRa7z0VHlygXnS
8h9k81/GcqdkBZMc6fivHeFR68e09okh9Im8u+E3VmQKBoukal6o7eXWJnP5
ZJiAxavVRP3fHnCeWfzhQaXqES0wvixooum8/cdfjvk3v7GlCwyIXsPXY2c0
VkLrupBQJab3MqyxstjNc+M2rQ/z9Wo1Ujz3CNp60nfjeXqfU8/pbGqjdSeh
3hWTNT6Fk59l1cCnYqxYUI2BgApclYI28jNZSlPGD40Tbv3Vak2kU9v326x2
Fw8sOCB0eKgKXlVdzQ8UEJ8uVVP3xWhTveR7B0xr8gRo7ZxkyeeK8jpA+lC1
UXkFzvMXwPeHwmaDCzdwdvtzvQJ4POLtuAy5lLC1fN2ZP2SKeqwU2RB7rchC
zcFXXlpoXQ6sYL3A8v+bpD0HmAtQRDIgNhFYayteui9hDYE70auLzdxzSSlS
DtLdS3zyowqznCJH52qCCl6WkY5HuBz+GHUvXzcxF8epqOI6tYEMsydanzcW
q7rczeYKNkj7LVgIvJVJsLZkXrn0JnMijPc83pJJI3Qa2NOTS1dMB1/B7iA9
rTHjumnFFNAiouE75S/XdEdLUWYmKMorAEj6rcilseJ5bKRe87UYwuWTpZG+
dxrEjQZVKYvY3yQf5oWTzwFfdTgbC+txD0jnk2PplyXAe+soZcyc8/ShuHtf
ijuf6NXFpl6cOXyAotrDh2nNaFBiy5cZEKATz2JjyUx18Z5OekXJ6AZdc3tO
kLU0ehUOtBdIgDby8mJ+oQLttQHdMFvugCMwf0+Zi0m+UuqJOHoRfg6VKRay
qkFiWo/mdynzZ/5Cm/yBnf6wR2LHjnQjqlyz8rfCuF/+as79c+2/vSnLPxYe
l97KXTMcd5GUsyQ0bqG+NKzIme2gObCNkT3UI0nWwZgzvJWqMBmtjX42C4yJ
Tv8rVoSkLBIhUGrcRpxd5R2hVz2SHL3s/s4KDH1M0D8qz0l+/LFEaN0TIptO
7SCFM7kGx4VzRUY5F5ARIUDG6Zopc1xZg042qSRqE5oYkNuNUNSyx+hwY18n
wdwu5M602eYy5gPlfss1euDG6QfkbO0TFgnZBBVLcZhoBRQRDd8UFxbyjWI5
IFp2Typ02xC9wNCA9Hqtf3NUlAmFULnlQe96WnsAIxjT6pub8PzTNMmBH1xT
RMGHR1jwRbU2l3FOGSAzWNf/evIDAMhiT7WMVPUUGkcnY2BzwljZRTImpDFW
HFD/VGJWqJSFC/pkN4XcE/31ky97erU/oLMEk/+5GGFoflQC7jfbCvN4EGsu
VvxbMaU0fF3TuOi94GSUwR5H/JPm3Q6GNeW3cMw2kar0ntOH4jEnifgtRMnd
lNFsjbkCMfCxPWilNe4uxMYNkMGDjJMVM9rBQ9ZOf84uqFRn4H6yc7aWVNdZ
OHZq8EorP+vXAv9YxsfBTqJb0BZwa1YJxfFXBTB4d6eFGY/GkEVlJA688fwc
lKTGOXXY9ZraBc4gDm3lhd1npMKUfAnjAC9O2P/AT5yXaIa8/yRi/GOH7JUS
OcEmVukdC8dJhwdOg672ipXhSTu+04tCUrS0NJbFlXSR2gWM/5DX92qIesUL
1pkje6V1DTY7Eow+GVMPE8W1dBV3Z8d53GTAATJX37OhD7nkdSZyvFbvyTo6
yDUY8csyKA/xBMlGSrsLYsribCMObcSzlDNqie1t9BdDhSqQp8Yvacc653dc
q+gY2bluPWAFVk795qtqpn/02Z/OwWZGsU1uF3If2Fm0b26+YD/ewinsOBQf
SQupAg3Z7h2QomckvOaMYPV+Sm003bjarOkqdt5S44Lr8dU0VKo9ZysrQ5LD
EHhpn1yGOSc2USF0N3+rCbNRlYeqSgETZpM7xTXCTeG1FJqkRtzygdy1JDte
mLMTnrrfW/gzoGVhewX3q68rDnzDJx1E3WwP6U1iJU6fCP0MIzDPXEYv4Ad+
SdnoAoTdHd9OEyUsjzq22qrFL7I3Bbq3qiTQZK1946xOf2Ru8QDmz7dalo7D
XAUDqyKmwi8ExvHh9MLQRmFqqdJM8Ue9L4AkoiB0kPmHv1VSI934aoobmVJl
b1ulNxrl8y2w8HUdxohfHILYjyAmj/tmnKQrMljpnht5jXR4NiHj9eVE1CXa
y99MJ5bHlZLClckWkT4HBC1SUj3a0JIFMCu+icB3eidE05BKibWRpsCmucTu
3CXWuzsEAMZgjgsHc6/RI9iJL7VqpQLV2aAuwd+D35tgIO+ghy4zxzux6Ek7
Ka0H0picB++TixNL3Ipdx2ynxLn3IFej2TbXl1wWBSOtXgfjMMuu49WR+cNE
QfNctEDfPvXIbzpZhLYR3q+j1k8nn72+K6+iMUYr4f+5+jdYZyXJ3vh8pI2U
IjYLvIqqbAccT9cGLUlclJJEGqF+3MXdHm1rc4X9FjA4migR6EyTSRazpG3U
MDENwhtmqVp46blGVqxzQ9eFkK5f9MZDqD6swOeojkMPpQ1gWtr/p9v9JhuS
jbXVzFOIIy7oO9wDmP7cyuYFUymXizZdTnrJ14WQxv7s0Kp4wJtsGtb9mGWL
HaHXAj33OEBjXBmamqNINru1zOl9Y1Q5jpQp/3t+guxhGFBgGIKfKVFVXY+g
uRG6CDilP8qprLfiBVg+9iU8hrUHvnUdxqVycDkUIsrLAI4EbZeEjNmtUBW2
wPNL96w4ZfADl6BSaF9O2I4gDXogXva6ASkRYhmq1pNhkFT9XwzIPUqS3Gli
e74WAz2str+QCQUvbXVaY1bW9dv7lEiZQkc5F4JmTXlagz/2yfATBfX4L3UA
qTQiiwzfPnTxlae5y6uM+OQg6OJu3z+PvP0/t6SGG6QJvyxSpjg0X1sgM5xn
N/6mVzBgs8jWMZGZIsaf05ydhRnIh5NSTRtt8tYLW9yim2Pq/Nd2EE4Q2IyH
pVMLRoBQMwTCEKzrrgk8OTq4AqhhTp2XtY1torLMt/2PFubGkarbK8AlmD33
3vsu73uGZHkNZSGKiia6D+BG9zky4nbnosjbrttMbHvoMeoSiz9JyWGx9hKA
vvFYfp72wQR7Np81+tMo/JEW9QG8lR1x0boBXSy7Uu3OFTdyYdMtHM+6GMtw
mULqU4xHJo9a5dpaYPphsyJPnKM0KZdwhOaAqZU3fREOsH8dzEbacSgnMcGD
dS0fTnRpgdh8/5bK5Xw6JhXUOaFrNNilvGxUr4dbKOKDtto5tITL3aYo702s
UIq+8HXbS2CqCXq1X/9k5IV7MiDVEZb6trXGa3ZVGIX3mwCqg0rg//6JQ0b8
TmVcmMNqrWnUpr+GxtS1C09iwoG3as8RvitRg8AqnBKll397RyK7zWJ4rfb/
3C3lUfqP+OzfRMw5CCo3Ud0neSCs9dbXbH9HZ6LKduQNS0OKjT19CeIZ8aOl
hEr0GYUl3qPyPzaNh9M8SjUizFWUh72NtY6Vu+asQGGblktyM4pig/ISRyxH
MrhV2M5IXnRUwFnfMk8/pxvcz3f9bIwzR/iPThIWbveGSxzh+aJH4Qi4Z3ln
fOhmtri86jT4PNyLlubqXixo3qnxHiTvAQiuplhYLCS4vrLNg/yr2/+K1f7F
H5p8l7wHyC3YG8T5ribza1Eght6o3j5YG2cPyEb24O0hecUN/63RFaoR87Jm
h7IMcJicoau9HrF4XZIVhA8ngj24ee/uQsSNmeO03Wm1BTOQ1w/QCpv4ojQz
vlji4DCPxnG464k2Cpprzo96ojbxsiX5Bz7G9M//TNnTLzh6U1P3cMcMcGP/
dN9xhnCjLQx8HBjBGwBYLu8kpcfYzlvdwp0Fq6q+O3lgpPfY8X+82DnbNwyC
faT+qu2h4+O2FxQuPiO3PuFmQvhzWDKx+o/x2/l+RYYxdlfnPj/iFITtAmFi
0sb5XB/xJILJPBUN9d168gusAKdEYuVTV99YqZ0k92WWZ2sP/pKdfC+5bC7b
LS0Mszw+gELAwa6OvFGaaxF6SsthZ9Acud7zNRJ1149bOeaPSMyX63X9pubP
KioScxh3RY2X2PLL5v05lPsuRmz7ECz7m3z9KmzhhjxbIXxynOrVpBtGMnqG
OudwhGSHbeFebU453jt4WSP/mxvFxso8Hen0geVTxzlzeuB1AbjZMwE61aom
o871EltswbVpXPdYp/2UqrMOR8boNvudziFWLMidusS5DqTH5rMG1mq3MN4V
lRX4PziFxeH4HBHhwGr+66klmKg0MHlV8NIqQXFLKdoOHMmck6b1ef8xbKYT
abLf3pAAqYShGDLJqnTaSfQD3xHasoxyX5Z/OHM4dEAdy+0XXcfjRE2LdgMu
rpuHfkpwTB3iYlvtTrZ1X9ZK+/CfjNjbaixEGr7aquN5jyRBh6lHFCX9Q1SV
c/Q6hz5/gxCAdEmt0QjP5nAAINZeXjrP3kg6JXH4RcMAemI+1AxDvN4g9AdO
12REthuBw/DNJrtlq1nJFM8JE17PzF9w7q8Xq155Vn5LHGi4fP8QKOFY4cal
O7pifl98cEDTmkqA7ACMHGAYy2Cv8rrWOL+FzDvkHGWv8xT9NflDlobg0P4G
FBL+E0fmLSNhbDwZIInCNKVLW224Bjp3J5GMYDGh3So3oeSlL9DRDcgz+UbB
SzZEyjzxk4u5jqQgM0tnFgIIO0Ha9zTpWLUX+vvZcrR0SoIZewpfUgN6FZhv
kYOYnp31W8WpyTcX1rZrAywhFQUKt9D1MeiuVocpbEC8bL/yBoRdfOhgzesv
XUMNZ25+SKE++Y+LtKmjzSV3BAIzS/0cnCRcvmDG8ak5Ne0qkBYdLJ6fjH/m
5tbtyz9wwmoMWTc+HE6I0YyPYf+dPByLgU4h3++JM0VUP/lY4IlNwl6H9rjK
v5kd8PTRYFHBcTrmN41lIY6F8A2tdi8Dw6LdumfucP+uY+AHVYmrjncXWQCJ
OZWsBN6LPDrPW0JpHOgFDMOSdRuVt/cB73tgKlVFbOzRDIHorDkMXy3IeKGq
4+vJ/t9h2fMz452VS5P2LAPzdnZ4ZQJzhbzcmhkiWdxAHOi0PaweyGFbRuzH
0xiUTORQVIv6v9ipoi7gkO74ldFzCKYaftGFFhb8X0B1JyFNlTUG1dtUMb00
+e0W7CZalxVuzu/ZW1fC8PIpxiIze6ulMe9ivVeWSEy14VGrNqLNVjIi38nD
885cp0L4by73XCH1agAwcnlbJU+arVn13Ctl95piI9IGDSyABrME+YbZ52c4
7urCqum83IAhjfq6GNyXECp5OM9fSnRi5VRwQky0Y3X7cqWQw92AY7E7faov
8EDmMcIuhXTHJ380Lzm8ZnomGVZJ0QtUG0TJvq+9b1vkm3dp9q4vjdd1cD7i
o12YjX3+K3hADVH35Ab9FuhITI+dmdD8nBr0tIU9ktRcTIJ6kGIAsUaUhZFS
A3wh2XK4i6LoYa0GqkbhM5os0WPnqt/Y3rQ+/vydo3+bGZTvTcswLROh81+V
4KH285sCDi6lZkGcwANoZ1Qjj7Ltx+QrRdkEilI1aBFDvbVPDJSjBAwLHHjL
DNfTwwIfsHLgLbOUsnLGCPIoZ5HE4k6Qo3QYpxz+NsuuJIZ6NKEYM1Pof9yO
2d3qkEJpx8jbbhb/bRufLJUgfZNkLqIy0iZIahcWsCMz/GniifzDjVHkjpPI
xoa/V9H7ijDyX7d7mOwOeP0Dvr5oPt2j8xohz3YlQwLI4OeRwAZt7rYXXo0v
whJLxnRxprmWGfKK6UNikqt356bvgHVTT6OHp3TIW197la9qvVabJzWKDRwK
3KDmZYxAJD/eQJaF2QY9Yzfd9AeUHYi1qJI8QLVYRsjN0KmQLwh+geNdsqzJ
wwJ1W+4dvzQjWJhEi/5GklonpiEDM6tM01TH+urbrtptVIU0sNz2F/Oe4s/e
Wia1OI/U9xIQaIiOTjv0glAfqNxVzJ7Uc22FUcCmm2Ftz26vgjZLUMoUedSc
Pj5JDJ25sRS3YqC1gq6u7fToIEvAKdGSwYBYjhf2EGFRKDFpzxEJb79nOq75
oV0J3/eLhCTh4xQCh4fnXnQi6YjK2Wl984/2ZNWlJBCJERcsCqh/RP2S1JRa
SZplYkaMFkHg84WWT3b7KdOF5vOoEvL8brx0WZ2zJWnnJqzrpMi7JR7Yrzwc
rznpx/dMfCGcC6pTegfo7ONlMGTdiGz8mNvREtq3EDitPb5PUbKOVuf0n+qz
CQ+Fh5QgQnUCJ7oRwD1hDviXnoCi4Xr9xh4g7DQmsS8OkEqUmrHfk+MoYjb+
zZAk0WzEavVeqtgUugCjv+tUsiKJ0mVyT2ysMMCCubTMa/WHXNorOZHmerap
WA4kBbypMk+zpYWew5xwpfoAArHievu28z/48yDFO08Dt3aoYlD7Xf3LrboQ
1RzStMm8+yxL2+Nsa3xXnYsDECBNC3wOzyLCO6QNVjUc787m3W1c84FNod6L
92lN6ukUUOXdK8zDjpUvT2LMP2KwhHAff7W7xhmvpOC2dx3VFOHN4DU6ydSt
+RQ924fIF18fV0ZUY1cM3gu70KS0RQ9ZgNuT+GeMUwZfaMSqAFh8OR0BBeaD
mIG8UEaza6x7vRwsxljwRtQxUcSFoyEcZH571Y6JU6ii6Qrrk9K0PBm19F1o
3aFveEfslXCqlwvs7iOwWcfCiDrEkTi3FO6FotkdPFM7nennWE+o8OI1uPY5
t79edCS3lcccI3eVZPlV0UxHP6tChlQvQMGSPpAb++1HHPQWUlxKGoZ/34Xc
DVgJsUK1xgqLL9m1rRvTen9+7z7d4tzQH8oEEX84IunJ3JNu2lGHuqMQrcUi
Rpn11MfmWsBlvbynQ7SufxFkJiN0pLknM+tim0kfggxzgsg2UxLErLHNFxn7
M5itgIRMLM8cYqz3KRJWii0khwnAWfBh/AvRKBmRzMjOQxHbHw/FSebGVmhl
zvY8YWAKa5SLH87EZ7u+8LAhiTnBURegvhrilJo/cc3Hb9W1Qq28mjIsnJFa
LceCJI30uiUTntwaDWLsCwMg0XJkvdM7dyDHz/55AeB9F4JxEbRraYsYMBzv
0/s1gex/j2c5X9AaZlmgDpit3Rz4mMbqcDlmuexmRe7JM4jbh7SR54XjdiQj
sWBqfW76VMzPLe0gFwsGbUUYO9VMMyoClbFPHw+EITduMH74gfcEbtC1TQRW
QMd1o2eJhZJnmSFs8rLj8inqGGXuyVG61ufmeGxwbjsrdCokD61KfHPsRO/l
zqR2/9LGaD54bdLa/QsrYRCsJ3Bw+2eNMQU7RbGr0IZpMXry2Qn9eAdXT2N0
1030lgLXKLqsrrLQgFyJRuNdiHyX9lmyeG1+y2oXh3+AyWq95JiUmYQ6f2Pj
o5xB89Uo8GUtcawFP5ELi/kfuUPk2ENjPzOrJgA7KpZlu9IXvTwlb8WABig0
S/bVMDZqi0pM3PlD/X2f7G9i715A8uFu6rPt7mRVAraorymmY2kVmvHAHii0
MbKANOQFbpX79qv1R+i+4PW5QAAYepUPSZyPUl9d97JU5k37yMIOCHUNYnP3
Bo3SuwmiWT9PXDWFquOaVZsCn81FrDax4h2iApPMk6LZWPWeAWjcEMEBLqTd
r7irpEn6BGscvl4olNEb7M+ZYqTKnHaMCIAD1cV8QW0sPZKxXaqrl1mpKQJY
CKhGLT+NPGWFZTGR/eMu/HfKO/Y2/rr2t3ulR4JypzQmVe8fgGZARCaE4vlt
Uo9poO3ACJ14dhp3arNYH7WKhl78QPPD2tE8eK7oY7cz+3NlS91XhUlfgNoz
FsA6HAGBOhtOIs2yMBxOVEV4M0sZ/9NS7+WoccR4x0XclxAtJWFcbf2MFHPH
ucM3kjmi1nFhXqkP9cwKk9OgyBt+BiG7CTQ9e3Fj5yeS0uA8O4b5l3S4mutX
npl1wNwyyw2oKL6eZ86o9w3MuMwWSKLmfDPURvRYHr8HcVbDuLjGrIt/OEp/
fYQUc05hh6GZawxNZ/RuoyLIhDg1fmNPw861nqzyFFnUf0g0qyQFmuFgFQ5Z
OeHfLdWsEUYeNMlEcLC5rdifeAO2mi6FTI0tfP6bc2Z54kBRWLb4zNyv0Sz+
4UBNU16NdXjwFcVHqRGfXA16terqxB/fWSuYWS2pF3yPYH8jc6qpOTAAEFOc
Dh/Ux/wheBknDon262fI3jsPVGeTqJyq8TWEPBcprP1gJt8g223YR2mc/Dnr
5APXnIISPAER9KfVW7cJc26+Vw26A2/anvbJBpUniOJzt3yFa2uaEQJ2Ztue
DS9V5rFa5/Y3AYK7MT7AQlRn2mUbz8tlQhCbmMiAmkKg9qPpeT4r0ZryvBzH
gkU4leMklpl0qDI8Wj0+IyK8pbraicV/vAtcE9IexKwHI7sCtWv6pKlBKVVu
Fx08TbCv534j8OqgexDE7wOdC93N5HI84ZlKoA13a/8QiEaVZMgcFmPYnh7c
4Mmyasg/R9fpJ71lu4RFc/+lsQZPu+EMGstAf2UhjvmznABULZcSfJGsS4pz
cp2fEwWKe7kZTFm0vC063tq+/HHp4Y4+lVY2lpUfnJmatCq98ZgYQXOioUc1
bNES6QRXguP6BIORHcifHwmtQB21T1REe2TSmDSR+aO5WnJwhcdH1ewNkHHd
sftSuWsrHIOYxsHjqQvMvFzZyDeI5jibs6+ckS9LxZSWSCKU9hOLuG1d09Zl
aqyo4BCGPN4O/fpOmGgkwwfLMDxXsOiLYp8ysq80oe5yhgExbHBFbljDlpqG
igs9yOWQfARhP/Du0Qg9rxE5/iOGqEHdLUhCwiFSrEieWXcKhiKcVGthSp6s
QAK3VIaDfCqIjPbHMNYnWvdwW768bnuGkXVaGdppHUR4NVM+o+FU2XnWDiXj
zl2tXtO/krN3+gxqoTRPsw2VLg2/GU9q7ZGQzD83ig0y+racaiiYJNy589Xj
QXsSQPxc/oOmwkxRj8hfizxbLiN48iN6L5QwRqmvllO6OCYh97zXJcTBIEBh
z+mqOpmRsc/UFRkcDABTYTMLrcWG1mDBX1MuJBwt7nGFSPIbhL0OL3JiaLjR
VJyTs8BJzaj49gXAjA8QAWvIlgPR3NAmLjkYo/DD1nsf3lWnkEVNDtnNLFv7
jo873ddrZNSsUE+kDDBj6KdpJDRDyFOF/Ol5Uf3UZ/yCfJppwC/+0w//5jgf
ztbY6u2XgF/ybGjdIWqexiVeYXpgNDZGQqV5tPdIF04P/IEeoiX79G+TnARp
pNbvobyZ9dAP3chZY9tudh5NX3gg3kRg8DfcF+hYLvBzp+vp61mcW9KuYG2Q
N0CrA2uVeStWm1nzpCuMyYWWJyH/P37zwiDLear1/5QqlchTnDWIM0MR9K2w
/O/XWXVlpEEQ2EXgLu+8QYtp5379qvGJ878fI1gMFMfprCJbsRJvY/MazP1k
4mRxWsTroLoT5ysWH42rGfUWtL4HiKDkE5TeqodpEvkY2ZFM5TnJT4q/8jSe
uEedcMNTSx7B8gEbS56FIgGgA1AgkN0uuXqz1wDqXa116pyrhpjJfJnNRgEo
qSAY1VhplrNuxJvQkY9We29DabODicliic7cPAG1y4fyvwemp9iKf8aeols0
yct8v57R5u33Joj+yF5ztd1fUfVbWEy9KaHvA7oQH0D2s/bewjDkxvoTTvhC
DIgxUzsqeTo+eFFiMxBTJX/7Ku2QVQ/5E/U/owlX0HHwZUKmHTxM3uDHu69E
7NE02KfArLCK5nPaB5krlOE9GqGOrmyCmcNKf2PAUM6dY7NouBQa+zHtcjgi
oiuGbCyrO+rAAeRlW15ujEmwIoZYJUNzKJU/WGc7oCa/FvCyMpkZPngD8YdU
x/6YhEcErU0N0WFG3q5RGemQOoIU0iOHAOTPR/2iH6FoqLZSavgJ2d7gUPtG
FTnARYDemDuWputst4nH4gvWiiMbowuzmhq0LDMc/PcoCaAGJ32m0LlfOkwR
OvnlrROCuKvhReZdQDecVRPBebVtJLH55rKuRkHTzSatP3fq6IX8ufj99dlA
uJdPlvRREgGd0SrP7EoBz4NC1jWuSjixdLbnh21zCcTsZooilOmqGOvvgWPl
LJ8Qo3BdhTrl3d8t4ETaA3cMh6RKFtP1i3qfQX9bdxBCZBXiDrtPlVu4SXNw
fQujqrG7gZM9W4UxDTWnhVENxhZ1OZ+05Zy92Ej1YJsadCsEWKiMcGqB9mIz
LzdgRUL0rHdj/wZy+Mx2ZUaWjgXUh4QlNS1LScdS9P502PeS0WmdHi7UHMrI
Vup5cCrMjr7zckMidLFDp4mtfq0rVDOeezFMMQOMheKUMwj8gRKwB54+WwH2
ArodWne7D5scCKW+Bc4SPsLWY2r56ijTFdikUDTBh8CokQ6ZsAC74OC11cwu
6tLmNVf2tWka5coMvfzs6u1KB3l7B1rIPVLJO0Y73ORXQIUQujO/SNrM/ZJ2
PejYnJxEcdAHLvy6XM3TZFo2mFoLYgvnbtnpBh1vvlV8kjYZ1jPqsvi7rilY
1waBqz4WkPXNLhz1YwB3QlgqNF9ZuZY+xJXlOoZv+qTmTqfhGjmbe90Zox9w
j165crJx63LsNdrAS5QEvbjBqXrzpngyvjfw2Ev/v7l27uKwiASrGIgOcpuQ
bHma3TOcc4Lpg00Sdnl39JKe1NpBWk9MV7WOlS9NMDFBFjGnCTtFoM1chEwk
ppCc34k/gu/l1+d/ckfrNEzttuUvs+vM6jePBEOrSeaeoIqeeBke1xA3UCrZ
pxMIO+uIODEgFfRUsSIVii5YEyaiWWsBiCPbWylm+J0suNl8B7jk8Fu594EN
e1SIHuWKbnekxf3zJ+yo4ubOIdkLZlvklf2uEwm0Gm0wn2LNGrajj/dpqgym
1yipaK8TaECPTVW19IGmIlPecnmgJJwaXs8JSUWpkUHIzH4S/uvdZAgaMnXg
LYD1uP21tnGzzJmHsmSJ/qO5EKH1IQ8payHtGqQOqC3l0/TjCPKkEADgG3uJ
E2nVe2G2X1A2QadDl1xGPCR6K7xoxpjhFaLZgwNm8v5ryYAzwzIkimySQdoH
apD15hzLpqtB01XUVuumzFo7VKlJpFYvmN1C/0JIkNMaJK6bBjGG/J9NpKA0
AEhbXuVQKU7BXJZL/bocl9AzjuzleW+ooH15qLJq/vUHzT4g90xLNruJOTPH
kViqlQtLrC6AKm17f1AyHTsZO9wys6X76gnnQcWyO2Ez+rFlfWTmhVPP/lv5
5Y2rgjxAB40ssXyG7XMckwvuxtqmNrdH5sadk1qZbBK1ZyaQ4dQntpNFvq+6
e7JwzT2MSCwYul8OWfmGB8d7JLrz4h9OX+ArCVLBjL1SmQY3TFtGGbSUQkXt
awnBxKHLbI+BCbwaAoxA+3BpZcV+qFD74/eUXSZi9juF2Lhp39WlPIfoU3oG
3ZJuXyg+TpepN95GlhPWjQx+S7Di0Uh4gNAhrHIXX5++rm1DNw9SaFCI8SvD
SatqblKYcUo1HfVChcUznq6zDneH+PvYsYnt6u6IxhkQQiZn0umLWoGb2j7s
6IKlkjYrKOUvpFLiM9Q7jOMSiPlBShVtSpD7PDCIiqUyIagTiToQHD+4DOnQ
vuANNO/k8OUZu7Qc0pZ4Bw9befXYlNB1WY0c6sEKwp0mFXPXAWLyCJ57lJNb
637bI0326+Kx2QhAPv10aE5krTsrn9L9nJ1Axwf1P7LHkarvH1c5R7vofyiU
y91TPQsRC/vO5VFWIfhGv/BjFGx/Y0M/alkF/lEYRjyQJnbMQm2/MAaBIn80
E15rKj+7Shr6Fjqce7nHe5kik0YHpkLtsAsCYLgPjXYbr2dTAnowfukVMNPw
Exd5rNUJkntd/xEy5fR6Wp0DHrGf2VXChjERgQ9us7kjNFOBXD2E2CMe0kig
IumNATxjAMsAv0Y+sPmlGEQAZ6nbAzoK3ubLr36szuHV4e4ttQIri9XtPFDt
iac/ZTl9lwXlxNtkT+TTU6MufoXuZOZB8rH4q1OP00aNbvTfRhiCWfLK0syX
knQIxdjkQxlaelDXb3vKTAJvM5pzObH9izX6TKF5L1M4S6aaEs/LtHBgxEok
TMcX0pkQaPxUkQpmWQOTqHz5xwhT8kDXrDa5oYaUYmOjKHTzh2V1nqVj5rs1
Jb5Jzczq5w+L05xJClTwvXkjFelXrHQYJ/tE1HXtEDnoevu8txV9k+9cehOc
EbXja4gPuRyyriLTaO9lToXY8MthzUSdDsH9zsjulL4/Flk/nPFIX5QKGV4+
FirDKieDnPHTeqaFXGIZsm82vSD3f+0fHnJVlQ7Ub/8EtO0/lItNFkPpS6DX
g+LulUbMdbbHhGmS2R/pcASBxVUdcbx+FCbMUM+Ximx/ZD6XcCp3AIJmLTqV
AxRJ2WCFs0Wbm/n+6mrYdrcUcGVRJhADYEGlQSTIowRJGUej4QcP86dr/ejP
VZj+j3VftuRIphuVvkDp1tHc4nyG61gyYvrpLZsxlRm9jV7OIue9ijU1YNiV
KK8Pwm9DQ0Y/LdbSmrqTygkrHVWyl4J6bXO0l+F4HA6KppXH5KgVl9s76Pif
3txbuTXWOH10KC1Rpq0ioJzVjQTWR9vDh0tQxySpRGjp97t8xexBFN6a5rQD
rBnNp+0b8N10X6715zeT+8obhffQu87QCQyS/XUWhrzIdORCH6glwTIxcn8c
OQaTCbbvN3ckiYNMCRfk51ePVpHKkJlP774DpO+w9jlAUEwU6Zl+sx+aGqse
XOcIx3NLpkHWPIiAyHNnqt4sYSxYufqS5GQSg/KKawjb/0WJB3+N8NUO0GqK
BRImX+0maBo/Hm6ePOm5eNhiX2IrWBmVUpkp8j3hXQp2GLJ21qGMspblS336
5NEEOqWYo+FRHzjpCJ/c8hZ7HSb0KLelbRjA1QFKh1Fzoxtb4CIMXhhp+Mdi
cZX7ECLxrdeDS0x83e9Q4U7UufHJIEcIof2SlS6AynJerBv0qn+w1VsUIV2H
LQ3f/xKvdAr5FF+/6deqV/npq3LQ3P0LEWtAotHAVyPePtvc4yVvtBgxwss2
XXgbwLZL4Ir4I/0UrQDz9+b4ZPSlf7A6JE5PFECBjTNqPgrAaQ3BbF1gmE15
YGagDfdHOZ4or9BM+7+Ys5+qJEDHcpw7m4VL5iVSM/fAJmIBl0XmPLppQl9o
2w1chkWSeIuVx2oCMWpYbHiyhv6PW8J2pShtui3jcGK8KMZ5FJ84vixKqiv9
QohvS7DOKNpFZzYw9XoLS4ntwiGqDcuZRveq/J6lACLOAtMMi4RLuyC73H85
+LvcPIHjO4kM74EYZaPWHp5di7PI2mZanKaDLbjv80AVxB3QW0aFeF5gOTsJ
8emy9jZWjbeaiZoYhwH/d+vFDhJdLz4QiczEpSuCW7ngABiHs6OWK4M9SSUW
4T84f52dSOYOMMFBALlpY4JTHw/9zGJRkutoosAIch37YNBxGUs1+qrkQH2x
e1mjtK9CKl9MU2sXWbspLyR3XWyv5ruETuYclTy4yGPgu+f0cwoN1ABtxGqA
oAxR9cOfyvnbZEgbNuzGUYGIruTdbmkTr4oeYJapeEFhbl3hgbktD4gop8Ii
WLGdhL5fFIOk27kZfnHa8ufYAghfgAzc6qmspjNzLdmSUagA1leOc1oHrcJU
uo8Pts/FccrUT3TP2XENXUWkGXu422cnjyCmMEXoK9XycKsAkicmnErLP19J
qcnZiqkn5OS9/JRszk98nQo44zJKBk8aKfIumR0dtDpozn4mLkA/a46vUZ79
AftEu2X+V3PKi2OAJ1iKZ7jUcYxw86eRSTG5VF4pxgD06mtuYs2YvXDFMRso
hkX6VblfBweXJEoj1fkoYchnvZa4BeiR6vSYivsDGjNqzHZq0cDxRbpolFCX
yFqJcSkht7oDxzUfhirOXkfnn0XMH2h8nkuk+YBMJ8u1rgXqhgd2kB4skxCD
wq/yvk6nKIh3lQ+sGfIUnSeUcUY9i6lq5+gHHkSgj6bqsw/TtM+YTM3rZqz/
HD90n61V0rpAsNWMOn4t4S9zsaGKHRN3Jcfb3Zto9lxERWLco3A6RXygBPE2
UMQZ4e6CuDZ4rWcLkZatByuWnZ/4VBeb0uUhA7JhjmT1JcNZHBldA3y6vKlx
tguI3MuF750vETkZHWvmRVe/L4cfwWphmLfRPhqmkD6XSEmKJ0RYBZr2RVBC
/3jhLmOYKcPELlVF2scCgo2DVNNUDK2/VLe5+m6E3Crha4/09zlZFToIIFZc
zkxrPnjXr5tSJn+46gJ7m8Hh9EmPzEU5+uxpesCBeD3s1r7FtnLfZruBSN1T
Msg4//gzCPPPGnJhQ9M7OeGUQLZ6u91LsMC/+ZbmmEcFHsfSwuMcUjC+jn+T
LvKfFerpqia4GHdfpRbKFvW2lMZdMnA4fa8F2TaMeuzSoDAW39tBo07mQuHF
g8d0ByvOK9TLOM/OyQab7s+h4eLkQA7pvUAA7jn/hGocy08nIa2/lEeZ6OdR
S4SXVGPdkjb5i55vpDo9o9laBmNGE1cK018XHhUR8uivwk9AIl+sqtpvrMgN
4B73DFxzsUBK6979CUyd9Ab/5fVXJn3msln1s/WFrvl5cBH/aWOvEz8cLCkm
MZWqGhdRWrI4jnxJw+3N/Z9KYWd1V8FVle+tp2DQNYiS6HIz6FquxsStV3sg
Ukzu6F7MVfhIzWGTJ3GddmhOfvYkqdvEHquCQ+zka6Z9ai6qzB4bTahgVgLs
/WanrT+3NlRxNL5alT6iHIA7dRC3SbTlzQmNmZ6nglGil1hqprMZtfZKYJfm
7YxfX7tYsMBVaPwD8yhll9X1Zu1cjHmsA84h3zsKTtFSb2/9QuIpd4WtAyYx
2oV8iMQX7/Mro3O27T94TGRj9tVwA6m7OsY6gZgOlPUAj2+I957Lcmbv0+kU
sZoQkCUKLP6hYcy5KlgRnlKti5TqiU9ur3dYxFLoyaxpItHXud8/MZGAjC17
KFT99RSFYIaAcBQ3APmUvcCHD+8PIG3Xn0fx/vHYVbw4aWjBxrSLLDezixbK
9rX/zROpy60qqSqfin0YBC1OCSsRO24Pk+Q/XDaqTZmdnr0r2TCpsjL1FxOu
j3rROmaQglN69lyrTgbSw0Kzgym6qM4x3qq19zUkTg26YS0Y45ecskYH+lep
I9OhAU6mJI2XuJaJtxFDyq/hLbcJXNE5OOP8c0g20iwOqMacClxaOzvSKr7L
E/bWvTQPrxIzdmHTWhxSrXqMFmAe852CGYHBbtMQL1aqFI+zJA4qWWvNJLDw
VNz55hznCsDJPc3LAbaF5M2lwdYhatpjD/aRdNQGSjM87GrnzLpC4ohsJwXh
B4eKYzqXX/0I/nmtq5UA/GEcHtiX0+5VSw8L19rRtVjSoqHG9min9oW1bHX2
qhtPo7nxSXUcjWvpjHl/guGjR472ILL1mgs7775t/QYlg2nRqxsNt8qOi3EV
rz0Pl6EAGUkKW1PrimSpxnIGTQX2rUpL1X6xfkeOdXsubUPWJqMSAjir5LNw
f6vZ6CXikQHtQ8MehkZTMdZpEHqELtu9wGT5UL+5KjF0jDQ4OOd3VU4HXc4o
BV4mviGw2t3p2kA1TIoL0bO5KJKw1cjXlTzFUvfH1gGeUFgas2QMlJYveWtc
TO3HK9yKXeXNeQdSV+i8MsPyv97NkdLkUSp0X75TwpRyLHDDF4ywwNB5Twd+
YpZecJ2nSYbf2vMrA9UOgmgKeo2gAKAgJ2ZIcLWgSifFTkMod0SLjEZ7+S96
FNGt0gW9DtySQIwSh6+/hD+mHVKDV1GF5TV4Sa5wpLJNlB+3MlaaT2pTzcXK
j6NLqMzZWUefCXgBXIhYuGzihrcneHryRHgsAZBug+P1vna+rq8V4+TORE9+
nMUINmbeYMRxWqK+IV7iuQR58Ke56RjLDULHcZy+edVmtqN/0rc8Xj9TKcze
u5o/xPq1WVTbR+RyRYGNJgt33HbrHYsPwk61rcuBrsGOBQ1aGseQoAKeccIC
w2DEu/8q/PEPZ7oaKmJoVeRSDpNFuq7uhndeYf1cdVPEJYNJUMZSqK+EBvA0
fab9MKRnP5Crie+fZJrnD7y131qvAGkxk3ok5PYlI9mrjMOf1en0JHMU85Hr
imDU0Wcys4qQNMIcnPAYLD5oxfcvoEbI5RpYDH3SUDpMcrTY8tr2W/rZsUFC
cv/1XTCOYwbfuwxNW4bu/Da7ZYfSwtuI17ZvUQJpWriup6LKV2bpWGSCO+nX
KWWVnoWRNWV5REFDdP8RwtRpacaoiuE3APvh5bn7dvbvRU+cJgotSwKdfFLS
AYaZlSpCIiVywturSjOnETk/kgeY2/DG3bqefW8ttZ73k32IUbfR7dVYSihe
F9iMm+I3oDBajxsIaN2PgdkyaCw9FixRXs5xfJghoBisK5QaAvD5T8ZnfFqo
juVivDSPrsSHtBtoFvvHSysWUmAJX3fStHEX/jD1achONO1ldVFhjLpy395P
hi8SiBSPwZv7kCA6yYtwJx/g4WBOsanLoP6QMbx9yEUA0WHvgSnVu1Y0o3Mp
WkoRt26wZunWaS6CBT/hQ3FAIm81GtDe8dE6tTE5lptK/QwwSQHj3ToVnTL9
4CcZDh3Jg9qWEAVIcSbj06YQ/ptUZsz5pW1X0JpShcKtJ3Ylq5QQfhwQDXHA
czJa+EwCz4PgnHMqVXDKwJo7PHxs5gb5CfaGrkU6fpiWRtWa4fY883Ck0vlm
H1ibI8OJMcHERfVu3ruXc+qoOhmW/FWXlusC4QHuiB0mLatwjaa7UA9wCKpO
5FlMUjumCxd4IOke245x+7Tc8vg6vj4tt9UfmtSUkK8WhWm91ld5ruJ+NdPb
Vt8pn1sNVTFQ8hFuqXOofaDjd3bQkXQgM3XsepSYwKuTsZ3Wdh1nZ2C6oH3K
21JKL9wmBGrKaX4xx8GzseX+DL0EXwHRL9QuIAqUuqIH9M3u9sAcmvh6sTgg
vEgewi70ndwZAq9+vmvnwFMPsZAiRfbaA+/Ffnd6KbZlQj1whKHygPJrkOcf
hebLdd4e3xPNHG5jzw6wqE39BHSmvM9t9JvnNLO5yNb0aGseXHNsbTe9cW36
AihyBf/C4pa1ngcC0LjuzIR2d+vfbdXPRB+ybSZj/Q22mA71ByKJQMN0SILj
9yP6xEwAJM0wI7Owft8boQ52V3ulBe4hOo78vbvdDUWMZfOSGI7sbXzBT2gJ
Olp0qnb/Wa6rZlww16sCd9koRbWeHusL4LOlCo6QraH1z65wBTA5CTFpyoAt
0oqev9hbbi0J29I/4q9oH2Z028IGRJ0okJ7n6ye5Bjg7fSyZDQ3f/sLiubhA
KBezrhwQRZh4w0KIXMGciTP8Uq2mQ2UW3j0coSVEELeUQ1Nm3N26OY6HJNSJ
6xqXuF2nNe/J/NBhBiyGr5qTsMh+1q9futXf3vnx00RxXHUdjuKrwg6uZ+e3
Kyc9CK0Wjj89nnmLcpdLtW5EuPH0m3BShCsytQyqfwEA0rgUvyOTcrsu9AY6
IbJonnXoM+0VQ+YRNuqXWj7H19uHOHlQZ153/AqmFc1uWStGhwj0WlvZzTS5
bxA0OH+c9W/8kpyjm2GW34OkSMzXvUUWL0+nV8yBWifb6rga5vVOHqYPx5F2
v1hjUHqc8Expif+JjE3JswaY7HEFrMIWSu+QXD4RhaYmiYejYffJ6Zd7TQSk
PquaH/r82ifClt+OJQ3bJ/7Bis2UcTFAdFjA1fqdIEkLfpJuKOdhryc3meNU
ULIUw3coCIox9UTy1CH05/+gtMGTVZlRhzD6f5dqixHP/s2xmfeLZd4Qb8k7
5a01y+04Mguv1QyakxpI6RoC3QVUB8cYautPdSiTcYhxhsMAYmlBphNq4zJM
rBASrWCFEJgDSnAv4k2IDKcefi4v9dVecsCMN7ZteP0m+0LEc1M1GupRTnrE
/q3WuKr289Vd1Fc+m3I/lGghWNR6q6klfY8gducgy+i/WomZ91RgJMqIvdS/
OzM+F6+wkdzdeXOo3Y8xusOyoBJHg42e/8YjPpB6PxDbYc5zChesKzPtwDpz
N1+J+YAMJuKi0pbtqGTeSWPbRmwNxLRji/ohwX80jqSQ3fArFezDi8igMlNB
AjwMkhljXhv9s1LfVWLs2/wzeU71Zjh/Mse86rLMjysDsKpeIwTEi6QsGmoY
DcVLjLqz0+HL2Spvz9oUVz3+i7WB2KVvgdXeW5yp13fhQvS/TXMmIMYGd9/k
ScqjOkkwcZ1hHMQrY60GR+6kkSVP0J7NEqu56ym0iDJ4Dpjp8poGS4fqbSD9
Do4OwBh/u3Cqo2LP3PWbgEpTrRtLim/W0vZch2Ih057kysoP4JVcT8UFGpYe
Xu+S1hRG0BcK2Amm/Q6B+jI80KZDbgaBCThpfiFpd9xbuk5pyu3DHvQlWBcJ
CbX08TTIp/thcrHsag8SCRAQSx7A0On5SnVswfs688wRiBORO694uTK7fFdj
0BW9ALvTRe9cVIo8dlwdnVoaGQncHdmDsS/WwoXIX4bWA983Xf2vnA+lg2tt
Il0PLETMiK8elLvysV7+Jps0eBjkoVwOufUA58S/lqKo6X++NUCwwDl7bqH7
WDoPVWcPcKjhZ9gxlLZTwRJTQO96Ufp5WONRHBY6e0ujLDOXzKDlnnv89P4O
Yxts4+LhqvrW0tWMM9+ZVXWhgyKKbDYcuZjoXH16UsJnVXJ3u3rBMTrI14NE
PuYhTJCxRBTdql2A++HBPSLRTHeyXOb0HtFKInpSv9MLdSxfHj2XXcnGEap6
cU8SAGo+Lk7gRf9lVA+3RdsjqE6R6U0nVnZWaLbl2A90FsP2gF2e36+aKS1L
HQ9XYc6p62HZL/N0jZy6iv7kL0uvUwBhhuxQMV3F4OpEkZms6qyKD9FNzEFT
V1t1IAyD0oKl8ZRmBmvtKV2Hojnf1a0Rps+iSSO5HL9gvNs0qoXmzu6nLYNB
bPqN0GcoH5DJdKusTpWAOo64/LzlBCCwmHMFUynztwlAEpw/Uu6Dayh9MvJk
ohfx5iQO3ZiF0skcZ6xXSDAbG1s0oVbfkbAqIRFLiMVRdoEdk2Ul3+/jHz10
Y3O7e8eNQPtKprvU7NzLKr+uATSQlRGI2LxU/ZqSbLwjDEJXXGhKEqxrWdmV
GNyU2l86goi8z/fBcQH5lX160AG4bobW2SmluxJWZA+eE2dzuws7OmCDp1vP
o/HmT6+eVe+9yjTUuEA4eRDDsyvwf9N0YFnMvCLqOMTQhfstCkxEOK2GnQNl
7gaeqSkU4sfqNzPCFqGdyfya/1+rsCtBnOQgmhzA9ziRFuSecztjsicGFvPT
xpcGrw4oT11lM+a+tsbkpsxAL0UPvA7X4fVUhlmZDl5dg2P2pRGTwmWzx+BL
Bogj/nKXikAukYMGxeWrSynTBWrCHYeeBbQhEJhjL8U4i3uwg077sacw619h
I1CHO8HjlX0k0xdCfjor2IfdK1fxc8pt7808GCrfEl0JlxtMClPxNsca1Z3i
710EaO9SchUFxfMEaCmXs3TUwiWuEB7pzTXW4jZRcSpgXG2o+xao3PPideiZ
VIVTDZZZr63S8TeSfYtAtEKyz8wLtuj349Txkl2R/rVf2vwPOH0kzpvVYY/E
VRRnsKqzQYM54QtaRClR3i4yAM4cv59kk7NefQr1cnGOKsqa5A2a1Nke608L
GX/H4UhO4vEaQr8CJ5WZmGX3cmFs6bV8IyuDGxGnsUeVvy+/2JE+3cVEM308
rKo9F4mGwcd6pQ4Dd0rM6NZDWfEp2qlVKEPEGif0Ot4k8EG5AL5Db09G8wUH
qENaWNrbEhLPRJVBvM5+uyupiPBK352bla8CpVbqNHTGAc1NOphKccJlOdpK
QmKt7sZ2C/xXfERa+KmJS8JKxBRYIVHcN3yZ4hcWfN6cljvqaIuNQLSwkI++
x2Iu2WjAb5DU7R4QhGHsp8DMmUxT4W94FApS4TdZhb13gT/PGmAUvz3WFznd
v9vfK5EeMg3Y4ZwtSihLp8Z+sAyWjA5cXeg2B9a4uEIL/IizeNuaBinwVDGB
mZH6PWdI0xFwcku2dXrBE0E2biZZvlocpRkX3tezQxEW6VBl0hJ8LWb4mX4v
2GQD2RNZcgFMZecDQC4WjcIdSh4EOgC0tc/xRLRmT1/Zwi0WRiT2tEooxo2w
R9yD8bcRDkv4e2vsHwZH/sXys+eTpg59uXgShyawwhcP3yhh0l8ioTGWTM/O
8ef0L9LZYZG6TqoAa2MnGHU3Z6Of8MnOcnVevnEjROpz+cUhNLrbOBG1sHZG
/fZIWHQieSFLclP91hso70zsSTAp67HKBQo0jTJ8vcb6huvOxJRml1hk27Bp
W+VeUzG5Y6mvp7Tl7KkP7YlxTDhhAE45unCJXcMWrza4GYI/5xJfliQbAF5K
gxCWr9apzmZE4M+ULk2wWRgn9fnGxPONB7ClLxs3/0xBkFPAHdG7+ocUznWA
UtVe3Vk1iG7V/gYlatmY7gGbKsdLYRqVqVdk8W8NhrXxUNYPCDLkTenMFE7T
aPex4L34dFdgy9z8dvMGniyssAdbYhx779rEl5clpL771a+CmvhhygWILPDc
OR4Rh3mVYpCYffSyt8AHvc//duX5kPj9aNSRiBnHdtNGV4j1dnAzgw9BmuSY
Q9rQSjclEZR/gDCYOWSzd4zHztbY5ngXVejtK7YM70xL84ayyn/kHt9OKCeF
+aY+/Iyn5EIaYsnsUvtnRB50mpaXhR4htSOHvxCSIoJ1rr4eKGQUnjQY3Jj+
DsBtnNnKt3zJjp964hzyZ+XGfA5q0tJ4sJVSaRNK7w5h0zGG5U15TN7z778l
X7ZZNi6WI9k/Ezf9r5hpxa9QDDln9tByeGdvnZ4tzd3iCYI5deF5np3a6R4a
SCPVzhQsYYRvmPiG9qXzWhKjBZAC2l7Q/m4SKZxEmlebJB8vFQ13ZRhVfCT3
it67ujpKVAuxJhuqdnwdV+6fiqxqWr4Bmr28QWXnmmmrCZPVl+zxBh0o8KUx
NdLft9cIINd9pSkbhqHMn+tRcOVlrJHwl90WmfxUh9F0KpC9VUmkG6dzZmBo
EZwkauMB7Ja5WMMRoQRMNwYGvgh3xkvZrqXUr7Z71aYZbItOr6Vvbymm8ErE
SlSxTC0L06y6a0IndatHQndrucnBN1YOcRaCAL2DULtTDM0GwFrijtFLN28L
zcT5T6U16HIxI4dvWtoUMvQVFLJQ5Ue9ZU98wHQbyfVHR8I+8nwozptTLKBX
RvFAIPReYWdBiV2l94xgt+a5iNEJQ/EkuPpQU4k22nyiUKeH6nLMLFpoXLU0
Ir/dzcmmU1GAG2ajbnp1hgLuB7kM18sQ/S4J2AQAdT4U5pUrzl3xOfooAV1D
znwF/YJ71EHS8d0VT1uvYyjAzMkZ2YqwR6eoHbCGks6/GH2H2cRiiXTTx7RL
28UbOtg77PgtWD+tWdqT/ki+a7DrKeecoLslGKe9FP26Ouoy3SLi2p/swvNk
RFHua285dNuWggrN+gsX7lSpxyjMdAXzHaN1C+tWpnBG2o2XLu14adrG/q/y
7GCODnZ5Qxzyb3wXcD4ix2bTONwL9yjIQbwD1Ow5s4VcVR66kzd7oDqfz/c8
rgs9rhjKk4crw8aT4gvewgZKRku5VJR60CSPAyezwIc2O0CAtYBbqFDR+Jzp
NmfOzjo9D4peVHIGET2e/E4EHVbHuif5BIHMBNr1HY3Eq0nwXR10pmeY364y
E+RIEIT+aSe3RGvZ3zIVT97mt9v0KMISTdv4gjD88cnu2TL89lg5/IJ/NfA8
dykILsSKD40sy3EZFSW1wEgKTE6tKcqGNiYKfarVB8ATQExfTc8sj1PDCZ7K
82ZEmiUxduU4xlAMcE1SLp8l+8f12QwqbnvM5Twz32GH2NFQCqNeGioIYTKU
lfrRr6BiUvaCMYxuJKnX83G7btKilq2hKAU5Ksu5rhu4TreHxgAKnBTwXgVY
N7iB11BwJh10jZ3FcSzH4k57Qy2l7sxtFlxmW4Jyi/Yf/f0CdppbmWLYPdJD
UrutvU7SPZaF59rkVt8cr7MCwfJONOge1hZR2dowGMScenDNDUXAqede6GKB
mZSBS7gFxkdtTCtDe/WmMJ5SagcExYsdgPozVNAAQrs+C7YPQZmEy1BbET5r
kNrEHt16qwHfEsrXxlrD+KU4Jp706Zc1bQnruNxGakVXyXLonLQY0xeNLpdl
KqZPBsMP/W/dWDYbuZ+Ba4jeNrPuhECXSIjuG7ktb6KyEeeg+Q2nm25Tsy0q
udY2ObGdiYIMSktAgpqGbH/mmo+0EGqk20USP8jlw7g5svb6PLXJ/AARzTIa
heZyubNRvIROdxX/wUdsvRhMTS2podElpg/HjwWLuo/Yoc4VxBmTjVWoN30g
R2RvwaazHDfOXzeB2iiW8pur3Vij2+nJ8lPFuYw3iSJLvrbjNwvO1b9xGvav
amuFVskBt1cGCcXKlVlOUGA8J/j42zlNxDICRpGVKMfCCShidwY4rdHYu7pk
It2MT/cziSPQd6GgTSI/16AJHIeph09F6LgbfATmbJ0vXQvYji6ykuSOhmyt
t+dDLbqe7RocLzrddNRVdTlmz1l8dMB7CFDieL/uvh0IdJ07WaMEdaFWBtVn
ueHgifas9LM/PgK1/zDN2Cnpeg4fVIlxheD5wu5NCb34DHujldXJTRawLISn
Umb8GpBnzTD1yX0c7rZvMj4X4o0ICnTqcTsJ5WyELbEy6LbVwXTiT3barZhx
WiW1d6LCZLp3OwW3HBqcCB9LUtkFjKeUq662w+vlQuyWuhSBEfm55I6IHLtQ
lNLSYfeA+Zw1Putgq03nSmxWcbkxIboDjCqQ8BZ4PArSd1WQv2qCBNIPrBAi
DHpQT5XoWj2F1DrztgFn4TXoXbj7i9tFUA6q9ixAdH4nOf7zKzIpIvGjsq+d
pClgVhvLA+UPZhdMdv0DBzgURplWBQFnUINHo3gp07cTZudEC2PusVgqg/B1
ysCEDreOZOehdZcGfAj1rN25O7e6+YlS1XcJmXkEkRUJ3pJUNpTuSspcZs40
CP7TG7pWpMH1oxQqQK5DGBAyYY7eAzc2uiVLQpay/Rp5BUAYzGgzJL7zTzMu
1CfZ7ZPIUq3td4CZTWNZo+0eAOroX0SH3AWLwcGmquFAKFkPVQu3g/enxH2n
QZlQYBcSMZ6V6al5aH1p9nltAQm1KMUtQcvr9+y8bwDcHXmnATnNpN1pjtsT
D0LCC0LUyUin/EkEmQDApaiS1QVsdSwMQQdC4z49rkW2sxR4TFRr7Kviefgo
nmkpnGrSp/WnRg8z4F+OjmAthzDnATom06hwh//seqmQ72jBzD/PYPPqQ4fQ
ZJnwqxGGiaBwYSDA/V759PCc1fU54jMSGybPmTlhJ9rW6mL+sM2CauYYn38I
8NtuRXBXUdPsQJK1vPAz4gL6MkHLyrXnjCXYiKgEM9td9NgVDTEONt/SzYpS
2o6okNTfIaR5Ena6hiuqBr/cYFUZ+hCWHnxgpuc+twPgwGPBFDHXMh0NXHIF
rolrUD74hXXPX4t/x9jbN+wK/rOCvTKE8VA+tSrLv+6mrVGF9Ku+26cI0+aI
2ICkPBEg+fxWYKQcOfnD976rYn7rB5+3fU2LM1+RjOQEmoWW7/NPtnBM96pR
H/7Tp2LaIZ9fgIK4WBbM9cneMd7oUk/clBC5RWH/M1Zl/FJnFsNshZ0EnrnA
L/sx2W1c0+c2t7V9aN9k8wGRdpPtKfIU4iGx+n28jDHt/JlFN9BwZZYD1WSN
WZITIIDjd9/aI0Jw/rZ3eHRyiU824ZXOA/mxDgh9c2NtiYTYf0CyF1UD7DpW
AxuWiwphTt4lh8Ulr4Ln9pz4rM5iG1CBx10y9xS/0jnX1+pverLQNA/6dEo2
ryZHJgIokE4VHBmgrL6oUDA0w9PhB9brtuIhFWFvYtWUARGSTCVfqr3xGJ3j
OPanVhFT8yCPC8KOd+kD1CFVTYZginClTGSqb+WtrKwwqHjN+gZOqG/6Ll4K
n3zq9OCJpmL9v3rH2f7ZyIETCGdHa/KmOGLEVN1fsE7fk+mMp17QmsyVChO+
d7ks7in54M92mZa/QhKjrhwOwyLvSqqpKS2kS5OWEikMCwpM8O3t4YMILfxw
rGPLE6xN7/lMFunWl1ciM0/7XjIwd8g72IvJx/P0wypY+jTzZzh57QPRT3OV
5PH7+TsGR3rcOGYAxv2wPoyfDznvCcIKICVlCsq8yb6aHze2nhQUIWlpT3VZ
4XocpQXZ5A+dvVzksEAeaShaw2SXU4NoMkybTGe83SETvsbSniu4g9Zh8dZ1
rs8yd7IytwLPT83+mSSaivvtKg85XYShu+cJK7MJJlaXevPYDE1IAw9qH5t3
eRATLKu+aT5x3UQh/xlAqsYHkQlMytJBt951HUBWIAzqow+1ThkRlOKtCGyt
TVAogfK0YMv6QepYQOHz/7g03K6FhIrRwgiVq0ooF7yvBeACYrLP8VyGfy+c
gfBErn5Kyj1zV1rWwOv5UgTlpxrWsMa+pXGd1SzPBAgyIIOkuSHVZMAByKep
iBevd7goEYCEJ//Vxheycelmgb4mKlexoDSoF0or7XrmjSWxUfoBCBeV6l33
51ErYZEgdpJvJO2TFVcBRHFVvCa0hQXZUU+segTw0R+YPua9IznEPVqWWvVG
k7ggV8mA9dqujWRjU6inhI27Fon+kuCVA7hvLOy4ujNkZHobOV5znLUrn1fx
dZJngRtoD4iK4LJQ/QO2TDHrYtGntYu6QeTXyaEv5YPk6ktyNR2g3HqBQ+lX
JwqcmfXJLoaKNAFOc4NqEDvBrEVkfZcHJAOISpnJqPTYFEpKKqmYMNe8vuop
BoVFuQ7NVq2+y0iw3AVrAoRcZ74Oku3X5XGZS8Vqg3CtNdvr9TtdaGK8QKKv
PZPLjrypvjfw3LIYfDlnzh2p8rugYK/7C7bUPNzD/ViD0LTEx8Wg67zIbHHf
LPVs2KWovEqEnaIQJVHBQ4XQaFEwO1LbNlJk/KiY3tdgGWUbGyRoDunSQAqd
CEtCDecQVzTUBYyMQR88rPCe5tXOeVA+fpgPOiyAHETVMS9/yBZFR43v3Dnp
ag22m/zNBqLJyyQvcRL8RQrKIoIaizCVyqXnr26FNtRk5E8qNOCKaZxQdVCd
QnBORFmH6kvQ6gzae9WY520do1uGHqgWPdyo1sj4kYLqrO6sCiWpIEVOhYnu
VZZwoL2ZHI5nfmFudMGn7ZWHW4PwB38TG53EVvY0/f7TRVSn5plqt9rV/Bsk
7sV3y9fkeLjmC/IqM71f+jx94RB1rbhrdXjFd45y1mO5j9ffX/QCNr0s6RzH
t/GLYRRftCw2pnksh3WGC6wMZIWzm2Qe/AyHzS73vqTsl+v58pU/9zWEWpvU
JE4d4pbxz5+lGC8YIL9iZSO3xdJg1JtH5m8SWfbltxEIBaiPGK7FCwktce+c
rj6P6GEWtaCnJBPZgb4GnCgjdRVk+3qzRfXV57k0dmIIxe7KkDylt8fbfTCJ
ILYQBJwFCzBVoSC2ErCHgddy9W62iFhB6JIcR01KUF6M/WOojM7KkBj2w1LD
sDdYFi2/DMBXC14rYm7pwtMSF2OG47v1HV1xFMMWL6o3LRhg0YqBLLSNY3+S
t/i4AFvn+gB9wAplyrS3Lpk5Uzj9PT9XI+DiMV+qZTE+omyF5+PV0Ls4/vIH
XL8LLE+NTMBPLZ4Me2rorDVkZ+4qa8lvYQq29Ens0PCdV2S7nE9qBaCA70hn
+9lV+bTd0PdlZtfY33YrfzZ87sd308uWk64tw44gv4UhJEF4cXr6gV/SRePb
4easWAi1THQsJl3TeW2MdAZXXYe6UvwV9yzl4SCVsRJWk6j8xYAY3iobxcya
IE6Cmnp3UZ0i7pDMB77WHCEemRLA1FxWa9lLlqBF9MASOjv/VuAdW0U5oXXz
+Ry90m979HcTzMMFjAbyRlI3UJI0Ii6iDgFn1EMT32DC3bU03jvM2DftrO+U
r9PIb986B3FqhXrwH7iR+cCFT/tRAalyuf9mV7x8LuiMxFYN6EnML6+mCtV9
RocyljcBaaz9wN8yZr/zNw3DR2s2SCModtHg3g6FPIkXv9hMRw6q+lfAxZhU
7FrqsFjMPnETzNeT6w+Pb+XPmIM5v3c8VosBGkWBsno9F/JhlPS79gqVT0RI
SoJL0UsN1pHGFzPDutRUsXaeaRjud3IVlmHolzQJEaMOGZYkDfk7c41brREz
++5HCmAlfpXHj4bI3dv6nngUgVjB60JE9nA69WwmCkX1+Teex4SK8dfs4Sv/
F7eR8+7BQr7fwcyH0mMYzn1Rqy59zbWoUgAcDzcf/Tcv2GB+78cCNj2OwzbF
cbgtdT4DePhFady3KrTyZnK6m9Ec2NS7PQmmuR++2Xra6pLpJG156Ze4/2+y
LXnTk7iQKF7BpT9w49q1kqAVtrjYZCQ2RrM8bTI4eYduHQRYQasmS3lvDVUj
4KY5YVmacSCuZsNBMEQ3zqPf7Eb10HuEMzSmwwZJJdVC69cSUGACZgTTt1Og
zWcgBsDV1jzvX+NNZXdfjDULe+kUoVzWbe7MkFSTPG+9BFFX8WKjhAvK7ir2
ucd/kL3lxGgcXf15oseaBljdIIWZqvZkzx9bYqc9s2leNgr55p4p+HF/1My3
qWJQQK8o/BWrhGSjanalRtTymmo9+pM9J8rc9XSAXW5Nh4IrIaFxdGCo+wHA
TqQlBXqbhUEEMaDzMgO+W7xRCQ6IG6ugJ9KfP3NtUZH+RKaOLIHFdCM0p50p
M19uY1g74lN1jUbrBWGUTxtLrXrmINPV7txNxQpXezi9FLoCVrPpXgJq7hqQ
nBDMJqztO+rSzlEsCDgFp8zMyJGI1aLfPWoB+UrEJ92K6pgrNMnIfM5LoPON
3fORAsHgNevS97E6DtOGRyO9KKpiCi+R/xWEv0ajyY0TSjA5PW0aZLbPuvwS
Wh/zfTgv/395qxjv5UqTGaN+Ud4VfyJaY2iXlIPgaD6ZxIdr93Ua5UXnQbqz
nWWJA/QJ3icyS+gP3Tc7ArWs5BoGvezTU/qUwhMx48g1f2YFvtF6tbLht629
MT5z26FBe/LoaxoqR9aE1lHYEppLRgGsm1hjoszc/onzUjMq8/Zp5KMVI6nO
goGbuSccixB9qYS7QmafSLyB1nKNyjMe3d9K1X0URwKG5VwfHbmGaPAdZC1E
ohyIjkeMw/2oaJg9HGmd+oy9cUZiTBbyQKX+lczwYvenKgmiULmV/xXEIOac
CsSgINM/+CaQF1zY2Ic/uOP5zoMkjiEx5dZpOprTjclhQgyWlpjNwOxFglvN
OLFOSyW9sN9kEPo/s/+LGb2oHUGmytOJ1gOVTR/YKULNfU7viq8iXZkfg5Sw
s0paF4EOecES6ESGVi7TeGDdUExxgkAfP93sSIMc2m8R7Yssg1K1eDnMyp8D
6z6m6JnYz5o8cPcbJc2YHO4GP4AEadfUm9I6Te6kAi97CuICvS2GEzOKzZvu
HOz2zWPAWnoHkE9xSdFAoFs0yyK5R4Dw3SmWktRqcQMLrlzwYG4YLZJ5lh5e
h1cn0SLuJrCMgst5QiSWS2JEhkhOxPRGAyFY35t6ovtXlDUFfKbH//cP2yX5
xLwU1LrB3/O0QTk0XNej4UAwuahu4+CeoZ3dVNR0LnaxpDyHLNw3Dz6syUlM
SGP8skFXgJJMuE1EqVJJmbrLlw22igy6bMwXvM5vmAqENlCW5HPcXgHeUuZp
So1hOHBn3Vc72NfSnfjkA6hSo2TY2pGI0+L9FAZVqwGhetbW2Po3bXyZONHO
UkA2muqmsCyblvKICRf75ARO/kc7PujMmftBDFL+bVoG6QRRdVXelcUwaEqS
aoQIxleWpObz43oig0ULS0ZYxr+PZI/hhz8v5A/KKnqcEHNQJZ57/11hsti8
FyPLskTFH3Xo4oQ0hK2THOcPtbYkIG0jGAGt/AQkikj8Qh+t720nPcM6Kny3
yFNd080VlsjxaK2D+wRycHcW90gCg0JrKa8435c4UgIaijzCMeogdr+sCoTr
7CHN0G4HFzSyreysC6H1w/b11tM3zYEzGAP5fdAibLcyL94fbFVcLBYK3DvK
iS8thIpO6PPjkr7htln6prNSxKWiFCAdTr412MlQM3H7C/WdHWRiv5Ykj9hp
rZqeS4/rdnU4xYBgSce9HMnErbe6SsY9zJe7MM17MHeD/PvDhSAfsqHCDOIU
q3+giqPmOkjLvV3gCub8JAWR8gXlqcj5TPpOyNy/7cx17ELtoqvPwuwTJ3D7
y+HiXPulh0nA9R0vqhBY7QyK91Ure6YSDB3+97J15he8b3HZV5X/qLHrwz1B
gBzVI+3CBeteKJIcxMo71tbcxLyXUIZHGfb8pckVLpAcvakgCW9qygkbUkYx
opIdt2EyQrqpjg3mQuKGKu/F9T8CU8oz8g79mdY6S3FL92VNkZYnuWVjlynJ
mhmabIqq79/muzVbe1q7ObfPLNuXPcDVy/ngIKesXqwQfabsKfK/SrrwGp2B
sV3TlC9FtEmhOVZjXVsktdgf8LDBCQFxcHvtxF1N6LQS++kw5BZp9Mj7UPtc
8TjYPTDaSCtaA3SSjkC/csttl2MIOj4GVOOBDjy1cD8p7k4SHnscPxjnv0V5
s4lY921ZZKq7lZr0FOseu8WaLvuwTOc6U3gWx0TgDbHOGcQC8W2JUGTzH1M6
JMaWPAGBHsXH76ac3INSYKpTUZXbh3rk2kLqM6E7kpYxhD2TmWaJTZTp6EQ+
ZgtLycFMofK3HKztT/UMZjG3CjJWYFtBaCKSg6PYb13drEht4ok/xKd/YfNS
HzFk6HOBhkJDQn8f31MdBrT7AhRbTjcJWq4nlQPZMl1iyA8TWbzJy2P/V2yH
40j7UZRNRReUkm2V7jU5bZvLwKW4tR0QQZlwaGYG41DlcF7kRGb6On3uJ1LT
/Dp4MTIegzhOmb+7IT7N4/Ci+bt/dVpaO2v38xUq26TE81OQxDVDKRtGHV1f
nb6/xga02/o6hUyQ0Z9lPjdJlhgSZjdum7688FHXhGAgJ9gNyts6GbOsAuzt
KRiex7CQE0Yuj0WeWjpShmdWdu+8i20L20tAj3HN52aaR6SW09863qtH9Y1X
/pVBSnc0YjveZK5L4c946NlOpbSnG3sTfD46aqDkGuoWVIfrdajQcGqvg5m9
27/BeHnLPjKKzr2lcjkWrEngYPNZ603x3eBF4jya5XgHQcEZwjG+Jt60g0ot
9vUotWAYdKzvW0h80LuBenkBBhJ4rn+ZmfJViXnxcMaCr3AWuyFYcPbOwb/+
ecwTCw2f2HVnuLcZxi9a6OThD/uK6bHjs625eUR5bKxsNzsCAz3VTdHbzkUD
4Wz2mT+ywFDpZzRaB26SrPKGlGnShvcrKvp2xu+L2qgl6UwQpteA244nOfSU
5Xxft2hd5M0oGSxZ055sqPmwsOqIg8aO2PYlMRe5eiNtRJPw5Y2ciNzovMDY
ZyZGC5GGIPoL971Xs6pTgWZRzs8ZTtiZzLwAovNcRguPtOYolb0coQgaIvhG
emrFjdAW7VmCCw3ZTesT48alOu5bfhN7y07OA/DfW3X2RD/E1h36jEMcKXc3
KZ6WAKcVlPf2httEffRJnCRh6FkvP5dMaGlIZl0FUGXOlO7hl/JFCwHQoKgL
uLZrwVbdSGhZb0Sg8iBsbikntuPOEQlY29HF3KMAraTW1Br9z3O+KBR8NDM0
XzvTEouokb4PJrbJMnhxBJAf76UabniNI26wrab4wbDSsEb18r6y6Qml84xO
++L7rrWM/ginHE/JKd2eD0F0EyWo0Jn6+qCtr/9xtjIPcE6oeheZIw+9Xv59
lyW4EnUnQ/fSnbQm1lixsSZVzkXd7ICQDULqEk/3dMYZbHxI0ILNBGxuPQHt
rtlIA9PjkuSXTja6qh6p0X18BWTQwVkFF0iEYktI7Cgm9JE9VESRFm5AruLj
+L9Ag2Lc14+m7KwixAZuMooi83dFHaLlmKawJa4YDYnFtrw4enu7UGEJ84z1
FBv7ZS/TUZxCg0mlc88vTwvljulvfwX9JXgnVnB3U2LnVTcylCkUtgZ1GgtU
uCEcdJZYaEpMGANGlusaW/Q8z0ngGrIyt894bmaoPRIFaQnFrGjtnE7M0i+C
UeXJd9PGVQ49A3mOs2E+zeZNNRq5OiUIO2TcE60AFK7V9CIMB+9xXqdWewd0
iCW6ZCkLpWih1CFkArJ6MvaBMEhBkz8m17s/4ohmdmiojIcV1xPnBdlXJbGL
TzYKAMNadhfhY/uDTz5ZbnbjnJ8vpUcyCofQxnZUJK+SoyjtVj4kgU5aKrYa
3uwPSiiV9HT9reXNYDkHS9c4QErUmcA3zdr5mY8CNNN9ZgjBT1XteDiKuRtq
PpNiuqkh55U2IzWLtOqFGfIV8uwPxEzQJJ3X2wJicbL8CVMQcClI3bQdXp/6
XB3X3PseA7mnB8laQZup/pIj1/EUdmEX5yx2ra84PoiBnde+Uo3ZSFC+EuNs
I2r2JO3CTXznLPdPRCzrAXp9RNqWTdLEhZdpwsNrlA5NBnwWXoRL72cieo88
2nWyHnEO7jbWfzfOxuFP2TidXZH6BK7DaVKplgUySUOmaps7Va9eLEpoYAVO
hwX/0TmbXbyfoLKSggRw3L8HtKD2fSE1XuEa0CATQop2AT0Bd+RfoELBl8om
h29Syl0aq+DgUbagWpfUq+zR23gJgEYS/VARlLvqQqlMJ2l9TseF1O9lMYwR
GpnS/vqzSQw7t+FHCb7wg56WI47RJ4X35FEiYQbfVeM5Nd6on9LXpD5fRnMW
jZyNwMuv3tp1FgH7iSWtaNmNiTUGUPPzJn6eZNZgN7QwvY8W049hfJ/QLdMf
TKX3KoQAQ62X6Ir1OmQlmGjaLXPxuk8Po2f9yPBi9H47nBsA45nmHEq8o1I8
fYPxMo9jGSPZ1pmdJuSudDug3MgS4L8iU5CEQ8szZ5pq5SfWT0YXJNyYM+KK
oqZQeV+NXV4ZqFLvGFsWPdobYPqxGOj1/AqJNPoDoaeBLFJz/vK3UL+IkEhV
l9L7FET5RZXCVH0Wx4K+skJ5i8spWtu3tggkh6rrWHr5azTvFFUAz6tuAyYh
99UW7RwUJmsuz5pglQyYjz9XgoAjIp3gyxiOg1r48oVUQxYbAj3oNiOx4i2X
s5YY7lUhmwCYkHDKFs0ynbelMBunpe5nlnue8r4o4sueARCcSbSLzfcXG9Vw
wKKBiHiQPvCOIkil5uDZAgRjkfZ0M0NsdjDYNgQnaRstn7PPOPPo961Okw4M
BzLZ0dYhfpyhEs0zNa5jH3zYCVuDKC4RKfaCrbzpR1pA5FpH2uq8HK1vIYtH
tTuUd/weD1qE/Oi1q7YwlaQUayui6ZLMMhRkJOd0VsO89HdNNgbMVbuEltPm
Tzg47/L7h7zpSbgDZVneEMEPA7GXV1hPnkuiuD05bmw/t83O/74uTMYZfexw
XOHXpDZfGS4lUqZPblsAvSEU1IUTjYWz8qj22MoCUCi6lVNPk7SIm/yVtNwi
CsxxqeIgWPylIHWORfrEUKMS3ag9c/FT0hqy6DpYO1q2nrX3qMB3rWJYs+lo
gu3nd9r7NurdaBmIUZLpsca1XnMxZgWzbix9JrJ1HD0vRyBcONR2QY9/Mh0O
i95JimPayfgOWwPujTCxEJU3uSauDLwKc/Wfw+HAZnxefV5CecZZwQuTyktv
RBmDp8CXg4C0A04usQ6l3R9ds1UplbZuEn32yoTUczyGmy6PbQu7RiyedvjU
vDRexHBvVJGkyLS9t0tIJ82DUr9PEPyKTWt6l6hj445mwOf8uAy6S4Wmx9KQ
1uQZ5fX/bV9XAhlKyQAlu0E0AFab1XAy4GQTivpq/uekUvrch7rBzPEhIr2q
ugKoraY5hwkHfGfqCFaf7D8ja2KHnW4RmX1ER9Mhx3Z2a348kCm3zJxEBJSc
b3JtvAjItuBHvLU8YPWqvsIfk8cee4vPO2NNoAbAnDoVV0zKUUZmr/pY9COr
JRPYRXP2FPPXHJ3zfT0M4fpe7NUNTxcs/hUYPjl2pPCeFQ8AIfi7INL3NnxZ
OVuFDjOrVZk/sgtUeczSJs1JWrC7EL6l3gplCYKK1+tVNuVtTJvhbDQOMqMQ
pGg/Bl5KldNAddXgMG3W0A8bfUYEUTHbmMouO8W1YnQJ0mgOb/m6+gZDHLEE
zKmEMRRKUgpHyIfq9j2UdQYcarmQQegOWa19EOHm7aZhNK4eTr1CR17RnRnV
I/sGbFq3EFejRGydZpAWfyXY+RuKGN/XGBkDPCEZY4xr0FJHl+sKGHjuXbzU
5jTUSpqeEjpiuG9L2UhtnUAV6MtYsGWkvkR0mw/+579K/Bsoc28gvzGEPzUI
4Y3kD+T80hIUA/6bYpk0gV5KTz/nF/IpvEuO4107brGuAGR/2JU9uq+8Psfp
JQFq6HI7KLPKzbxBHnEcIwads5BRrlMAm7/B17xWC3Uw+Cxk/7vgzPaZXD9U
ogHchCYsgJnLGR7l+8nyfapAWfdKAbB9kTFhX5ixLOuUlWHJQte1oLMtI7lR
A6dFjXE65O7tJGx4jIYSQECQoMy526fWbuh0jmUvPrgihZdb+URDHlvYaA6y
uD6ol4xoRlwoEl2BT1MDlBcBh8MY5xWEvOMaNmRgei0zG7yB/JoJZLgz4cWG
KV2IVd53HLy4O8X/phBbuGkIWntV/1A6GtRSzQgwCG2M+hFfutsx4tsqNkrA
YLh6Nc8XurE+wspXFaj+m7xfHo3wbA8JtrvZhlAQtZWgBdcj8cMczt62AeXN
InGbpWVV72XQSVezR2yTzf9JVyjYy6jcmBPwaEhU/mZsa23zHUMNS2almZgY
G/dqndKrtzHcW2LHwOVSvWVAwgYHuULGrLnInWuBwY01a+D6rCpHZVzKMCF9
LVrS4Mm44cbL0NO5GfDNhHvsg1l5F8/4l5Wj3qc+TknDriQ9CC1tZFhPeRwr
HgXU/DpwxYil1a+ZGaoFPRddkpxSO6JPOP+OmqNoEHHfQM1w4801Ad8sLM2e
sdB7Rp0PcyXX4M95xyTKJxvnwrM0CQG+1KaOUIhCC+lZSLfurlIJfXIoWFMU
M3EIgEpGtbEEI1cC+IkAslK7VjTVV5k0kMYd506p7UWn/vTp70kSxdhD9bKu
YIUdTsxakEZtnGm1ZzwaE2ePrB1wr1m6k2QO2UtEJ1PYSE7DD17n5rlRPdDS
3kVWrIBI1LsjeLtRKFbTrT5xd2Y4h3QP3zkygAEDcY8xOu8ABXd2DFKliorA
pbH6vkjNXNNfV8kmd/JuV7c3PxCpMNybxI/rI3myjBJHmY5biGo7D5pVlBIx
H0Umta1JKvw+3ulMqGFdDh0xtzB1iiGmGbxwKG5Z4LBMn+oXBoIiSUvK4FDb
sz6CBQLawdC10dAUHjMhelHXZx3Ait50ejB8u+H/+fjdIENTR2anxC5hXFf4
khnE+LeEo3NnlhTgGK4yxYTemowX7/0wnx0IYRWWlAX6pQSaiBKz6rH641eJ
4UyItitYHnB0sNy1wGoyFGVwCBl4sTGqTOcen8hApBIWT/HeZuR49vpnI9FI
jCgqrECvmSxB1tqxrwUmBQeq/NfjDkFuLa8C5V/m1ipOPzFmDYK8hKNu60KN
FWtkI698+cBKKW/HYNEpZCY0ZEuuGlBBtmwkqieULwNwtaG1Vogw0GLd0pq5
4FOeUqAlKbISUZ/AmznQe4UkipEU0YW8vBvL8rW2gk+98nCD+vYmgfMpnhui
PwoNmSdWvpZFMklNWWDgvjSFHlUWLMvsfKWvqyCAqRTyO4sDiDYlLryZJZer
Upo4fVB0MEVZpS/dpfYGrS4XZNou7FjliogSKIYZsbzWLI0gSfR3XrpyCRlL
zn7uSFiGJXNk5EiiE7exmdmInE0ROS3Dc6UJeie7Jw6t/vlsLI/VxA342txk
sqJfrOenQ3cMxwawXDX3cnqUCl2+jva7uaf8rAg06UPhPVPDQNYVO2G+9ppA
OJ1FcRRTOrWb9F1j+F9rKdLRGkb7ljT1DAke3v2ABMECLKNBC1ocgMExKs3p
N7VZfhAOlBPeFV/0vdaPXipNF2ZzFEwiCg7UjjQNzsNlcTjfZVQBqJMF/v5I
cBorI3eUlpco0jeWU3bEupiOvJuzXpwVb6HwgldkxVYggEq5mBju9JcEXHI0
ay9Bc+R5a+aZYKescQ0egQUxMP2FSKWks3rNWKqURbF3D3HwtQmiZDssatr6
YEc1H8wawSWOcwmS3FJfZrRvz3FqFhcC/u+m0U513IOrCgF7bv2sR900hoEz
CI4D1HZia4ELC7MH+wPpVPb2q+MarNfGE54jcYnI9dJIq3yWqopCvj5A9Yqs
GKbPRCP3MZD8X47x5VJox6PTtlzIC6DSZ0PrTpYCxqTtZZY3nzlZvn3BGifI
GdWYoCUJ2fV98E3hj2giiM5HorNltUrPYAPwKlEoLbYUdob/mg22a24NYFa9
PeAiVhPFS4EczXRDsjyD3VwZ+Tn6tjYYyPsqe0V9SL4CVVsOm3Q6POKSgu/J
lgs61VtChk3mzmyOQXcCEHREgK99zpK2DcfGlN3gHQg6ktcqc+5U2d5lPkGK
AK4Wf8yJqVxvZCOkCMVQ+UMEaUy+vD3MzDGU8/NiJsJOY90JX/i/T7Th/PzN
4i3U0rTHklY3tu+kbztuOfTebPBemME7J5l/VVFLiwZdGvrUzef+S+cYk/zX
vgtkU8Z5121vJAADEk5UNK2OiAyRKqbVCFh/iXyinyu4rOPZ+xwMEZYvore6
z/5PcWZgB6KGr8A3wrg4fFC9icwXxSJrU0b+ixSLanhQtBWpOkEXSG0ZdkmJ
gVQnBVIMWaOxB2Kgne3rvgFeC0hBInD7MXGqOj9FDsFtnTWHaN1AG38XXLhG
YZbVEQPMUdCM7UL3Zeky3F6r7e7kQL/mA4Dlrl8wPfqeGluiP9C9HMhruxdd
iJUWxgwtDdXLQic0I4aF6W/CDrjPBO4S6MU0vLjRj8h71ErMbXAEr8LcZb8C
KGcvjM6pmBFc8ONCkKfdBvFNLZSmh0JMs8JQ2LKUoWyltJxYeNNZ0esP03Kj
WY9KH6m2iY5BZiqE5Fn2mki9NWq9sjuJn+XNOUjvg6j8NVBkV8TF6MF4nMOb
wlMQyiDyDTstTZtuZC4ExhFR9c1McOodlR4OqhmmsRXv0Bl+qPLkliiaZrMd
HqnKUVDdoyijFmwqUVy7gi1iK0TG06WkLv2BMvBppnuhILzwLISAnl6Hx1AE
qUs42WD+SuJLy6DQ1UbASnQSQM6u4t53T6xHYe2YJ+o9PC8AhDOgYWXjR5Y7
p1vZcxPzOmj10VOwfHsZsECerverGUeEUXsKEniHmLVOMt/3QZr1l2804YJL
6DGdcuurs8nqPrLgb1Hfwwz+7KmrRA8qrxc0RExFIMgM0LQZHJekb9xdbZ4N
LwPnjk7mOIWXjWs3a9JBySpaT0lOlDmNnaKwc/qzWzSMrq++RT9Ie7XwfxFa
mixrttJ6stl5XZPba5b8JehCICdDcihUnXJ20VwYwHqe3hAPm5yJ/3mHJJvU
RLpS3MGd2xv5pxwHOFmg/W2VEHvCVKcm3NcN1NHyNTRjPUTqpRzv0YPdo3LP
TLByKHgnT6y5CA+GY4ao75VRRewg4bvkKnToePIumwsvGufhGjsD48eyGs9F
PMAPmwxXDEJ3/Pj3prvBn68zxOmui5i8VeqZrnKGEPoOAs3F2tjy1fyVZlYB
rqYjpcpPZgb6kukbXi0+DddtZ1wwnBgTfC05z6n+vwdUVbxcIBrQDYqJ3Wpu
Q357mjSoYlcExUHs7ySBItnASkGAJy1xBVS0BilyPWhlMwf7ysVzVvyudZB0
u/DAfXWjGW5t4x4fCq11+L8NbEnOBqAz3b+oqPQf6nMyV5nWFdstZoHs9Q+q
w8JNPmP1X9um4GCXjzrDMG5DdsK2g1eaq8J2D+QhmhP9phHtC2tcNA9IzHnB
T1dy/F1wNPZNYimfhBoouSALhvQVgRBUig0Y0LnkiNMg2ycpOdrylkloFQoP
4Cm0rq5I6vRvAU61owp0/jYar0GckzjBHv5W/dle4EfcbZlZ3tTJcIw8heO0
U/pczTdBsTekZAdoF3z+o3jWlEQivRZNvpFbeU2SDaFX0t3r8inBX4HEQ8w+
XdZ68qLm30FGSAVeKKRJM8rwUV/gFzzeo8QpYjX7TJjZL75pbYmhEhpn0SB2
2XAxX5P5I3OsA5xQDTfbyNPBjE/yZ1vDzBCteaAVSm4M5Fu2Ezi6cYoEF2la
3iZrWCo2K9xS6DC3plP2WdQmieMtbgq5H9eNXvuj3LumSlsmA855qbtNkJJf
NJT7GoBCcjoXsipS/liH4SVBfvGPTU/s5/dHVNQRS1DhSAdMyPSGQxB1pBgf
rsrU/8jfJ64XRiMWZvJ4ySnzCMdwOUYiE0v+koOcSTusSlFsm240rY/XWDzS
B32meW5/oYwebKAj0Gj3gzPMl5M3svHp0WBk3fbeWJui50asBYE4YqQb7/F7
zOHIUypnQlNcmT97iN+CBqFimY/gtYemgjT+dOJWu+PJtU0C+v6HzhAV3kYb
0XgclTOckujghTBqtxj/1EV8ELarecIR2nirGdUfTfPccDsqNoZxrVD32Ok0
IHtSS/oohsabSD+m+dv2OfUjJ5vpxoTHiYU4RYbixxiceeC7zIZz6UuDfMRT
JxeVyFGbkmuskniXf3+3psaO/7OBpDMWImHIuN42BovuvTF3irS0cwKTlmHg
c98jXhFC2guXY5+sVaMmLGY7mhjOpxwMHQy3bs4B1FC0G0IEppA8gvPXrU22
WYw+RIII0GVvkqLL98YGZRmtPI42YHAfCXspTopcYamqM2JuELWwcZMKwJ/k
sI5Fy1qS4JtR+HMjT/OUWGFa+dBbLeEc8d2OeAu8SM6XqjRV2T1jiCywRukh
Jv9Ytns9EgyFo4V4fk/xP223IsGvhAFlV+Y366FdrB4is2ck5+pVnIoZIm9d
X1uQZwU/1tJ33FhchTvSjI+J6MsdEWhRnFlP4eBGIV6uzx9Wm9GU5WcaUd9T
A+lwc+bpjOjiQjT4o8Ox60xUa2KmCi0k5/yTE/o0yYts4jZyBz1guDWRw1u8
pU0+hzW/TuFI3GbcYAEljrEVJBAoaR4EY9nERs0ardTkqU/cOJqc2PaTY/is
ohkVaPR7LrmkkY32zOYky/NhKyYSpTbgNa1ww+6Jpwr04KcfmLkm9Hoav/23
TNaAyMHyBVlMRitP83MUOUHTyq6HSxGvnbqnwhAgOjtMxfOzO9vW7sFmaJGJ
zQBwaBFeY5DDBePzk/37bifLHCyhObdYkQTxF1FRbXIYDSuXH4e7BGLZ2Gsn
A8E7G/8/qZ8U7qSlHtIirjHsiQCGNAMGagOdtKYLDEwWj+CbSTt/085YGXnC
iphYnQrZwAqOBy5Mr0M3mBDyG25dBOWdtVpdPeAilngEslW8DquhBji2XcTT
NRNCCNs1YWlOQXl7zlfnFtjdDtLnOHR+4gDmJ2m3wV+BvTAADVwlGjbJKDOD
4PW5aNXE/ErpvKZcJ4DbpJ/ym+a0dnh0+cq1XtN80iMqqBhyvMTkCFFzozIn
ovc89eTBB4lt9DKiYEKOPEggsYXLcNNFe/QKuPa8CVldwIaabQCDHR/PmlxC
Gop38lAzPDN/tlnf9WyJFJUPkWWsk1ZjFUI/bPam0qjBNECooh1MMppNKX34
zUvyFgkE+IdYs/2Dk1RO2yqyCz1O71kXz1f/BIbStvf1Tn/dxMLeYWsVAyn2
n5GUznoNvbQsPbMK0bqRsURcEg4zmn9qk+UYbYwf6M8biHXcnWEeGCyU59ix
HbHTKepmHwbQtLoAd9CYIVeOR1w/9KGPAeTes1fjN2F4WeOE7MjR9D9OaEJO
ZucIshL64heSIKWXEchFDHTZhrbTRJQFP3twFoiJjwnLiGtElqHmKcaxJEba
HtMr5fWHVFpSXLM3UcatYgIWfT0jFa3iYol7fjuj5mOXPwUG9Do4QYTWMllw
MPxImZ1wjk/5DMGbl94n2iyVogKhsxWWBjn6IEyHH5oNMMrvoe0N+2LblDu+
BL7Bb2k3lyPn/AtU09Q6FGBQ8sjim7kBv5/53nTfNFgBiAhRGSUwwx0ap9fn
2dqoKTUbRCFzel3WRHWf5sYVWZHMGia7LbOSRXMQZseQEL0DjKF0J+Uj1WF2
UwGk9fdYjzBEDgbAUXP7HraQKAl7e516mnNDYSZ0T8ihMecXCKKya1/0h2KG
77GMtJfN3PKNRok5BkNhweX11vbvplkZMqm1gxz4nbXe6DKMnsTJk+wceBQv
V897ZVFcHfJHrZtzolts5/3KK9ch62vcCsJAHzYrOvJm5PWBDcQpfWE6B8cL
IYj9tCDhqAIfLQut1Q8APRrGUrH2BMmq3KLcpe4K3In25XlN9O753FWjM5Fh
8eYXsqytXxvINHDv2e5A7OBS2mH9R3/8SW2NH6gvwCka4wzWbocJKhNiKyec
kck5NYOFf0AVRaZsWA/sZ23vPJNCanjlAid41ulkUX1BxDbDRAlmeBjip0X9
GiYDlw2XFcoeMETDhgb7eY3yLMo6wlFB6QSP2YZWdl4tdJTs721RttB4ToKS
+wJpQBAbud3jji4GXWP/0vvGjF9lNeK/nu4TMDqctVm8tEjrbdczbMupKvfb
TPARIRA0O3ZEesqpwVkZAwOWxK7AIAHrRM4cymBAvmORi6P2tab9tCs/br4A
qimdlZCHj8FRn6SNqBLdCiKG+3wH7Jb455576jnZuXSI5x1aPrggFlTqdwwO
iwiPMM3pbQRb+iN8dGVMhHANDN9RdGfKk/azxvSlf54HFeym+o38HYSzAn4w
qzG6y33MljOsXnHBcLcX+zFU3E9USfjvbZsTEgtNEUXJwOE1Tjg4kpTMcjKV
OK5kyfg3xFIjReWm2fqlrCXJuKFgGPzqaUoPeijBHt8ObCv2i0rx9dvUdlgJ
4NmsFK4r0xhYppuv4TWDueH2h15q4AA2xzKUlLAhQrAB3Q/u+39lpR7vFpEL
vGrs2c751UOH/AUJpRRX47mJicKYSEhn+HfWZH8pHcOSA8i1jdRSkeZbxnU7
IIhSfcICoPKgcRsgH0FjZgyGAUXGD6PXorfaw2xvdU3vsJzPDIJwHBDYvhBW
Dep2b6/NMhC9hUyWuASDXZnpoThz3/q3UTUmnwfL3iqJGhqnODg9gSwvZ42h
TpYU70ERZVb7DkYGRm9NZt+QDb5WymBTcso1GQlqHlApk9qwAoSnJFibf/7g
njsijNNXIghfm2GTNORLBC44l+8DEVKpaFaLYhy8Vqu1Jv957ymGZwDask9f
oymOl7bsbugO48duszsZ3NqdB8YE0xWrafT4qQTcU7ytz2MQzsHU7AsxxqDu
Tk1jLkb05an0eLaswjzBzTEIFOfXHLtPwOoXDQJzAzlDvsnrpXOECJPb33/k
oEuIT46BodpWILWG9TrHDIPj88m32RCizQtxH5O0x3B1Pw/Cve8301Um9WsL
rW7n/+xYA9lgug/CDKfai5GD8F6w+GCopsfx5F7+JQXLXy3PoziM7KfhFggV
UBiv78yQKFcQ17B681fInvFx1/lO5GSODIPqdii04tAQuXmixK+FsvYgf5GF
bnWrWil9xuKht+r2pYRtWQjZvChoOeVJ2TDYB6ssEfUPtgYTOjlr0dMxLxrn
pOExzBnDlv09DppoFLtPIxWEadvwv7Aye/v4YYrEiSZtz23Sjy6BjNR5Q68x
G4bO3OpMXhWUJ7OmFhuY6iP3uxK3S7pHxxkWaXsMwbDPzeW9y1HBUoAeobsd
QJ1UTgQ5vB6ACvPawdS7Y36ohNiy1EOsIkJcWEf75OLM6lsQ2KXLOiZnkXPV
SZ8nCtqUr7g3wQ4t3Fez4SKAQiMC8QkY3pstM6Yfz023ZjvUuqf2Pwi2XkKo
rEiZiwwMneGyOtwY6hE5+vWsiSkOMbQiq8mH6Jd7b8jnS3GeQA7cf7yRG44W
bK0ksWCpU5YVsDqeg2SJq7FxYZPJZz2IeoqapCk0LUUzyc2JODceAmfp0KoC
JSu0Q/PWEAD+bidqvgK6u7iA/Rwz3JxMxdeaoMC27gYpZx4cKddmQE7C0Gar
jhCMJCxFR26gqtvC+5CnQkgCJZ+SajzvpmEiJXryQK/oVd2Wb45xonFH4iGo
negr6xIJWVMqY6awTmicVK8gYDANZES8wO6l+lQh56vIQQ2muuuiQR+z5M7V
jbvpvQwcGGS/Gd3OwsqvS0YjKgENXWRx+so3EZHCppM1mAkk+fqnGTQf4F6j
fhU7Gsq4kRY/db9PEoK9ahTypH+MOv2ODy2EJV4j8PXHn2Zk+4iuwoNRLC1h
lMzHmtt07QMAoDLN6xihz4WizScMg6XyYYr4Ajww2CWa76NxaLqZA6sxi0SD
rtsO1R35DGCtdcQR/rZ9sd6sCLe/t1l7pyORKv5nmSG+DeNz2trY6+KQfK3C
tybfgk1+CniAVI/emtvOZ9//2qozPycHxHl1fRHCukro9N29BRTNeoZVP1+N
YzHPD41cUROqBX0OnMkTTBAepafeBD3ztAz1exhzwglvZYcSEmtlYo4F8+BC
bqecnktCpPyJF4HyFyN9Zx6FXjS6dqWovRczBcjeqJr3sRdyUI6DlGMrNofM
5TKi1hA3ysOtiGwgMCDiVfuD394tWKArN5uSlUM8Pb+8mYKxoQEzcjH92vTH
3N+HpP/iNcEu80HjkwyZY9Hktu+5OaDxyEfesVyZYFGh5kROwG7Ez5Zuoe9Q
1if+VJ+cNZjvnGvRNl+yhm2pKBD+HfRp9tAAgGdW+LauXrm1w3OVncVrq9d6
2v3BhFud1rXoxvtzlJ61g5SDRjDdOhcHrWrzmzgKrzEYzJQuwEgsu5cH6IAM
Bha39cu1UU0LcYkaptq9dgP8x6fAXUxAf/TwkToom/AZd65z/2XvszeIvjKM
ECVgA/nuOAUO1KetbExMEp9cA7DWCLdqLCx2WWkBch0cQQCvCtYIS0o45zMk
BUMUuedpEwQgBkunbAWEka5H7RwfVysZ8zUL5YXNnvNYRAsuhPrsEpJw3BDu
oZWJUWMDu1O0+sGagmJ33FnaBH3wuCp31WjsSN0XVBZq2zSD02P4NdLdy9gO
UUl+ljhG17MSKsznS/Iv3pPw+SPjk450MrR1j8DRBg2UCBfc5gJDbCi6nQrh
FAXS6ah/pNrzrRbJNSt01tTZFKF1DAa9IiW6wE9XpjV+nMCyPFYH2aY7VbiD
SmOpbdqOFXHX6aLjqphFmk0OtBTLphK/pJ5YXphXIjZrI/KOA81QV/i46zNa
qPs/EmPTggQ7RIBawF4MXf3vLDl4O8KD9BP++rXN7yqctK6cWBnOEjTxHHCT
W7a82M0AcGRQ0P41zizZrcLddRo2JoJv43FMYbmbSdhoSIchPnPi5EYqKLPs
Zt7NgX/mR93beIMG/4ovhqPC2lHVMnC2YaibqhFnzo6p+i9f6cXJaXYJTsqH
eA2JZS+AWfdibvVeLk7JpMNsslmRup6P6CqXfp7g02dHong3ggDRyO6+Txm0
sTedb4lZmOCOpReU6Q04P53FpxXq6GD+URVU+v0UAo7f0SaMF7D3iPTOkkKH
5rWCdJLZ3YmGxB68+QlAiej8XFNlZ1NKHgYyvl6zoY7bqr48h158XnCc5Fko
PgaRTm9KPhBkTg7Z1eEGR2DQEarzeZNXcw4tsRX1ksizWU5LXpLFkZ+eWoY4
S/jvT2+Lvbb6o1uwMZmg4j/S1mMvMfrs4lYKB642H7zICdNFvNKqFcIeQ4G0
Ul8KkfCCEBGSnKvn2ciJw7LaXAqdzK3E+gHDQDueT3afxmwhqM1fFukZNrGd
bz8G4VVeweWKXN44cW6mDg/ORy0uP6KaCthP1qOhWzUPs/1bD61XFGGLPP5Y
IrZgcMIMiTmatdW7f45i4EHduXim8JRu+dYPw6eU2yBmBU4QE67zkgVpjO4a
yoQFMJt1+fr0cJ/JjpkfjGWIdAak/JGTHSvj7AX0jPCNPUDw76xEqPl/OYiB
T38vyU5wpQKtJETiPizVUIwbEHBm5ZhsJXf8EqUAJlcYmMM9bh3T3Ddmii0a
zjFQt2DFxq8b9zhZSbbw9mAEnTLaRmkMrGh7hH9IOwGs4Zv4N6+5kBF7tKX1
76fqVd/FyhP62F7fdaTCndbcyMe85hPkLO/Sv1oz/A8/aX4NzXpdVKv/Rn0v
wEzA93GOu2ocr6b4uLY5050c34YJxQFlLG2iiM+kmH/VmQ6731d8u1zT5gf1
/gflZ8G1VvnHSSfnC0QDbAbTBPdwbpsruTbJz8zDZtzAecAkQTGNjTdrwEaX
UB10YndqUu4gsrgD7wFELlAT0L0pIydT2yqhlh2qkRSRqPVrn5LCjiRFW/8V
ri7eIhBvGvSCUwfNGsoI4Ap04hs6pn7XlQgEUURq1GB0QzdiAJCufFTjBqU9
dbtFR0MADiilwDvWFHAYtwracQWXq95gw8bEJqmeSto5JWoO3XdDMRjIP/mA
8A0ZWwJ8GQ8hJNalV3K8aAyDzmJB0Xx1A/vl+OMImFbFN7lX1fDg6CrmisJt
KvqjD+CEKkA+7HAeWe0BmDkOyMEXqGaxEP1p/g5RhZ1XqMz5VAMWxpaRS+u9
M+jemEf/vIojaIjjla4IWdY4lULFpU8gflAlEIMWHqseY9H/IqxK7O1IEfVl
Jw7cZe/sEk9Usz/45wNlOOfwEB0xmBgyAm0/6Wm28NA497AV+xNwjyDfhOTK
kd3phs/wTBy/tfk5kVdw4FSEO+hGrZ7wOSNOOBQiqXE33pbFWSpV9n05pZT7
i6Ty82n+GdpfDmQj9ucPYGXSKDVa2VqJir/RMdmbZtzIRDQQO5AIXZ/Jojts
hhrK4FT7HezqqI9az2BNmHkEbIPQysVR+vCNWUiq1DHQGHo9Azh7R5wFDkyU
CJLOvrX0wONrk7fpa0KNrbO0caHY6bnQHqy7o1iYnjeO5j3Zy3lNEW0M0uPV
xgxTuk/1Ii955qsk/zjXsvIH+lR9gt0GvTT6mRjEglE8YkUmi3cTw+KXkaIp
GRVpY1FPlBGVjrxkJfoG6ezpmKDBg4Kb6ZE4C46SUbQKpjU0MuK64Of41B+u
oKxX8RCiliZVIdjatPq8rk/+HtIKrMPSN3nttZtDiEJrgEG6/5nhIL3L02/L
K+Ulq/YME2RYvjT83rewfVkixi2jYo3iorGdH9niIRrM+yW7rixKN1PdM2zZ
2GLtOSXagCKkqnYOYanW1WOYuPKscyU+42VaF6xuV07+W+Vx04vYLzawckwy
vYXw7dZOqM3KjBVkov/Z+uKGYuBRuE9xK5IftCt4Kd+Bn2zJQxL1510B80o+
Oz9O1UnKdJQnKzKul1+d3UEj706WOaTEyBG+hPR0sSIHJ8RouUHLhhqRToSc
wxWzTNeRBXdONG36dRreHpLZ6SHHE5zI69AzLgGjXKkKp+I3rryZOY22jtev
Q1PhlETIaQBRCv7etKOiXUMloNo7ys3V+WiF57sTj+ob41Ayyjn9k1r9JWqM
8/GMQWe8vuikjsuMeC4qSOcKy9uRaHL/nkNJqNnLqNSOd2eq3y1SUS3XlfzV
fLVsnt7o83KFPGLUsOz1NYwvK1OaQK6W4FXs9lBUj/gWR0mVG0Zw1OYMOIXH
ghyrPqSWV7FM0b/HvGXdRSJxW/IVpzAUWLFOvGiASHAiETbaNqgQcDeui9Xa
jkFjxhxt6Kvta/irUVq6eMZI8YojgPWYkYDRmcathxbGOSnq383U3tvMkU+J
UjZk9NvisEC8CKuz7ouf6G6jcp0rYvGXVDomwfnbDNPesVyOQEbn86ZL9RBb
8vA5KDaCEvCv2+0FHdGM7VglbFC56QwtX6mwhm3MVDhCPRvbF8ViMlvkHyG/
MYrrNRGuWH2uznu3rKFj8Y6LozUAegPu+f02wyCaAIHfkVpAdjY62c2cz856
VG8trRKBQyXkRd57phLUp6SxwqG9TwEfQQ/+xNVmYfGpJA+uwwE/WXxyti1b
0+dQVp1HYJsji3MsV7F8bYdP02M44Mz/VDWqt3BfXfGyDk51pZYSeiGgmRnD
7gwG33mqtW3VfNZAroqeJadyULgRqJ4ldSZHzkRQbcu8XwLGcqykGT33yuox
PkGnl2OBz+6PIRaN66mQ+WX0YQq/H/q7/O/OSVbcCDx1A2eifmxWHYfEC402
TSQOHmJeZSkSxW+QP+bUvIKIvXoAZV8TiCEx4mC/84h1CmdzCerp9Ekpq6vw
Hgq5NyYSWmWMall/GZVEAUvTgtbVZOdN76DFiqfRsO+d0xXIwgVu5Q2OJ1Gu
Jflc1W/u/cFZiAH5777XSpPoEkyaH7oj3Eyzsek+N7z4In2W6rUbN3C7mFDs
oDXDuXcQ6H67hc9uw/Il1Rd66rHTiCVcptUSfNhO7mypGT1yCp3QSgqGK6GD
2hMkNqmLLp00VOPfDtme7fGQgKPd4KJzTdMUlnQvutY1MpLGTIX4v+g5GIxF
YrVDNm3Ejowec+GNvcdtX1UQCnbHFvyB0GCG+JVSpcwhGbVZpBMnBn5g0Ptm
uZGe2TzQZSdLIgmCv8gJw7tUi1F/98ea98Je4JgkraM1O3UYU0VLUnR7r2+2
J+0J05be8A82ptyMlh08cwWdgP8071twLKIrnjhtlscGPm6+hGinq1OlBr2D
4me3Y7b3WHugX874YuCmF6cbeAi7lrLhGXfxTH+J0mgf6PFNl0fl3/kcoREW
0d96+9ch2CAsi9WEhFM3/rQ0Z6thoPp8VaKu3EMAl4MSHNiqinS0pKkKsmUz
UrCRUl+Hot828P+U6sqywpTZaf+2+TqbkjdCh22rh3G2ROUaRJaXXj+IiCFy
OxkGqwaetYgCqIePkKBZORgG5NlRPP9B12TBPdWbRVVe3Naq0VQDjUc4/4wd
kFh/BeXaqOpreVl0xb1HLFKedQyS8P1A9T5vNhl34+mEFvFriTcuFH9NRTuS
jrkAPcK4fd8OPaFDXl70VFWIju1O1nCMFuA0st/2NpI7gBByO6P+VUiRNz9k
py/hLJ5MILlWXQcLzedAY+24MGn0RVmciMWRRRbamixZysa6TSrrZiD7Rb/g
FtASp6djCfU8jllWQteCNbU6zDgFo58DvMRgQCUELNBoNlIktgO3i10lQC+2
2NVNSfyDcllScHm/nZzkTdO5wq0q6L2uoNXNG6bjiYwWK9I2jqYGv6NOZSYG
cKTNRMbkmuA+pAzfPLOR+YDtY23C2epzmpia+RJ6GsgmcgQamb0SXku/oHL7
JnTQgpniPqxkPSpDxgUhG2wFh2sJhKSMykh41s4YDZ6FVOOkuxa13e1G7eQa
7erAk2JWpRHyv3H+hXLaUH8uVdes1c4hS4Kg7EuzEKNYLP02rzOmhOb6p03R
4COguYDVfPDUPc71kqlLnp7tAqpBV2KZmNWEUjpgsAIlOLMUcQBbMTKUL08K
bKwkyc3XZ0ZvLaTEVhI3zTJ1BeGKUIy6iqRPEw6iGF4jHrqewVowyYqihJXI
wweC85L6PRUvnpUkyB2h4rNxZN2lDakqAyrKSOf2482JN+Klfv3hm48s70wW
5jUzu8I5SxqR89KtyO2dBsqr4ozn/3GW1NW/lmKwz9ui9E+t5ngXxGsOYX0A
BlmBcl7C1quKDaxmDAoR9CK/ujDmWtrOo+hOEPqC9MNZQCJkoXte1LzJV4G/
062gqDn+vGgVS6MVR5rysEtkZP+g+bWcvO+XCHBnyzUaJbEDU8i3FNFK98ZN
wSBkW7ho4yrky7LaPwteQAv3SUiSezCyvUx7D5bCmFrcSQdjr4NCX5vYX5fW
tYPsmzWqHprG6FFRgaq+/sQxRdSjKPQ2aJGIxfu0/uPWNbvXYbi03zO+20qA
dVdLm5mNfBmRdTZ+tHHg3R61CfdQ/YM2tRLvu16PumbVWM3Rg6Tb2WeI4+BX
lLRQm73mWrq7TPAMLPUNwCjYkMtdCi/aMoiz3P63tyH7OpjcxgRsaB2MAzER
Ugc2gBoijCnc5dkNV2LpzxRK/g0puOx9k1xdrvjHpzL3hUiOrMixsgR1ZpUH
BSOfnnKLNUcUHzyDyLrp1+Zwfvx6RWD+67uITeonAN93JbXj52pVUpMAjooI
9VVo9f1zzFQdKufrzAwnwzmQulKaHc+gD86ST8lwqSvPIuqPHCI4C+DgPA3Z
XBK5HVCxuDICFTSumhIi1XcCq1eV25udYqA4EuHGpnqAz9yMk4qxZZbzfk67
nERPCh/pkAlZU1Zl6pOl/9JnMiTZ6RPESptnipDsRxfO8SoOS3LUMaTCDaUw
ym3GqMxw8mptkzGelyHKqMrg7MKHuNAmgvRQgAsxhAh7Am4L/U9S3wzj8RIq
86IDGGlXG558GNoyDjxKMGf7vYfrDxSVARwsYND0lujVJEbrrtZAC5TRKfEz
Agh2hbcf/EPgy4obA98Doj1zR2yO7m92EUx6rZoU+iCF2QPdXsyUqusQU4US
QgRBkcLnk90pIwIBAZDA0xSv9N6FOGfNy2bZHrMd48WBxMmzUa/WkG6BxBei
SisQ3kiy1iXqaIHstK0AQxeeMHQKDsoLVTfWQxctf/uFm3oHATSnBP0/PWhk
TTyxffh/0y7f4yKhHKFZXaAQtagwvLoNEm5ODP2+VsynUgo5XNbjqsvQ0ASr
lqO1E+P7XrHA39BUGmGcpPBoIZMdlebVpD/g3AduUb116amlxvgmFABgt0BN
tGjqMDqhbeD4cDh04iKOHm92yDO3LVCdzrt9kaPtqdxtsV9oBUKomEGQq4W4
Zcgw9LH5O/YCCJZ8e4uskLndh/tdIAE14WALD6Gtn26riWWkVXskeIWfRmDS
14i7XiFBh0nAA2e6YlaEzh9XhPF85QtvW5ENbKgwr9AswkQVDcSEg03aIWPW
rZqgsRlmtOFhDaHQ6busRo8UED1L6y+mp6LxTIo3Iq1sCek49E99s0E6iG6D
TSd3iXNasMn7lCTxPkejAAImdwDeFV9P2kdAep4C4WuaW2UZGlHnRwGgig5Z
EpR6EniTuIpoyCUUUnZB/Iy5TdR22n1b8WnFpwmCpncn05dEwQSsQaNkCyIC
9hl4xXzgTMZMgvm80KxME6PT3NUH654HEm+9oW8hGGPwfZuOMIoSenOWUwcS
gRZGy7fWwsv6R/Z0Ww3nO7PZpcK2X3ol3AKzxVywsxSQ2b3cv9CllY26vDA1
qyUrdnzswycTKDd6zQceO0wrrd5OV19z8x2PMVGY66cylDOnpXS51KZTtLGX
NA2vROelpwVvgO5YW0FLTW3RG1ehlo3HdCQVt6AucgaWSSv0byKjWNWAuht5
mA5O2J4llVB6qiyJBZupEWXR396lIQQHhye1DHeo7DCj3ZxXRvx2m7v+qsCU
grulbpVKBIoZlN9TNtLedAAVMPcP0Q/NmnV+MQi35f/qaPoQC/YR108IEpo8
/OOT9igjmAUSP8UeijImqL1gSf7ejA0VPC3kbFUWZ8aToED9+NrNUY4hr2eK
reyRU9srGw9Hlit1YSacrYuAr4PDcRup+6HfVT62qiwPzO2OlJBNnpwoa4bm
dV2GQFXUf1d2WCoSdE9Tv5140lNTZFHaVoDB3suhw0+pcS/cf4+08Qntpm9p
B5qI31J3zl/jz3KfweENBRLOVXiv+46LWdZ/OpgIgcWh7dS3AOTm2O/1piLi
da6+KOT3YvXe3C5UTQ7LQ2B4fDaNxFKlaDTohwCD0JDNTthvlwSDoPorNPP/
xiCSjC5sqPuGGWM7qkCro71UTmnYHof/CmppLdD2cYM8n1Gld5i3W+jy0cVj
o7wlVv2c55PPOtudMCu/uS+vw/AQgBzpKWekN5ci8GLvhbae2sfnqfP9wE+Z
ATJjSwz0JiJOVBfxSuIl9kCPSDQOhdZgmyMRqdBwNC2soulEL5wnhoVRXwWv
3Ax5rVJA2EmpK/N1mag3zl4cAQdAGgLcATv101XgSfWtr0iN/v6g/BD4aeZT
pmQIlCxYhxTJ6JS4A4gAo+nYlKZ4CDX/onkhxkA2gGtKGlnJ2hkA/d/rVNXu
xLm3TW4/yU7O0pqX9iEZSL0sZfzVijDY3j9Ac+4hIDFS56ZobQrREAJFs61d
GfoNENdZ/3Y7pdzTrtORJdxSYizqXPQ14e0pJTLiB0/ya6Cm6sXE5hVFfFWc
tN0dZmIWa5/Hls2lx4D+Xsw8542Xf2htc63rd8CjQQkGOqx6C1xOZDqS43A6
E82QxFZd2bFnkyN4ToSmk+rRK+S+2KLfOTdfe8tS5NqfyAYOjICJUhatCoBj
U+dKvjj+P7Nj4P1FZgz6JBKlawYboYMM+Rtn+sZJ/D9QtjeIxH7TIoVOnDyv
Y3THJUW4Ht565xY9PI6ePJjlyN6SO1jErPNEIEaN9reMsUgBPg3wgKz/Iu7D
buvmrYbwa3A1490YSEVXypjocliWJvW/s663KjrZ7hwcQEqHhq3Z+F6fl/C4
R/2EcuJ+HufpG1UO+OsGGPHbe9dywXlJwGBSs0yCJChlepht0+ee5k5/SNNO
uax7YtYJaiH5pNRA9ZrqWozpjK65Mqjl9B15zCJ9xc0/G+uEBKI9FJlI4xV6
sP2Vwt+VHmb6Mio4Hr/zOwfFzyX+nYQyZusvkuwlRzDGjEeJ2FhDCsKmTyDC
XnkKj2gE7GDjT0qMiLcNpNxPOQ6ZrGUNUDsLoqJpkgJlR/tCrAqzMvJMpplH
cYGtJ7yTczpPHUcrL4xhRHZc4zYjY3aNMWWPiSNQW5rrCcj5ReCANiuRl1WE
NeTc+7/IKNU7wNh7z80RH2vd4I6TgO56JXkX8W+4+b28ouITSayPV6fEt4zd
Cegc97ASowoVO+DlbaerAbfVcIRzWXWtpuX+3h/F9z9TCSdNT/JZIuofRcXJ
NGqu6iTsFyGetqB6lZ7zFpITyfr2OpHoE9mfpvjVEF7fGmGqeLB+B/Mv8PWX
iTZGPzgAlIIqQPpgGIOSlp9LySv+0IXudfiPIDec53ZNJjst2yNYYZAMqG5g
ihnrkS/zI9c/SiG/8OWGb+NUU0ZWOlagWWKuzQhaED0Gs4cfnEhazGyEfaJg
TlF9GClE9KkQj4w1GtHy07uIMgWTXosaDyYlfcB5W7u08fHWJiSJcC/DECK4
SCFXGUpGOCAGj9MBGEQNiEMAOxJE8ouRJzGZRjkRi/6SU8/BgDnISziLphnv
EMt36Xi0fu66ZoFcPFDIILjDwkaW8i9chjwL2JG831CJEYdDUaPz83pdTEiD
fb6hZy+bCA4gO8bcWfmZUVrF1lPT/YAu0Hb0PFM4Z1GCqhhVJnn5WEqeHuP/
pproImo99luWgDX4BI0HMzYDwfLprWdMHGB8RbU8GEzr3LLdovso84EQi5Gf
g6QqwqQ0PfrKsvDvodE5Eh19gyfjdssFK/Whv3idooJMM+2Q4F6ZweaLfMq/
gdnan8sNLeFdDVLNdg3eBfd7gNhJmDM5NzjqJc5Gx+Mmm8kTTZ3MSgVoenwA
YqDs+fC80CZ9WdU0RmP2PGUgLJKZJ+UGyp8Sq5y2+2MAUr+/ElEkBNFIYxN2
S9DMBag71k9l6178caoSMVZdFe0bsH7kZ2IKc9fAe3m2TFi2qJYOo586F7lH
yv4aykTVA73pSDUeUGUznoeao9k9iWNRnd1mnofHQHQ+QG8kmqXakPA/AT0G
IuXb7EKXxGz+sWnZ4wiiZSzAaD+Z3/DyZhWsifXo6nOASaKePjGo+OnxeOxx
5REMYvO9uV0q/2TPvCpF1U1phc1tPFHY4HOCizYQjuS0QPhj/YPw52s9OBfv
reNjZf2PuDIPGFT2TUlScBXhjajW81uCf906cm8RJo6ktZNA55Vd0I1pPara
crpO+Dmxkl1qWaMVEJ34/5EG9ntgJjTyq6263tgigk/nUxOsiSri92sVUI1b
Lm2sQ83MwHrFHxdWLqxrrSd9sTPdajW5mw8OHGhCPaDr9r06eYmyZIqw76Q+
EeWBESXvcwyz0bEvtMDNpa0+ZOelGU9M5qWGQ2jk1cf/ZtHupIoGvDM68yIS
vkQbf8NTL+/fNgG8m6Nap3x9Qep+XMUamb18HIAqqXuyY0yEGXo15qVLf7UJ
ovOkAo69CgPJcgrAUzp0lugQu2Rl0AQa3ofPwTYyYEQr99Bnr+++IVN3lvDZ
B216xZhScwxryrrfycBWSpRIkJ54MdvtGRIaX1c6k+ZaT5WJafHYr7Thp2KG
eXskXcF9A92j/cRoqpHymkNnzhSnVTHCNbKzZVvIlbYQH29FF32l5X500yVj
52+6k3GEQSRpU44XKvwcODp7FVHl4jmBH9y7YIFnpWJhss8MclbDR4eQ2h2I
3xnRihjbAppyAWDAlcW9NCniLwIdwg7k5wa4msmJoCWTUapBrlZpbkwTrOG4
e1bihgajBoESSpuwGVFrLMOg6rWIANtZEfjW64RBzOMd6jKGkTzovrMtEPP/
d6ohjjT/y2OFMGD8LDhBKdYCJs5GzpYv30AB+0l0xbxqmezNcBgQdIvLVevL
L26mqkMsyqxgNpFl1BXD0tnWYL47tj9l1rBKgkwZzcx1FJYfJtP37xJc8XJl
N3Ikleo4pxIaBq1GDRC4CkW/KIBfKpAR4sVggLqh6kAiSAMUWElIVqHXO0Kd
XYb12gjXuK61n1cE2RspnqNgztNgJoeSn1c6U9SCDBhRXingDFti+cmPZpzw
kG/gR0kMrUydPynNVmTA05EID5RLB/rC7PBExiA8FMf1eH0pZFR50G4ozzmL
OkT1mtMdKO1qDyZJ4ax/fi5SnrY2S9hZxSiTwnnzW0NkcbOKkIta070EOYFU
IIC0/3EWBwzJ7c1An86DIpvhF6039sUJQ7JDvKkt6ySL/txxZ3e39JjP1tqO
Kq/QPXLQYedFYWPb6t9+60tIUscA2E3hFrFv1oDYnt9wGIHF0Srn0mF86Dst
WdWt5nrK+j9f+sjIDjyh3nL71b07PrtdzJyTmd4EbIJf1sDrqGx+H8K/9VxO
XryhfNstvVHhHZEcEa5Ld7UrcLH7Q/zYO6eXK3ZH4iSryBst/AgXvxnBJpb0
PQ5Q3fvQ8dBtQYjCwHuNg+dCds295M7HKXCgyrjkHTFdGrXb5usYwF9anwpJ
tNWPKPPDTzuw8yqTPZwf+W11tnGRMrFesVFNlg9h1G9gNSvA9qHxwx3tkTBy
mkACQZibeN4auRuvsXULQD383q+IxE6m6Rzw7scqL0wOqFaNUTRtWmsPuW9E
98vaod96lu3IadgnmMmFktA4/pnRdCIPUMP8ErGK43zc257ep+AvlC8F/PY1
/vJtv1cBmn6nCr3SceS2qQDpWXkt3B0YrvvBEKXirK0fV8rIWsrK7hsxH9Bf
lG47YY01QDQn8CtXDP/8NYTG2c40+uoL6LmKqp1/wH5gyZZ1qO8hYA27q564
xZPj0eiydDj5xPogN5EoA/uEFRd/d/5Ny6JSfauZ12AF1aJebvbuanbS/dO7
PUkab4DdPmbW9MVM2Y6w58nmHUiFYWBmcVMvcH4ONm5ILHvHyEIaiXNVHGh7
2y/Iw4Sw+QIe54hQCPgHaRdO251ozAk4f2Q9hxZZNXwGvIwS6kfMkonaQTs+
s46g7vFKFvM6zOXWn8IOM4Huo0+qgE1nI0gsxpFXF4B+jYjTJBlBZNT5kdqe
98X9uK7d1Ccd5o9bErtapK9dhjnD3IkXSZyRoyFNJz0NhcvLZDPwZb2PNg5S
vd8wJNkfaOVI6Vi0ZCnBHmPVhn8K3NDiLzrlzoE0AJV/SrRmo3ZKwAWn2C1i
JpiXlOBR3sO9uoup51Q29Jt5ArP+yUC8TEn2T/mYBkhf+OMsXgSbugs5x9KU
JAIiiU4sGaXZr/zPFyC1fam8lPJyPQO1eVyETHp+0MYGVOuJoNbZH9Gh7XEr
yipCn1wtsO/c+XFDffrsLm9Hp4TbYT3WpTUjtf5NmuEkCDBhZUJ46NiTTyFU
Fegcjzuc2HKhvwmNzsYCovC3b6b4eKmK+biIm0yr2BFwL4qV+Kh/zEKv70cq
iyuokqpiQhg79MeIbcKng4d1GwjNB+kLueg1EAoqUOutGLHF6WvvVTKWgYTt
+L/ADdHvrgxUvXkEJuO7J9vzKLDpCSkhtazYwL9tcth+FNFVZl4fmmY3g4zO
jUFeaz/uWT64GRc/QteDTv4T7F0tRGpuLoZLFByrkUxJ3GaF3UCdwjixdSaE
rz6QBoLprFvp0KJfIuKAFTy70Ovx3eKJuM+ysSo6VuQO3ziLau6XzIlgGqdQ
tcG9s3kHMAInsQd4X2l0ZR4hBOgcGqXcnYWTaKz3yptlv3W0PhY7Bqvs7ZwL
Eq3zl/iI808MbN3yo+ZmtjerbwI6kwGlWPS6L2PtuSECqZyCjA5eHwEkiT8H
8wZlAJp7mVrzx320uzozEwsnGrmoJSotiGQjytSejR9SXzB6kWuLYmdVO4la
aX7twBQHSON6d5CjbhDhvGOg67qIUQqLAku++jLcoBYMmnhoCqrk70+DVxIi
YL4DdS0GQr9Ho39A8RgnwAYpcz7AyURYQJbsI1Kk6Q8MrvWq54dzZZRV720T
xH1SIqaAfdEbTRXKmP/LErsEI9QL18nCRgwgOrou9kL4Zq6hJ3WBEYbU60ft
lhOpiSkESPioo8gdd8F9wnhcg/QYnTG5lLiWC7vy0YKYQpqkDvPy3ZdIYSyo
LFNOOj3RWQwmmrwTOp+axBB3rXmITD1QklS3YZvQtW8JKSmY4MmlTjo6Nupl
HQfSUJp+1o4tMo1jwTAF1dXTiRThcD4Gl5PMRo6dEWDTnIXd52Am00oe2ibP
taWAr8f/eVgExO9k0gRAVnVmjSIsT08zPbssPAQNb1AyuQy2EVubpwWy6Z1W
+0HV2+4XIoRMP5nbmAVPbHUVwj6EHbBYVaU7y9PWOu8n9Noi8Wz8gz1mHhOF
0tpBbAH7H7NeUXAaXCCUNqEQrBIK47UTSpUxKw93gHmwyvFF9BAgoJoh53Rg
YQWLUQSEpDjKyx5vFcd2Iv9flME/KBPK7kiZPl13TT62dOFRZSuIAM2twvzB
1cA5mjhTfts/Wo03yMPjb0UA9wriQ50XiOtF3oP6K8HLH5baPi/hSNPFaoTl
tBgJbFNZTKbmrG3kTcOlv3NCPBLszJhK3pZqYSb3ZXKWIaS2rN+Zi7jkHlqh
tT1o9a5J+fzalOpwPl2JLsIPPV4w8yJq2E9FLZb7gxygKZACwHXyOpxRVPsS
HrR5H1wgytnc/kQ/MHBzlx1ox2pKqox4fjwKtCMjepStflc8oNQZ6U4rq/oD
OuD3k6WYQM1Ij+8ZbGYorm0QSu+Ow0dD05erWrvpHZMP1acNMQWJ4D3QtlpA
sk+nKrAUAbbDsV4qCMmlXNXMl/3ukfw/R1X3qj/0VLN++ZI8OvussWICj6QP
vGzfb4ZZzBFhc52SxIkAvmXX6ERUT4Hoi/8yG9aUSghhW1LwrEDpeif1ntMJ
dwkpgqyqf4GY7QvYyOMug1jayHFMm/qySTjDXasZaP4nFVPm+wefTNGrlwCp
FMtuuIplNZGOE4L3XQa8+fJNrFPe12yn4dMTLqPKN3+FDdSZS00E2OA/ZvRp
d5zf48ErCbT1a19R/JbrSIZJurycIw+CDm+sKuFTt3U2Z0dDKO52LAgzitJD
pIaLVC5wkPlE77dvf97pkZqHgnQ4MAUBLje6k25xf8IlZLLr84DxfgcAFZxG
p2ke3uA8Fwt+0nD/kWTaTad1/Z2aspWNVGcTVmGsloWfPmYJgE/7fzLnPHpm
TtsnWaeAILDYOSWWWOGy68EAbDD4PD+W6YMHVm62OQU+G3FLE/LQrSFrKxiW
hj7Zf1qxxBsURD54sNggUugpUIOt6WITPqnxZ5Hdzf2XiM6SBLxcofqitQes
TjiQs+jV2CiB1XN5vObC6m/Vuk018H3AvHsWFSH4CrSl2ug3D9+M/ZCRC2kT
mFP9F3jO9GiLtLmALhRJd36vWnGg0F7NcfEr8EZbqnOLnIKZfM/UJGHu0KHY
qBwqVaI0zb/jAnkKv+vO/v4lrOT/bc0OeihQMDxMDjv9+EfrcqqCplkEh4rm
BFwgMj3DeXULf89GLF+uFX7YHFFlKpA66vd8zTgWaRnq0WlLhCGUsg2BqMNk
wBN3VslWRXXnGoIn4KCabda2YfDIITHi5rUSBhhoIniYRKnkz8QgxZzvBoga
z1h97CzSIBQ88k/x/d35FsF8BrnwgxM6ZtHz9NSiBQxVV+/+e+VcARH88Pj0
C0euYyb2pgGw2iJybx0NuTmAD6BOcmYR0p2+EyuHn8kdhw8w8am+jRCYshl4
vBniC0Q2bxNf+d6VffaQzDiDXY/uizKX5DYa+qrxc65pZg/jKWrXZFZG07Zo
+1j6qWKx5f/FDIL1ikmGDJ23UQY+EIL+myD6ulwP9XlbZ//rsNLK+feFUJ/X
7o/kOeHsZbW2fOcMsFDXX7W5CWDVvsv6NL59dRfKOtdgnB5NPA7kiQJXO3/w
9vIADOImwo0Qo+/Wsv1LMSUERLidjW9pQlZYZ8lzjdvdjOIAvhIWCBUGKgh2
SHg5qPTmzJB6xR9Oya/Z11bulekRvvf9IzCrVKZrq1MLVDMkeQMaTYOVRg+2
yiRzk4sBCa3uRjwSorjT00Hi/bJ8X0+G6iEQtemcQ/BLkffoiM8x3EAK5A8a
99P8nus9Il7eKvq9xT4gzB5qAk/h/O/JArVfINCD9rxSmqJc5f6C+FtADnWB
QSZ7qXU2Rxdkqac3MIZZp0jxWZ3EiMrj5G5lnS+Nn5x8y5NLtyH3VdM1vsbr
DcFyi02h+5CoKYwgxRL1SnyS+f8Fwkuqw8r5cre0qygR5oZ/KEu/6TZnIUfJ
vH+Trt5IIvlJQ1ctmyB96vyNPjQs0vDn6vFTt5S9QKtq6v8w2F5WkmJL2Xjw
D5Ts4IeU7U2miExwtaWDc3vp4SKhzluZ+0zQX/p7T7TlcH9eNBd4jQikpaV3
CjKFMValMzrY1H8B1hgvvrLPcXd/0Q7eFoD02maQ82EfTmZyfFql5AvcWaje
uG5IZhym1zNAOijJyE6jlnAAWxc29VumB7deBlqt6x5zM0OIZZd5p+bTHnii
wPY8jtB8TuVXS98t2FA7Ym8f+6L1D0DPnNa6pp4UEZeWNgpDZ4oyP3Hj5YNb
8VsjCfDvLm9mF04/hJWgFTw7LbvTDFvUgejsU/6/KnqHW16lO4df6TOYX3J7
ePWCON1odHDplSXGwm9UkMduTspZr3x19Po4mwqGQ+4BVq/Tek6ZUslaRONr
Q25CLOlSlHh3JXJlMpWYukA/+ByG58pHG9Ge6GhGSe4ZXBSMGyGbZL6rcKL0
lk+ConpdI5VtXGv7v8p1kt6bcve9yn5HtghRGI/leq1+6v/R/BbJBKEvE2oN
78z9WVbG/ZtBYsxidsHdGXKUzbjw5VR8gekgzC258+j9Hz2hXbdpmKua4JoX
HK2pHG3ntQs9Jzi3KIC/erm8RRNdDWDp/pWB3ba851RR+SC1R9RenQUWjmbM
9Tq7apsnEdxD8W60N+GE8m9yHHLTlN5ToXSSuhl0VyNC+cPTaqhKpMzcUyd2
45I7LXmU1cMoKphEPzr6a7rh3/Z+TAFRM/JThdPvxyHEBMeet7d4NUw7gAGv
qG3xVZ69o+zkujUla5C1xr8U3JtrgdrBFQwQ6cxfDE4U4v2nyh8uOhJRBTSL
wLK3xJemiZ1YQwwO2Gfd99DJ8H/G/wL8nSwHXHtWGk/gEgw6Czihe/5ZulgC
+h2t9zAUQIoXPeHBsgmvxitsznpN3MkUk3RZ6iMDU4qaqRt46OrlM0OOWuxj
XtIlHmIZfnmd9AzL3ifL8mzuVr248r9bOKn7O0GnX5JBz/miqTiGkU23jQgw
gXgYSRmWYRqKrrQENYwOt3rhrIxgacIsv6ZdkkLcJys/VSREb6519UtzDRyH
QTN/bCPBwQjh1ZuoSZZzVMjbGZ5Z760hegcWIGXtFbptf3B7csKR9tJ3ipCz
MvpwJEWFJsMsWooSRfKFfxJARg/sSfolq8ay7vzoBft4/s9qlQIcllULyqKE
5DmLJydLDgaekRqowJI8Vh9TGlfx/M9hlsPO/XK0VAO59F5jwABOpXP7QzOo
SHrGaxT+xfutQYpTFthf+uELxQ+V9zBMmNG9UM35ikftct7EuXj+VPMfd7hh
JEICtuUCGLzsR6FVSAiXMJv6R//KUO8FIPgo8iGtAOm8f6JIusCInLpzD20F
Owh0y3HsxJxo0oBu1cju0LEVWv0GmQYoGxwPrRveGV2fvzBw0nmOyeJz1HH1
bTYMuQyNBlyzv0IgQ16vVy8exvgnRb/A44l/6jL2F94yRZVxuUIKysqWPI5W
G4tXFR6QuG3ggWhDxvQK8QCNoxBPegsovBfr6FAI42IN7JHKNm3PUuMl1QLW
n+A4X5YurZTbeXDtvVIDSP79CMlIG58Hq3bPZBaB2gdFDZMd19oKsKbh0pLx
nFHGxOwFNp5ee3eDxkP4Z9qjKWPvtTHvwcnLeKK+vc2NX26CHqI53Z2NHvcA
UeA38/wqH4vgmAwmpo4ETBelZncaqhZ4CllpU6kRTTwmSTCB95dLIDAlhj+O
JDASVtJUBLkruy2zRQaxgRn7udZruPk38lBYDTu1wwOK25yvUUNQhuG+HxDp
bjQYbif7n3XV9h2Af/Y1MvU2tJ+1iC4GvGGOh9L13zAcAxbpvMu48PF26NrS
DUUYKVn5s1oPSjWHGQjKqdBvqq8rddlbRASgclk9FvTJbQEnFAtMcSsFRP6m
rDoJzrJIgwNZfTTveWxT8U7OdOB82nAuXyXjqySb3199JfA83Vzn5SW6LJ/9
Emw1ne/nPty28NK/XPdmNbhbTRj+lwauSTE/1IwmRdR08StlwIEp3ME0VujE
Psvn9D8pWWhBiCLQBwQVizC4GY8p4QjCe7dMsQ6RAHmdVq52/FkOtdYOxWCP
QTWYAVRWYUOg05dH+bJuGunqX3G7EvOLwcpY2gZyH2CLNel69gslnXJDmE+H
ZIPvft+7TXoAoFAe+dyHLs+WVjbSdbdvhpJn9R8szSshdBD5g9hOHi4c1dyT
ERWpwfdDw/FJYWugfBR6D89yFuHkkDqatK6NgeOOM5xH7WVbQPp/NFJVK9Ux
OlEypV5eEqv0uiU/IiCX5lYbFlpp32UoD/82mF2eHLEshmum46ltae7pNBQT
p4B0vQk3oEtGr7HfYY8Y8lvT5YgvnrhMD2DLeV0N3o7b36YgCiTwZjNIcV+L
eXDN97tqEmpu0qe7xiYou7gWJnnUot9jY1lizuBg3NjlZl5moJOv7tD4Q0Nu
u8w0gaExwmEQ3cHh1es6DXiJIVWRT/4zK9d+sKppMemhNSJN+Kptn5WfDQbB
4sWJfml5fvnO0R4a5mrKiShLk/+vhsbZYBDpGt7h2NL20l1s84DoNurxXpgs
7hdJAIxk937tqbIzE8vLKZPCG9gxa8nkeZsxKpCC2W+6F28ENunEwD92GUz0
F5Y5jeIdQosrvaSfbA/JJdRdQHk8A/2D3BohHfgCriYJYew0o5FzNW88LowL
EpqpK2LkgPeoWF4bv00mphqsyR0Eo2EEzEP6Eqy62LGrOqT+lFmuXTUbLM0j
XP6ykNx3eqVbacFZKFE/s4y5ugH+PU0ooJ2eclX+Ig8iN70lxNFo9OJrcFlT
1KaSsRcdzdSBVLLme3qUvyCzyKyrwr441bJT2W6ZV40ZpznYiwlXV7+TEROl
mIt6k08COImgb0ahruSu464t60i+dldeJKfT/H9zu2U0gplWpEKuVaaWOZwy
OCWsxypAwCAOyss7rsOXnrtH5TJtMY0isbtYh37weY2gUtsdp7r2WdzujN9e
GFAtIWHQgg4WlZqecBAgr4G6+02mAeCxQVFzT1Cphpaji2T3IrQLuWkoaJBf
9fbv39zE29iUdQ00Fmzh4M0W8JUCDZcCOlKD/8RJcASyWsv/7Lu1mmDggGQB
/qCrKGDdlex/jV4ad7cgaHBU2IKbL2Y2crXvqBrwXUpGG9vfbd0zsw9h/v9V
F2m0OKv4X+x36xOPQMKd27OXXf2YJpjtnnK1gkFInWghR3A3b3J4sy6s+6fs
iyhdRI+E+zZw14Ba+fWWI9q7bBy8iouH407dZkVyAkHURfBNp4YzZBZcGySL
Ign579nQB2R9ngIlaA14yVs4n/T5BhUx5YIL/O/NDnq/WnEzAkKgmZx5Kj85
Bm68sgOupebQ8QL0me7PYjqVnLDI4WUNbsZ7uWPo40Gm20XFY/shGl+WbpiE
lGEIwGBgiZcFbzZqriVFsmqCChRyy/FjO0Ov68nL1Exy0c57dHeoBkQS68tT
ExsmJ/69fdLyju2jqcGoptppk5UfyCcaiZiVWYTEWtWBQDvl+cNUyZHl6zdJ
bHoTF5la9Jxh1cQYIyJtC1hJOORokcIfS+0vj0gjiSZG4LBaj2Jg2gXzsmy9
qAxX7Q0gO52YYxpMfNHLuVo/HSkiQ3zIjyITctNvB6ERNs65Y6gdH0F2Hg6y
vBfe7comaq54tEPdS2oN8gFr79Oi5R6yFZdBrAsYkllJiZg4ANwrd0BiMg6n
pFW/Y+At/y1A5T9+gHGJi8mGyTCCrwLldP0GYgU/bcIM98Z1kjEj27gzP06e
2G4FgMOnhhCmeG5Yf7haeB1fSfk+XUREIfg2hZkSUzuFr7hAMYz4jiA0UG6y
XhXh4l3/eZXGXjDtgJ7FZSAL9OtZzCK0600hVGKCB5w1phF1a6P3yfs7+pIt
zSUn/iaCeDhXHwCXpW6PVeaEodflaRdxzTK4IcL9lIGFqEYzUW8yrtvEvpqB
xEYoAfa9hG8bHpsI/AWe7cce4ZUyJFX//vMfQDtGYk3ToU4opEeXNHt/RP+L
CwallXzfv7rzC79vL7KT5x7IQKd+bVn56m5F0AbHGC8HO6dS6O6bXQFNuJQN
5jcHr0zJwU6qOvbmfE5NFldM0hUNrUXgNb7BHAZ540e8YS6gb17gFBScoZ/j
Zbeqy8lIVuOQIBBSIwjVzEkUL/fr0aCPrUtbl8Hl+Hr9PiNtjZ7r9CEN3dCo
vDRD1Is8jAEMP6RTqk4TP9bMHanI4RYS7whBZMY6yqqSSFIFN1/WS4Qg/uQu
a9rgtRDCmc+lidHAHU5zSC8brRYqBnskRnr+EG2e81f/Gw9cIliUEQVOezBQ
Kr2sR2bF27cPu8mhGmMCHFuvTKNX++X3igAqcYizq5I18Wyc8JyspgtnieR9
tW7tGX35OhRFNcWZ2F5J2d9SN5BQZKWJ/gtsxCt0l2UpJ4Til082NAdm3UPT
K0457Jo9wOCndPT6f0KbtWUa9mhl/DOVftTQVlW6CDqVmXIqK7QNeZ11lFdG
mj+54ioaYv0W9vbW9TgsHZSjASvAdtggDDI6Sd4lHocsnMP7Oet/KM99ZKeT
/JCsUYMeKUdNSGEuysBFMRtarG159OJHcagD5VZXHPE6P0pS8aZR+lDG/TQx
leWVk9DQrbSuwNM8rZ6aNDsl613RFvSurH64BefQ6JkNyqD8cN90cVnbUKUG
EpsVsq5JnfhgBDzb+/9f+nI5JhR0obMqoCC0Wm+tU9KKhk7S4rtkPd06V/Ny
c/ej3WlGcB1IP3cQcHxgAQPsARszeCHzUa3MoYwn5BkxH68XZNjneKM2NTI+
GpJn2fUBtk9svHj16Qe6syS1/LkSI8yDP8Zt4c+ZJ3oLy3iyck+3shysr5LO
TUiuAYzdO5Mm9gyz1R8dv5uZpuGKTz5vgLpHTlDDFeSGhQ8xFTXkP37B4DGt
jhCnEhWEdKjys3/dB62Q9lENyXjlBJ/Cx24xW13mp4kGevGfwAbEkgW+/qPj
uDCBcGs95Ez9XW5iMPp5sHfWQnLx/jvob3CUkjKBYkvHDC5h5rIxmKTOo9ZD
co8MdO+xLQVNeWcFksoTPnh4DZ+WeMfXn9NjGL/cCmlR5UD6P9jG3F31LFoo
z9q17+btD30Lvp7+9DzKrSaSOpjrMPuA77w2Ib4/LcmerMwnMygygTHUy18z
Do/HbvDs7qB0H3T7U2LfQANE9H6H4odaBrlA9DDnl1Og0tqi/CItpuJZMvVa
r8PAskiflAcKeZDzsGepHW30V1dd60y0dwaEe7VGeprwfEGoHIt0llZI0hwJ
ljTx8QnGH7l9/i5TIbw790HdTsQBmieQN0DUw6bXG8WxL2n0pvbVb6d3FGuz
Z2PNkAGiKI5k/cg2hayiEE3zNaPpNkkClWkLpQV5GVoRxkbBTmL05FmOP2D/
Usaeeo2I2j6oC5GujGt1v0W76vvHtIfkSZOs+s+53Sc81xhSH4rTmVSUA5xv
Ptn6FwXcoSMLQiBPWlyc2AVd83qWET6/GjlEJlc+1N6M4olUUcAiO1nvrqqI
0jWpBCR6Q36+PlsNtyfKjEieK5VT9mLxGa3zSC7iIvW/VIuuO3A8869InvNk
H1Y5UMtDRS5Hl1lEKLFSaiXzo624dN3ASC7Gmp341G6q4J78HhQ1Rb5oN260
EIwnMCfI9hyPsAOzE3kepbVCaQ+ZwsETR/MBGID0wDVVVyjR3P6n5H5VS+Lm
KrkCVYe3JklhktRyEisx5MkpL7JddbKMVmrzjxDIzNuFHkihSoCZAgZr37UY
douN9ExEPEH1JX9vKFLwVafk12S6O27AFCHp1U995oITzctPIEAmNAYEvR1M
ZgsBdqB/RnVkogEoqAoFcFoa82Ighk4KUaMGiEVlZ2CGd2UHZmiue2OssAFk
5gvwcEWsx/ECiqg69TWrk9XM1ygo4CrHdEqn7geolEkjQ2arn+LGruBrXbew
dS2LUWcYAB94gf65+HP3PIAxsr4iSgej8mTrV9x0KNLtSr+RDHgLXZCNSya2
J+DbpvieNe8oOq5S2vCSOeSIqjZAYzTxI/crDbV/eK+mqwDXK8UzjH/NenQN
xRw7CtbIwUryGzV7dQ0LwWhweP4vwxW/68zsHTpElZsY7/5un4j7i5Yb6Gu9
NGXlfLRWVADHByEU8rgbftHRLGWjLyB1OFtradL2TWVn4W9HWxBR/SJ0fltS
leRJtLLhPjeVOT3kxJJDQbnfcRhvAt6gZkmHjqLDV979cCOra674aiCnvGyO
CcMSIIbFgUtgz1PTgy7Wp6DHjYaaw1fxXoEQulkAq4hc2uM4wBQaPZ38BqYc
sOV+ePBD+2shmPV8t+ulxwhT1YmURNG4/tZ2GITkq5TvKyes66diNLjvGnMF
RUOvMnUI1rHjpZ+GwZ/2yYPbO4mjPmT99PCXCiXXZlgzUWnERy54oCz4/QKy
oM6Aw9xL7JGgEAip/AAA2mWCouDRN7w4M+LMoTVvo0rILQfkjPcHRpLt5Lh7
YWvJKe5Lcn7h5O56f4UPIzEeQzzBSgp+kFZaColwJSysf/l5bYX2xeGzlVzr
lXSIoyz2INQVBI+WlAqYvzqLEaIv+YCQMpdNBr4gNxNZhFXxR5cqdvxF6Cp/
uh0iDu8lAdfE+f8UnYizLHi6PuA0onlpsy6rK8pHKqbijfvHTxbWgr3g2akb
EA0K6uyO4TjLsX5xGVGx3r3FsNNtVg8mWuxH2d9tFueP+xY1MTVqV/xVPe/8
9z+7XZWo30ecoZgQ8SQ+iFDDF1L43yfgAoIHDipstUbKTZE0vhEsfaJvrSAh
XCN4I7Wc1sSYilb2ya6P2HfWxbZ1zU+jP+v/fFWV4MOH/8ELslfrq/QRXxxs
gOq4ok48H3CFzcaUAV0L4RveZQeW2YZ7ndB+JiPy7EZvArQoOnW8005JoDwk
+NqpSrxhMgUZsGVF1ss6rOOhgw3vBNRSL+1dK5AwRm7H538hXcP8VdpTc8cb
CvdA9tfHlvglxnmwC9gDZb328MNkswPbkw2L9c0dWhwGyARx/hHcJhoFODdB
E/7BEqC+UeBaD9ehupSOCr7JqQOZYpJyNmkKCYsyyv4htGQeXRb+UsuW0qSo
OJelSeWXiaw7FePQgBJFdtoxO6a5/P6yFxTExRz5SE/dybfUOtDpfDHWIeCp
080exbJLdYMOkC+OnjdYUlYnQ0WlSx5UbCJ+rKko0iZbZ8oMtbLW4dz97Pxz
rB2N5tsMQhZ9mlUc+t1kXK6TBBmsjRFbjCYjouXUsG3I4Zu5rlFjI9uZl91g
fcNllU8/eZjFJ9PskNtgY098Chy9G/5yBxV5Lvo+8IY2aVwqJrwfrfcgrOJq
HDAT5swritFviV+gmMGxnjPZB4mjVCG5fD0+UtG1jwjJ0vZoI5jFypJmxosf
yIkTncdRj4XUob8TQcDmZUqpR2ux9jV8dlyJc48q8Y4/wtLfmhECZe7YLw4a
kJyXM9lFF++ziGfYgKEzFCSZBiLzEXvSvEUBPCEYy0hh7uAS1EAipCCM+x2z
awT0t9tQ8cV0LXXbURu8rOaVclzdlDmz5o2nEWXMPAUDuPkIx6KzB2U4DTgF
swMLXJB2plzbLprIZK1V5tHpkntt5uHMRbu463zcyLvUbY7/xkJ3ngBdhpe/
HLdxpJttJ52vDUHVjnT11o4lhGm4kdKLeHZ6/Yv+YAElFV8/A6EFTKqHVlqR
JpMuoLtwX0UJGEAbvGGkZREt4+KsaZB5z8yY2kCXKOinRa9sQWGyh3qOIPMy
koGRnCe+1bSdFkciQssO8sKTy9rS49xgxREFHIUwDNwYWqEFX/JT2hp63cbu
6EAoORzo3ajKNqZZFf4uNzMQcVDymcU09m+e3V3Xgk54M59fQGt7MfHeL9bp
nmUq71mPlnowC7qhya477wv2+jLLqs0Viq+js5NSDBvsOUPqbK53SJ0h7OPj
lLTIXDnDAfDj+X0/yNR1aN50/gi5ilpjxXGsvZP3t7Euh5vB64PVOHgSRJcM
Gxh6JOAGnIu1YpCcpgehH2ILCdLgtc9nWB8oYDHIZWm+F6G2U1vHjwx+A4YN
oVzCm6orbwZ4yjU0/TT6BvnyJCGKlBGMvdz080EREDOToSVamGLF/Hom3yhL
6BFvruhM9nHpLsEJT5lUecvZKT2iD7sGN2TWioAGtnTB/XfCmpYpg4kTgOgM
yKUbZmxqpc1mAaFDQCd1IPIbZkS2A9LuxBjB/offViWhzpQpz7xRBIVt+b0J
DKBf0HLwq2rcqNdv8PvYSNB1rxuwSypNPhu9Xt46dNaA0EFLBOG/rXmnQmNK
kn0mo0hJJoOJpxUtsgBUZd5ijrdN0t4RNcySCOAo94EuM163/18T8XrFikLn
aBkBf3/3PhCjriHTOIbUrjKVsz4k7DBUmfbqJihJc7CTB5+RYFl/0TUlgOjW
nIQIF/gnwXFjHfGSazFRE0Qp5XualHcDFQpVFv/DlQ9+WF3eyQXRRdTf3/aA
gOnALQUKoxlxhYiQlqZbZblfsVoAJNPz5OlCbmKknaVn1rGL6iZq4mXPV3O+
c/V0cuqf10DKJ9EOobS0368UbfcuwPOsJuVSwjN+u8OtmG82rPjJDQL2dKXk
7x2g1vSImRuvUkUF45/NGJHDj55VjJqsphebz25zUo+bPXFvESaWY9/OhB7J
E2376OgI3rpkJ3t27BgciANeG4i1011xmejOn8zZd17lkze4y1hxOxoB9UXH
ZexqiTDnbaEt9IQDY1EdgkCa4rggdN19BU7X9OTrMo1v3Olq3XB8DT+C7hv4
JhMZmfhVTB4gPZg5j9U0BKEuO0vYg0nmoNgcIicvHUKIm+67rfEldF57B4dz
i9gtTGPgidmXvneuOuDc1DvtJh/adki8ghrVc96ztlln7ApY3Z/erGrLtY/K
yxFDnd1BLjELMeZELEtkacAwnipYKJ57/E4iSkPUhj9qOU3E9MzxyZX3PCIs
iMjgNChvgI3MmHfg2QucB+Xjk/zMThMNGKU6bZlk/7QM2lMObrZlMGuYaLm9
1IgdtthOIam4iTGIREXuA++EGq8QUTKnXs7IA6ynDElCwUI+8ySDLqwe+4nG
oxIyLARzmOTO9YH/9mpX7pnHPl68LPR/3LIFhvZpu3FlRSfTjQX6b192xpDc
0w1O6vAiOyGjVqIyLINNeA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfRKeqS2XcDBkkNXkBZ3YPciXt0K5oiPvvleD9LQwaA46/ky4fRP8IIPeRisIlYl+RoMH/KoPSOIwSGY+2RlAppr84Ty37+DsWf/s+jFs2rFkUmPeKVVwI0MOD4HHvmh2VVWBrGO80+S2aR9upqQv2/hpdhG+Jw0/MqDxqi6v2Ioj7DQr9lb5KW66nkISuP+hl8SJ1/nTDy6Ed5tEG8zm9qLoi4UgyfG77vazPPHUDeNjBgLC1d8DzIsWFecYEZ2ZxZwrmJJENtoNDFp7KEb57K31YNCLRAiY8ELXUw7tIHQxsqQXlv1n/PPKM3nVwa4fBFC1JfteXg5/PR97Kh9K0gIRMkWtTlw7goJWwfnBs2qQLgxXvtwbgk3p7oBYGpxJN7o8u5BBWIQRLTMQvQ/+hNsN+7FY/eDtqIVeChtN0EwHIrUo7ksOxlysTxQ80H99JkQcBSD3dxQjLSQCV6mBFUuSaXpBy9O2xYPgaUQzYFC/DvNRUSHGeTvAKUx85yemyH3SSxrSTFVeTYngWUxR+pniLa4i+ZtZn82SIbQPrQW/2qzOgbr+RzbBbsOXEevRwVtVk7RpJEYMcLNCn0Nr4OMfmhSGnh8+skTm05naaget3mSmaMijCG2/iMKBfkv43CsHAQjbPOivI/1vfxU6SHPj91YnxiLSCou28SevT8aYSVHeyhkZeAd2EQaraNwF2TR2cQ3YkVE9tE9UgNt9wFi4wtN/d2K6xwnBdZXy+Apb5SeN0hezr2hGht8WdHsRCEI+kf/HBPZEjy+t334DLAP"
`endif