//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
B6LgbOUuxgU3fvcfUGdmz3sGTPsNVPWdBWN3fRK9oeU6/yN1t1tG+eVCpJlJ
933nQFXfWVav4CMke9zCY3AJjgNxnkPwlGUfQdjA7GAgUjaNi+RxL+jI7GWU
tVl/oytL3izhBu+eldzbPEqFxs2OjINNzfwxX39KUASyn0LDdlVTL5AltccF
NY32Gs0S5CJ4b1Mw4B57vadM0SaMCsC3P6qNSOyPFjVZxvm9Lxt0lWuvnbib
ouxIKHJGGe5pR+2GbuUDYD6sOqFYx6NBwTkiwRech9dxnOW/UdyXFM03CNas
I2RhqleBmmfmOE1kxLG7Jjr8oylmSpX9NyNUa9WudA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hAzUFZ6M6GPVK7EonNk5uXXpnIqw+S7+Ws0Q59tYDeImTxc38mtxtmC/QhzO
BrKvwXbC6fHgzB0U2nrz/4rSV+WYlWAG25hGelccbclNYNFEgbxLslca0JnM
0bkebYKyXKKMu11fYU0TF5dMKsD19nrypV3hsg+ZVL1oQ/vxttJ7QSi86RHB
IDkLjFx4LkKy79cNjTCWgOBBc9JzAS9PjFEnyySTEnik52n9nJVpD/9eCJ2Z
yqSrBZNRN9lfAwrkb5EtWj5x2jaOe3WXIHDoMyMI6mVkrDJwG8IMTOnNju0B
QFROqpzy3htal5NPr6/quLEIbwkkFuqUCwpGtsgEdQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
BSCk2B7fTh5LAlRQCyBnWqqlXmRRa1mProob/1Rgb9VTdF1QgIB3sNKnGXfJ
2t4HREunnl9MO3/ldhlSTaMv1m/vKdYk2odUfW2hCnUosFxMKxaLBQlJT5hQ
SrXqmBIiuGZ8VmpS5ekH0aKPd4FzBZOEUeZP+MSRzCBcF7J1rQNjjVd4NbB7
DONj0dJzDeZRKlS2ddiUG+4E2mT+Oi+zlzV8uRWWe1PvsZ340VKRXNGD5Oe/
x3YqEc9FVa53pBunnU+Smxt3/WiBB1GPAzN47PfdwAvETGd/lUzhCvZ8By74
avBupr6W1RKjrBkNx5GRvD/8pHJvp+zPqMCvRGPFuQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FTXOwcKqLOU4NzX6YdXvFGVH8pgOFetKLXCGTnGuq1fpeZXqf6T1jRFGQEo2
somkqrFj0a6XMVQkISKKOdt1H/sfvphmgdkYPwuQm6QM9eAhdsQETmpfrq+m
JlIyTbNk26s9qioTOzWLmvP+J7hE6gJvzq4KkUevSaqzP97MR7g=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
rPcDWemkCuP+Klzp4Epbm/85et8Hfr8fC1ejsSUR0wwx3YhdahnOMKoGI5SR
WT+4HY0kVlNyxw4n3gpOsWvYH6c/y08r1gTJ+9YEYu8xeaGwkZUk9IUsGVxl
XE8vaK59LHi6JeIuc1cAhRxiwS9tyyYbvuRjZFOh3thXspls6Jx4C0UXl5sR
ol+Y8YWmvB956kLZ0KPzdKBpg08H0NzWc5Wwpo8Ri5GroD0lRF0gP8UVCgPQ
3jmsHMJr+RAfLNgtlrNzleqsJo8Kh06JQ+CvnzNPH6zALi5M7papqFpPpr8n
NlmaGQfX8eoW2dgSU3T/glKl/rGgQkfDa5kmIHmSZzR/VwyYgJUumfQavXi6
hr9aTJXRbFswwo15xKkZtujyFJPLRjSexK8lqt7+mpx5D3vZ/wpq0UGOcLoq
BmDx6TN07KS7tol9/rOQgTvJuSajyS2xO5pd0mDN433fiOWngJQVVmL9nze4
S2NuZSVTrrowvg96Z8HMiKhdW6wCPZaL


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ccDb2FHEiOFghINuQfeTq76e2rMOupK4HNGEs61AdTYYfv1y2TcHoyYom7dh
366QYBAbsaBJCjAfMmbh9/3Tlw983XG6yvOM4lvITBZOYGsNjdS8Jc3eqrIZ
tLsiUKwXOalCLcX1tVQPu7FUQgG4pAL1mkmqk0FqkZAh8hpG6ME=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XCU1tXMiLvTU/Jo80SMYcZH2g2SW8UOz6hmzru1xJRuzykyJ1akcSAi1d5Hk
ENBRtvSjSbb27lysOm+ZsLnPFcf6XYYAd/FwIGMB8Ps9aLPTTHn6pMpejvYF
6o5jtrDSQT+3IpAj8Ivkju5xJl5Z7ueC+GvZtF0wUAR2dvyaTaw=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 13056)
`pragma protect data_block
EkKKfeUXrHtwF1Yk+9bp7Cml+Wyed/tRKB0IrtWNv8zeu7E0XgtNLdaTaP+j
xs7XxpXiEPfhL4RXIq+aU64aG+kuByrhrb0228PphfBwfYsnLJrmnrJxzmSE
azdXxalBxafdq3+CtZgnwRjocTKMGwkD0QakQmcHFhtYRhRh5jHSrQz7LxdF
a0Itk+QAbKMXM2QYXMV6E6YZaZwn7ggFoAooxFNMo/jIh0g4I90FOXBE/Eed
c+zY+d2tqut/s85qDYxIjrtqiGvzLuR7qNemKyupu+DGtIa0aI0DLXbQmE5g
Lciuxx2sDEF+WZDIJQ9nuS9g8LFJEZjEFyMJWOsYFyciGIk4W4LK8mi+Q9cR
x7AocVFfWX9xIk/hzN7IcH+j95HIEGx1Deg8jDfj56tBRSE3P4tT4yl5PljR
jOgQMB2LT4068iOATKM7Sw1W43bO46MmmEbtvNZ1pS+BQ5fJ9HMObEyAmcaB
jydSa1uKuNh5pQnTaMnQw/4huc7roPf4SkQZUh0P3Z4TobZmex+b6OTk2xM+
KPun6a/GmE46RwhDz3fTJPthYt8BQjSuMkboaikTDc7e8iVlrh1CgeIss41L
5xAq1hmDPSurLmro4MlCVJZ6xw8f4XRdjJXojT+GHGiBui4/diZEp8SkY1pR
OSjXKrkZyrT/Wv8c1Qco5pZyA777WToZPAdHWGUHmw3bLlzhrwe214hQtRkz
Zm4Bvqv5TB7BmdL/IMnW8wANA4zSRNDko3TrljUJn0qgpgpcVDk0mg3xFZlx
mcOb9pUG6+UAlSxYhfB/Zm2nmvslcsFheGqIguFSE9R1cjYBU4kn7iRY/YWS
yph7+SXrJNuDaJOAXBJpDbzm+kLbLArg0h7aDxH90+E2xyKhj+wYGpxbSXWk
EeEveEQU6j64TuNTqu1C8qYZNyByRLan5ymPK19NqQj3Yb2p49aprFY8pSKw
JZa8rwoAl69Au/FnvaDXoCdoMFnOj5pPhAf1dPJtAH1JDrwF+vc2/FRelaKh
JMls7L5Q+7bx48EJTGNeHNaOuuRx6eEZA2UztWvKQfME81MV7Lg8ekMcWrv+
ch3u/DDj14MWlsqkgAkJGDGQQ3qQpLQawI+BzRjk/lrE88dKwMfubcFmCzWW
K7/G8P18zaq/tXYGVwCk9Ux0BBWXHab0TqQAQMsAMvuhbo4NSy+ZGwX+Ehoy
c0uPLEbOMQlTaeikEN6vKMiQc1D55SN1mh5O7lMZ3OX8Uu3qwf8zNS9h5FFt
L28QtRtEx5cF+861Zg32Oi0N3Yf4NRm6LmXoF/g//OtjGofY6DtoeI6qSKZo
xrOd63+GjMXTRkD76HMaVkXZKk3TfY5HrMsnyBXafWbxtEXxvjQwrLhFWons
z34CxRE4QCp/asdRqPNYXTqgJe6Os0WNRFnEUS5PiJEiUzhT6q3Z81RWkkEC
JQynyUvLfXPkjYFCYGXVm32GQV9pAcoEbTRvlmrtQF+bIxKOeQIDhF14CmPZ
d8PAvXRBcrygPC4Lp+ouTYa9zrh86+bWwbZTUHw8E2rsJek/OUEHLqoaUM9m
AUEmE+/Yb+XgIm5VjuvgThW7iGEq16ewOKohljdr4PbhJ9ywWfMcUKQRaIqe
Aw+ZgcOrUp4yK/oQ54ZcQ/ht5rcAziJcH4WPMHGP13qwr+EOuwBGHS1T/jNf
/mZOD04V9LLQdBrjqH7vNU28HUdVSfyENeNq4pA0RLhB0rt+LqWG027p+tFK
7EBLLS8MiB/V87yj9+pomi5yhdRZPJfbBv2U4j8AjNt1Kk6FlrDDpq3qSsA+
/8UGEcDIXuGNESgl/j6+Vu+gQItSAJBjlEHMs8kugHkz6oO8OMrkKB5Ar5Bc
R9bgduwMc7YePGjBJl+pCm5RUfgssqu5eCBdqqvypdZVyD+wx/6Uigv4bzTA
5KxpbBG8iIJsLIzk28AnFWXFYU4ChVPuqX+OghoZfhQIb7fuclYbdJTF2I3z
h4HKEymP/q/zbH+ISbE92MzNWknwZi7lxmvkMeNlECFnXdW6MlwIHKOvBV/M
dLMskFiD83Q2oCwYycGm7Pr1AfrGq7UYzd91xDwIZmBN6BPmNgOQY+A3cQjR
6OUZYrJkqbOYP0fDPvKC9NaOm8CLcDPLOKNxfYgfJdCYArxxwILxeJZqCuW+
ffDKU2D9IJ+Es2LbmAJKBBhVjiaLrOEYERsnqKoDXo+T3gYJxGTjIxTRcEUj
HeHrG+4RJQJ9zUNNW5Ig+thljxBv1xJtTbPwY6BXF+k+gkMBgUTg5TbFjtuI
C9zi1aCNIjadXtBE84tdq8WogFs0vIvC/6ERhjS07QheboZgrnsPSxLzirEN
DqUtVmZEBZL/VpXGxxh7Ry+P/IRHSQSph09ydhD+3hV1Tg+uAAwZdRsvmq8K
R/sYk8HIb8tfUk7wpLoU6lGOk7F+qFMRPhUw9ynTnMjP4xTyp4uGWdaxiPd9
Ig2BRU/1KumADwbP3dWdc9FOedcbGbp+X/KlvBPcuv2Nx+puAuef5FfgAc4Z
ROIO+8AriRvjB1HYVuQ/JWbTXiry+MAS3huRiJyg/OMOBdsPM40yGtpKvarf
2dKlg77MO/CVaDr/TyHDNFwaZfstpd8/abLbNdM4uiIKAeksEhq4+IbOeYGX
pxyOvPeqttctNM9ex2fIuK9pI3qxG/P56uRRtZmcZg0dRQaKrxUQTJDurc38
rezUv/x6alNDHbuRvkXybSc4r9kyNPOQRbUsL+zr/Dqpu0cu2NIvUBWoZt3d
1opgzwA50Nl3FP40b0AHEqHC8mk9Zg3INS/f3+BstmLff336559mIo+OGAdK
qkeSl9AGRIOn3kcRBh5D7OPe+le7jhsRrzjHRAq2hJrlMk2Yf29AkSpivkEm
a5tCOv5Mf4xrPHTWwZuXp3mbYF01BKCOGy4wACfLPDZFxtMrNLvzHvfnYAmv
fAgx/p/zBN8PWX0G0jtPl66rpzzcNkiCeB8aq9AS4QafIv8c+84S6RFcv5n5
LlNS+cylz81Pv3SvqGNtfOdptjGwts4m0Z/+J7BPPtfOIzfJQDATlU8Y88pU
m8D8HgZ/KI4V9SVaLTcGqzVytUXq4BPvY3Porj8mKcpeSPTE79HSHOUrCUc7
pFx4iFeXxeuKZLu30JWq9uM/QULdNRMvXz51bwyW6QAHXt9SF8grgrD4QHYg
qVdwrHVRfBdlJfAyfXNjUa0Jtb7yZjsC040Mgcvb2PBV2Bzg62kVGr1kZRmO
9X6ISpPCnfd24f/BlZMX672UjX1yp73V7fWq78TIQ5UEa2YyJLEC3E07mGmL
rkqwI+0GK7TeH9bKrueuTvcAvsUgLqcs1t6WkW4EW31n3PBeiQ0t6s3dgplJ
dGL8LnNWFzlrGnK7jqQoywgdHOHg4KrmgOMqPS6TiaQi44d9N5RJApB935jw
CNZ3xErd9sxRFGCmXVSbID/WG7Q0U7tTeYaWwxImJkJuCLYHmj5SgADYwz6F
MlQsVC+0RzwM8hNmzacCAwvaFerS4BTHDVVAura45zcLDif7Oj2cANy/4y6R
qgxIyQSUsAPLiFIyA4cEsX14NCAXlWdXHrD6144ZTsEWzxmObfuPsPZ2fl8m
rbfGPraKW+Rcgu8RzWo7+FxArBeD3+6aI6ehjbF39dGsczY2pjokywmtVD/W
j5304oS2W/ppCXCF//skfONM2bBAmh8zc3/S6JOJR2JhNf4OtzsRPufnCcGu
UJ2GWoCKAwjpzSBEP1HOWP7TPkW+PgsYctro32UE0O4fn9M5DzxLGIwZVkPp
kSSsiyK1K+2PtsivdmjtOhecHAW2SXv3FYIxDM3snc+4vVGAWl4yyzgSLc8c
2xD1x590uT4AFuxXBSjpywwjh+ToG1UUaS0Vbnf1b3fJpupwm8Q2BMs0pnwK
yq8ZrJRJKTirZjpu5snbxshrvDFIaa9kt/rnAsgpaB7C1VOaMBv/tFTLOlvg
EETH5nUYlalzrQn0mXnBEOBheGsAX70OUB0r9EpBscwBdj7g7vIunZEqvQ2Z
E6JcGiD78kyrbrDgLGC0OPvxLWiQxDxGF+AF3E7Qq2/0MAzf6IPT2io26OkY
oht5J5Ajov20TsebUQa5XDtn+kmWzEfbKOWWwfzLwDmF7rS6aka3sC8mfZaf
oPLyJkIpexStjm7g6M6jwFRP3qBhhztTabgxQGR8XfqOL9cUgPKyjk0W74wv
nMxgAe6AxuM7uwYvf1w2LrfoSMgio/YCbGG4e3ZZ0dZwwmsYtvIrW5HA+L0H
+NmUsu+m6BDFIAUZFpt0r/4rmvxPDUjITrAlNVlc3wkzw1joccLfNt/yvo0j
KuNP8yIzwnibUDEXI+iiTKhLMarQPLhUDqvnztFsCTGfVvv2kF+8nwu7EH4H
W4U5asVjjO5hE890+Ax/YlO7jJR2RZefjcGFhyTp0IwjmYF2FdJpZ6xCv8Hk
pPB4a3ePErH+pMUkjFDvhuU5pwz0NKzf6C3BruQYbImCGpaYUWa/ZH9sJT3I
L0g/jA1oEbziKZYkLdqssyC9XQ7pAGMkxoyDS7H+fkMVOA2CfmVD2xMsFHWp
8cuhESKk2zaQneJUFNIdJQVJFSu216gR1UUs59urZdFgKiUeTUuDf7PL9flw
T1LvuM4gD7XwOFPSGfFuie0YLhvhwLDYkdtDPXuBqeN2XJdoBYKwGkhbtZG1
ihhlsPDeccpiOqFnKM83M45SumX+TH2Dm5nxm/WZRIvKA2RE1V53SLtvEWfo
eIXiaQBA31cyg6/S4JJi4IMU+zGw75ZbB88Drtdb6JBMTa2/D+91Dl3Yx4pF
Yx5lSjQan9siumN5LUCk1tuMH5WPoTl0KVHSi4zLUQmziNEItQre3//xeNbR
x0xbPJFkDq7ToW8riHweJa0jqede/c4Tg5SWZ7rNI0yBaIVpzPAuvc51luPx
cD59nPzeO69uqGxtakX4ggWKT6GrR/ZpJA+LwEhimtRTyuvg6+exlKH/kIO9
Bnhz5nGjwi86K3H6zyaXBYF2e6fp14QQuJzxhY4vSNOIwhvx2akZ3Ik6w+b5
sBWDbdJZU1LC8Y4O6jcfJNis6ALyC6eWFfApdtUJVGETJUggmHQd+ZjUN5zl
nnp2ueTw5tPndpkpud1ycTtsRJ4+L3rF1ECHfFtXZ0wprJ6iteSFjNjItOyH
+8+UeNZP9qW4+tyFvZqKxmN5Y9JVv/LTq5ToEUjRLXGqOwPIjtglolrw4yOB
HviC5xOOsiZbUwQKMUxLK7+DZ+gaoYGV3DQxczE/WX4lOD2mm1a7QmcLFfbR
0cndIcr0bQVXI1XPla2VFZnX7ByINkT6kLcKL2G9e0onkX+YBb/3242BKY5/
7xTGzyKF5rLXP2qZH0vt7/762zlCyoANNpyw3lHWBIEc5/Tb9/ICaEeY7mfN
AdsiwU7hDvsGXAAD+Yw4KshzJNQAi88xrdZUksR2XvRul1gpsUCkI3KGBVkE
K9H5tlV2jcOwg3NsWsOonerYkSR1N6g/WdYSbRJDXdEu5kAL5VydnYdYOEwD
2aOnPMUyaeSXx7gI2zQFadMU8dQ2m5G+4lAa2zRmm0iNI2iWUQ/jAWGgKwUF
F41+2ihfTkEFTlYReszYkd98Uh38HjwvYgAHRlOWN000+jhaTSXd5HXSAeke
PO9VJTXQzKUYeDPNBqTgQ6/aN8QGrxlokIpN8w/wFDgQWgusxJeEfLFpOZro
f8LOsDEoApNFAcXvIiziMm1NUErM0GHOnakB29CFR0apVXfC7ACN4KWl1kXX
Q5UTQk3PhZc4KVm92sFfN4aeOWMUp/AIKUga56z6BAO0EuDjMcia9krk0nYP
oYNm47Z1XbS5I97GdEHEQ45jvooOTg/GlRE357pxD/tPw5oQMCF7Cwd3PBsi
sswJp0btGquj1cTGP/TaUIRdAMl5jTajoPysal8jEcsXdjKZMLIuEC6ksfSU
zpMA0f0151lV9CqroDKgREijSA8Myqjcb6sHiJbf6bof2UEK4Uiob9uzz8Bd
wHM1JhWQtpMJqWBUCARPcZ6Wkc5Z3UgbsKqAcZ5fHDvAI0kK+vHkrlH+d0uH
AxMC6VxxpLah/eGJsQtIDepRm4RTc2wsaeGzRRjYQuI8VCuZAjdqbsXttiOV
4sR//ULAP2BQ/379KIY1XlAOKAVzCF8iihzQZEJWOCkcFO/Me+Y8JSCxRPaR
FtPmP+jVNLxu6JYQATZc+ofg859KmTHpOFkAwmiqkwaa2mguEni6Zd6o7fw6
v220YLwObtjvEZ+eXhNz0N6y8ITJAB0fRWt7ruVUijyLySZS0L66MR20tsyx
8vot3CcsZtUfWyDFBWVhsizhEvAEbeHmxcTXSIzeTGKYzrWkSY98Mynj3mPa
AbDr6B1xWLFruIg5aZgcVpgsDOmx5u/QGFT2wVOr1CfNxy6HLb92JvodnXOL
ddee+LMU/K9UPtdM7tEksyjBGiwDG0xeRuLMpn63bUuBfwDEuJBk1WlTfT3Z
pkZ58bzZl6+l0O3DXNHSughsvZRSfTxCYWFkW6P4KIoAIb0H24EvmPd9ouew
cqw8pURcUUEfytmOEn/AlyY3Iq1HdagBVmLxW20lNO5mD4yHjHfT1rugex56
euvlAlW1Tqrg/lb0EMB0cfsN9ePwK51kZbV9Xb8DT6U/6g/YWGSHpga7t3Sf
lBvFL2K9QZTw5iNOl4HsYvS2/i/5r3V/9ebUi+x3RGIEsY5ABKwiUfmEz0dc
MtyzB83g0K1E4I8CimHeBkbyUcTZyNM036YlcPWIzT2yyHwq89xjlXW28AT3
QVuftZ0EXWIhE0UiR/XEBB/R1jsi/qn9pkbe1jlj1O9j7DnrUP1TrJA18BTu
gQOv1Ilz9ik6ayu+0XwWrd07J7QAwxDGfhhVxx0743OHjKfdE2DHz7n4fM+D
Lt+mxovwXvV0EA44GdONYDEuqKOyfK/OakUe4yFya6TvdgDH+7Cok99XetmB
UjqCxlvQaSVJ2cvseAL/1HPKUe8GFe3SSL71qtSfnwaGnNb6EWuxY3RJXMPx
tMHqqxd+QE0rsRsTzO0Iwa2oceiKqaiRS17xUKTsby1vvKmVoZtWpt1wCsri
pKj053p4UVLcKmaJ5nTCfQd4NF3oJJRHF2nUrn9f0pkeN11UMjNLx92qCNa1
Uf8p49RsDkKjJ13GqqGY+maYyx2uZ6SBe/0Pof+XL1xnoAwMvwY9uX8GmzVf
Prw21keS0RXZ/VYennGrArh1JhySte/i1t+LA/jfkq6tvxFMXMHP3fw1pwwg
2ywuOUKGOTxaEOEKlhlM8lgavC1xrH2lh+02AI0refWmy2N28hkH4tSdFEvp
M1+/rBCUhycjpBIAd+UfYLb+zgoCTTYqHFWPZ/hPT9T4XzY4bHpp5vumGBER
4pyIsZt8sWqZcnNXM/2bRLgdiIiXuL3Q27GlAWEhhQa1CEoq7NSitBDydMu0
11frc3xEtPIA6fKlu3pge6xT4Hb2l7qRvpYXlQZjR0ir417h16rZroZeOJ8n
bK9IFObLHCPm3fzI2fOwSfX5JmvtUyHJNMwkqfUWoHVPrZtzxYPfCeR2rkhi
56bazm9nWJ4UTVD7rl6paDepUsepf7L7NBb+Fr2eTummwp/UAaDa+eU91zNk
r5/n+tOKtrruj0emDfLFOYAIDSNk1w9N83LOICri8rnb9tl7y86f7WF/Q6Pv
zAi52b2K+Jrl6UnGDPT+KcI6cM1VsBuEIAs7iCrAlmqspwK8zcXEnhC1IpvL
xDta/CD3Z7wV6xH61q4ci3OLlRYxj0bg6ep7WZmwtKx1MTU0yRNa5LWDBIjz
3tNQuvFlTUWCg+XO3iIGekh0lTSmRD0aO5znxf9AtPJj2kzjojIZiIyUkZ3o
gjQ2DhHR74GWUnZOEqU4vA6T+I4ictI5haYYcnrGiYX6JctWVVO6UdQvtNFF
AonWfJDUgb/JGw4X0ZuB+GsWND+VoNp9/zqmiKFaQYOOm51xp2MFAei2hn4I
45IYQMRV7dE/4pwPZskTnJtgqJMqa0SNfXSBtgvjASeTEudAN1KnYDgHEIAe
IOm1T4rMfq64NLZZWV0djZtYScLBJHG8ATZ4cnaI8VDaCKeNGeKxmV6FLDdA
Rx38OUUmyvs+YDedCPpVU7fpVAMKznaxLSixwZbhH83wrFIThfgxSa4kQuQC
E227HvH7y4UVUPUeUtrjx4To3sFItQyNj72j59MQrVgHfzPUaA3ORLvgUbBN
8Lwa1ZmHqzJ6MuygJyx1x+m6xPwX+0aOwsNWkBDMYxykAAmx4EFEULjypaWE
P1VOXCH6cBwIyf+B66iVWKyIvebM7uEsewyA4vSxzedTflneAmSPibv/AIks
XdA+qK7nWdFu/etmLLogL3jOS2Cw3WvsJbmMFRf+MehwzdBJlud2OOz3c1jS
VmVB7voXL55mwVKy7HzD7Rh45JsP2LpW90hHydgP9tE95lb9Zrg694D5DDAC
OytFxzFfB3z3CqqqTbjY3+2MfZKTGokfItyLmVCbYCUfIkJwMKGrpnkTheuw
JsrCBwL48JH+Jh4G2xLhbTYabp5gh7wCfKwAFXLGQ7XqoBCnaOhsOJOKUcrJ
CR8/n0weqsqu9Pml8XxbD7R6hj9McMKp1vDZS8wEKFZEiWVp82fgH1oaIju+
+0totjMoC+KJNB49XPV8/OuG6ZbD7kgOQJLVfctcQUdPg65sIQJVI+6gw14+
sZAAnVDAY8ssfUKB869EF5cA6OyCxdXxY6uqGcxM6vE8lzmZQo/QtxEJeo6/
NJ6D8om2hRTuryEqoo7spFGg5mgBIIFSonQQltjOmb5jOTLgdMt1sCLn/1Z5
Fa29QmXpz7OQvfyBwxkKSzPyRNaBfJaxQ1NAH0lFOadK9WwQd9h0zJsiESzD
7g1axXU6OQImSTAM1qPngYtvbXomZgJlEY7juanq8/aU7F429y6E55jzio7Q
DA9HoVp/NOMldR/PwjGbXI5glVfYR9jBfsgLx6K9OcDsAZ4m1lTefHqwoMsx
v1BeYG2iL8Up1yem4L3lujczaAgsDKvj+edRXz9AtXvwBSXmD/2t6lMD/RUn
sCKMtkyeWujLF7/DoXG2b9uG5lyQmrC2kdzE7X034LkAcsSYnOZip0sFbsTx
qT2pilm3mIPSgK6mikwavMbmn6YSjMOthYCTg+8KAsq+6N1B0oDFRYQRezh6
kzX7tZTdL6uap+j5/p/j0gWyOHhkgc777K2rQnxx0N3pF6EHm7+48KHT4zpx
a5SV1CSQhjpM9AMoIfaIVQoTV5vE91wyqvkcTy5n9y9Tfu/1n695mOArihP/
2VskIT0dnXaYzASn5NJGiJmVSysq6cCfRB2nmd2zmOvIrjy0JTPN12RKFK5l
dcmoj2uP4tLNjVxgqqBpU5CxXPoQG2CY4IUaTLuyEXd7F8hY57ZNu6vUjYaj
Zr+vnXa8PyasyqenbWl8PAfw6Pc//aZRFjO83piI8oIC3OdPz7OM+bfAyrIF
NrJdSGQF19HOsfrX6PbXC0RXrFMyw3djZFwy5+nBhon13figtoXQCuuoMmO2
7dC0JpWxZVZLFpaXnICEjwTJ7YymtU7q8WNY/f4L3pClkBH+/yjADcLncFzv
aVSxWzhGpbdytO2nAkXpkiI1ecYqwomGAhn82lEuYGAr0NwoR5Le3Y/EcYVA
KwWMXIL4Riqh8MirQH9r9R9hus9IwKl+mNVEa9pkNQ8vsjNcfAeuLZZIdYFA
5JO4QDuoti/KVkL3tmQe6shE6M3dw/zG5tD8TXHei+aA4bQY1KMeKgcp0Je9
6XSoCtPykUrKws9TIuDAodWwnCKq1l6B+u70oB/u6iHA9Ls6ucKyDPTxrcoj
TK//O5FPFFmEtXWCNxkbvqahyrnN10DKLv2G37H0G9Q389bbG/gG3HKbdnpz
0JVS5Gs+ObRi51dGGasHUYzqfiza3qcWRzSHfNdJtEVCR/4v6wtDyCGDL+5V
t1UylW/+sxzpDbJX7mHdcS05lviqYz6hG3m+gpFAuLbhVJ+j0GVmh68U8qkI
qS1++g1sFL5LWu/V50+rXALfYLZMCjzO4PcF1J3sYE65P1pX6vT+aZtMM7eW
DEl5/uF+ZSdWDiSrCJhN8++fLaVBDfnCiOjOqUggkXLOxV4bDlTQJT/6TikZ
9+5mlVDeJ0FTEsrP1fS3b8Y3nmJY2g0jpUia5ZcihSD1eMyYOvr5PUnlVGv6
Sgf+5HSoNrwZTojuQWNPVwSEgWkz4idnlHfi3LbAOkreK5I+RedmK/PlXUJP
erEvHjIuWmAMMLR+WYulY/8wPve4CgBNwapel1ikJHwEZT4P93bVtGDG0oQR
F3j30QoaZBkLWdgcXiRzbhDSoaXtDQmuEK/Hm3oeJ7z/yltMEZaJOctfF6a8
/8E5mvwSBKhxXtcClAg4p9/+9GUeba9nfkX/jYoe3YZvM5NuXoIMUDFQQ1vO
1/2xyxxAAlSyiTovvjGR5ghXg8oXKgaZ9pWbskoUFNYJcILkT4zZvL+vOawe
xPBfebpvr9JxnRQ1BcptTGWZ6NnxdkCx0GDNrNv8K5lZhWGCk6IVQv6wnkX1
kYa2Z/OOgwK8g9bUEfA5SZk1ZLRkdP2qeAjESD4Cdli/9dLCjthahWHb6s4/
kIpwGh6T4Yme3//gCdzAPSzAaK6VL3eg4ikrZLrU4JvWKYatCob9mNDzaN4Q
vq+gKMDnG8RT0NKzwfilvTZgRG7jM5PyohUXwNkdEs6EjzDhT4ABPUEzkVl7
9HXpI+8ICktdBP17BQesIowCHm/R70hu30GsY3AqTLVzIekjffTJBWL+A4As
QQwy/5i972fQp2Ldo7gGDGrpqJKe7dUHCTyUECVISC8pLCW2cbglRuRmCbcU
+mKNakXiqeH9mmIF0cgEAVEhzNlpqS38xArjVx218DPlR9DtnvegoMBiR5Kg
jqBb5fXAXqP/UeRm/pI/ikuaxv1Jmr0hETr7nNa1l0QqnyOqn1cqFcOUUz2n
3HKEePCiyk2kQAaO7aM0LCLgCyZoy6bvr73VF2XtH/QAuhEGIbY6X5BGhezO
KIJxQs54/8jnw8mkvXlaiG9gTKo6oRQNU2c72i/7ycJXrnydaPfZ5QQGdA0S
gA1syj0F/O3RDSmOcCflUZI4WJnllwbQovXpalTz6XgZSrOo8/4vFUz67ObM
n77Ekbi9eDxsd4fNesi6yd9TGSU+9lqDll2eWRLDaOe440lkvkrUE5ySO8QS
c6CZE/Slblno0nR1uhallSsL1FLNkJCGqOhzcq+iE/c+P6Nqg49ous0SdcRH
My906hK3Cml6yL3WzaRawDawxmRNW50Ga7c+rzoVw1d7MaWU0jr2/LMTkVev
bFQXE0+2brn6+kOZR3h5wNb3tvKHQPQl2EPpk4K/06YvvxFvk1wHd9Or5E01
p49b1rB1vLjpOYN2YelkpBntxKH7mrb69ukkWBxrvnYNyn2oGhQgu05t+HPx
j3tO7s0iyWJUclvupMDm3JG+CFRlN7cKNFfF2lNpxQmJSAKx1wMjBuTCs/uW
h97F05KSTIbQbv2/q4AKth9DAQu8VVF4hKaWCmeJFlzbLOiWhOrt930uGG6u
8JMXhs5JN87scqDtP0mgTz6sLT2BRw6Iu6DwvPQdzdZQOAI1lpHam5JAwbEy
nnm3aM0GGAumxgW5lU8mfYtNXPqpyAQxub0FJs+MHcRvBooSNVJdF3LR9omp
jpWSQKg6ttqzvvb8H+TuCGhfmuVgokw3DVfJhljJptIewhgFeJJEjo3bVRYV
vrAPFjgRz+hEhAFtH4sX/OnnGWZDiym/b7DBTNeNyZx4CPEKEmN5octufC+U
ymXq3foMOkGcXJdF3YWJL+Zthb0PxpQtTVkK3ibpe69QbntKzYDASZ6DuQGM
J/3ghvbYvSFkpLe02I7YYtUm5chGgqaAInWnsmI7Q9cMSpB0ts+UdVCxKU7i
kSIewiOYL/KfygtjoIuNKAcX4k4JEd6U3si4ko0oCn7z++RYXNYWwNWOs60l
pc9AiMOsBCbyVQyJU/wZhnOQ0u0Hh8vuRgYO3UD7V70AxbTX9IZwdgmkmrrw
c8HEdsMWT+Qx+tGknlf2UWjTqisQBauRaMSV5e1QOy/fbV9T9AxkvnJZXdbT
vowuP14c1BvWc9wk9Go+F33hyP+ICITecb52ePbvpFIm9QZ4yenPxl59NEDC
42k07nClHmaR/rbDjK74m7adGWR/uCDR6qFZirGNKrdQbj3omKxnk+QisJA2
VnuftOTZIgUIHpn480V5jF/NJDWc8AfbgNbs4wE981o6wTqRgA8y/AVnme9Q
AjR60zhtIKTBv/0zcTQcxe623wXgoFt94umO0nSqRwMXSPd8GhHCWMNkmo8Y
rsPPZG+2ccOwamHBW1nKzOExarGMVFlWSYmAA+puB93D+hnN7k8oRQOmirVw
V/RUReh+VWHj+zc8SjHzwxUtO70kV1Lyn2oGhkUGT4HV/5iq9tjFqVyhl/Ic
O7W2yRTTswKdArAR2KVxFWPxzjdQvRlrf94BUOGUlaegFgZfc+SnqGmL8nuh
S3cEunrgybvz+g0Os+FpzCh1J7I8ZGpyCZxpa6D577ZMSDG3ke5YyXW8/Vaj
611mnFMSTPYrLlJMS0gZaPbUrtfQYGk8BV/4nT2P2p40I7jTMGAHVq7PFCo0
8vVjIvlhi6wGqqRSnD1XX41MnVPvHojKYORO60gg0Ir6j/cGhzfNzJksoPsk
z4TCCyiztcwzPzmr62QQsO2TSGkcIJEakRKs8hroXnzRBvrK+ivER001c2Cz
B3fjLeLu48xW4G7j4O2ygT071G3Kwi0nGWjHsdJr+oQct994Mb/Ytcvq7t//
Nd3lybCqKymUoJPiVgA15Ghnimh04ffYeaNwyikH45dFiahzai+UpdopS+Uw
OuWPVMvc5kKoU33xIgYvD35u/oZeaK3IsJmqQ+v0r0ZqlmKlaOZF2I5XtsDU
2TJ6CNzn3ROSYDF1IKXOzpI0itsnWb0ZJjj8R684yiHij5hulu7B2y6O+7RA
u1cTrt65XTud6SHqDJqVVTQL1F08EiKtpZFDFhc8WVTwt+Nb1yGKaO14oz7e
AGAJlKbJnfALxJ3EypX7UjyRDdH45dMEmFsrWorHYhmwqcn6g5BmQ5mldOm8
rsI/ypelspwXnmSvoOaTRXHlpUWH65pVHD8gKqSia+xLPpkI6vCMieOhWpp7
1LNzq8Z3WQHkCHz3B+QgmE7MEA/tavz5DKftp6ErDSmfw6bt8REO3adUqtcC
VuM0UJyQda58blhlPrHj0dqSIVxdiBNic6H4pdmYUvqKCTzyJlO+1yQ+FYIW
w9PoG8qB/g40BFlbrg28Qi0+MBe2NIyNvzv+I5y7TkR81Cug78y/T/34jV/d
u73uM3cvcgSH9t3Xv9wFIlR4ffU3+Jh4L6Zn1NmA+ptCJtBDKoTRgRMrNpqh
LbK19cy9h6icTPAbfR6kn8mIYfoSuxMRRICxjgKk/RlQlGzE/5NvhRo74EC6
68S9xi0FBuQrE3lzKz4/AO8KHAxm3fV3xHENYduL9zNciODTKzxse0ncK2Hh
/TvVZ48QtXlcaU+XYdxlgyR1Eon7HI698WNwaPRNlMO36D2/d9d0hxKZE/Hz
rQEV+XRDRA+TZurzxRGcJtzrU6CR59QNsG0Xflk/4TXP4PbyYXBFu8rvnWYy
qUH9nVyJgOcwb8RGUgdgE18MhLAAKQ6S3XT9tOEywrQ9pxbMBwS+BTDVojAf
II3x2Iq1XF/mVHsx6fakTIpnLD7wFr1+OK3eKxdh0eFS2T6foFxhPt3JwKNX
uqJnEjGFsNIEu0akiuK4sKuMU9IGa6Mr4Qe/4UvQvgGNorpyAM6dbWdWvkmb
1cjvyr9XlOk94n8GDnM/u2o1s93l5TVqxYkxmoePUASDVkDnarS4wU74EodG
Bm9cgKdEuur4bCOPYXngybzL/6AroaKN3Qd+DbsJpOe7ddxGbkI8hCAUt4Jo
4A7Nb3qIKBss9+57J64hJEsv+Rze9ii0lvQZjY43GIT8LEepKR4fVvW+1Ivs
unkLTNJmkcXcpYcKcBWW9aDG6LMDim+9VF7o0nKH+6t0ISeim0sIWlTtWjq8
QLQZhQu1ELQrfkCtEYAQBnKm4ZRAEqJ3GuCC+1qI0ZMfuH4E/emdK7HhNcbO
J+/T/dA7HifM7zgALsWYqUW3xH61xwyUbz0972Nw8QUZh9KHUUkyakMQ7cdz
8d/S27ru4V1aUsCOXD2wR9bJFlSPyODzwNEe4WYYruRhVJRr3Q8PUtdFUtu9
nS6U6RqmJFlRgszy6lHwkWvqcOiPk1T6v9LICzXTVGXDJkK5lj+eoB9DUflW
H4e66SezMyUhXtZE9zF74u6Rl4czqUN6LEGVsiOnf6p0ChMoG1WcUpsoDXTA
0RANQ4XwSqfIm/bW6qLsBgKFko2QPoSfGxY7p/xydAmdMC1IZicdm3LntqYE
ezxwAw7+LnwNyLGBebqEBWv6yKOA/Clxmrg+ZWhON/bYiA/cF9BhlaRnuhFX
gW3dsa01VYeghCjLxmFFmwx95MmR1qqPD0yjdf9v2CiAsSZ5x4nlUdmj07IY
2XhwrenuG5l5y4+JNaAnmaFeEUXibFYwIZoFVrW4yHbMNTvAQcxSXQscz9RX
IxituP+wbjKGmraE4DZxAjIkPjwibzhS7rEvo2BJ82nxmK8+Gi9pGgshnQHA
0Y91XurrzYMotC6n/saMZerkgIOlLbD0YJ24vqp6myFv9pUoQ+gmfuVOUI3N
qUMPEl7k3SMDRBUcy86VnlhjhqFmB5wYxf4lygzlacFh4tZWv7VFlpKcT9rm
YZ/+WnnnkDfNUcYgQkjmFvq6js5JzBptC3Jqjj8LQPTXZDoDmrmXVmlLHLxu
LT7aavtOnDI43/OdaSINH90Ok1VmBVBUN2ZF/8nmOhH9J7VFQUkLYuPnWw8H
615doyQ4NErF2Td1IGsMODYYPoAzfLpasZq1ugP7kc5WeTDvA7vi68dLlJev
Gp+R5og8bDeLo3Nf20M1CPqUqxFCyyhqdcThPlnlZzxk+sy6FVB8brmPver+
x6874r96AR47DiHfa7L+tIa0K0qDqnYnXbxukVNyPDqWNUyqdgy1tg83zfQL
0rBTzNfZ1zuKiS3gspAv/XV+daXuRY9MCHASPQFM2wKj5cCc20uLnmZh1f0c
hes8IpCyFhTzitiNLN8RzzkmXBBC7BMYLapjP+vlrMlX3wOvQ9igO8LTOlje
oDqhZbIuytEkBqROyyZgYFoM9jnpbg9zspZf5MM/A4tLcRUB4TVwAhrG6YFI
iw9jTylwa837Khrbvr2w6VhTbjOjdv78HVfmfD7IUteZqaRmijSWMJjSKKcJ
JKvw8NdosxHxMLDgl09PCUHjlE6pG8a37OA9BCYxNMmV1Mumg1tvYWyAT+V7
DYxP6rsCs3XD8TFBLsWhV1X+a3NtYe/nAVpvbFG7F5VmQ2cAlAHewIyD+lto
lsxlJxaPkmjcsibcrhZjTE2U6iMZQE/N8a5apzt//e1B5rncGW0lq30lBANc
ABKsvsqrsXgvW5uhdMo6F7A7kRarIUyqVFFO54cq3u+wuTxBOyt9dJLkhPvE
6Nu/rKZQZmTsR7AyVWHGh0FMlJM90HQBPvD1TXTSFfdImosPqox/Zfx7tcHY
M5lGqSftJKDj0FHoCIPxQwch5kKalNIUZUQDbZnEgEqPEczimUCHloxs5U6q
tSxt5PGBQHVQampOaZsQgVv+wC7RlBqafh6LG5GGizzjzqVU6weZYjSIvxdc
7Nv8UsgpQkXtF0Yz4jIJkadzINz8rq0VyEEOHRl0cR8kFZk8DhdtRHMW1iow
hRYfNb0tBoeSqWaCL6JYIluTwjlbfONEIsMUes5LeKTRxJR35E5XrBhbN4Lv
2BvCm2UAfY/8YdLGM4E1QplTW3Ch0GqrlaX8hUNm9942PSXVH5M9NL+neL27
FwRpyBeQQPvRKLEthqjSZo8gkOgPrkIr4AGIe86EhqHrXBJjiM0P/UPUwTUu
coTwS1UAF+UF8hmsKA8yaR8pUm/MTm7f420xi8FwUR7e3svCpeojO0c1jxQp
0+JjFTHANXw052NsvU2VE256syq8X9UMM85xXg/DtYiXaYU+eD0YPepmscht
nRg9SwXw3gjKT9XLFk/8UQGALwXDub20uBOySKh8ADTAiQ0z/EAKRXCswyiH
32qOjYJX2YT2LMP8jCJyKMyeYox4YEELJ8r4ZHnX7YeUrUhnk0MpxkmvaWrm
lg9XSsTp+izNoNC/xmnS583e6IfDM4MUPz9p9T3EZjXRhkehoiWguC2pLvm0
MYLwSzVIMTaVu9eJbLajDRQxsp8i/vDGgJyHvUTwnYohqf4Fo75g7LDqkNjq
VeQPLaZkOcnucdVSMjnc+dD47rSmP1PMYKW3zVKM2Ce9GK6eR8qm0z+nikAR
wjtRy/G4dDOuhLVm5nIqQQ31Ezr/egpa9Rv+Km3/e/q6Sxa1FUae441kHtka
jd7J/vy2UWciPg9DUC/v+Uptk5111OgYtK+gMvoon+0/iKeYi8mlt7pcJF8J
80C1Abib0qq0kwZvx1QJLoQepCTbxbf6ZZTVWYi7kJaOR2/SH13JCnIvIxhv
VnZQwtGlVrYjd8t+W1rKvjNKiCk5bnzTMPpySrCDI0ZvmFGTyvPih1cedcC8
TMPSielEOQ5OZ4lvNCDgz6mDNAaC//SRU3s6jYIU9htR103VH1/UnkvIpYLg
V3hetjIbOxJI6goRm9I5V8+txLXlji2AfTSg9D5NGrTbU+McLcm51wRYbhHq
IHlodcESr8w+CUO9UQytNA0R1vRyFQpefDso349GA7HWfSx6g6G2ltfq7Efj
NepLEelJkcx2ERm24Gxq0BHN8iR7k4pud0VuonheohN1VSiDKHS26qZtKBpd
rP4DPzMfOFnmWiCm8EnAs8/x5va46hqC8RNMomJfq2oxE/ONmnsUJHbzHWY5
/V0VCvlgZb/ynNrUyZDtvmJBqmJ3xdGSZa5zfQMqby1KPLnhl0xiJBozHSHM
Bvj0c2Adz4Vqw78pWhsEGHKiWdUt1u7Zi2nZvRQ2itJVqPx/s50r3KhiJm1I
gCW2gFmTDVLM5Po9cMdFU9ORKz48APtNZjTGghz0qimfr1toe10g8OcsOEXb
/K8s8tdzD8urcSGqW2zhOQjoYPwtvaT5oFzdUOTIGtv5KOz4+IbctymX4rmQ
OQBK3UsgqMfAP8ICbLtYwhKP+zVPV8yNpZiWQKN0oRaL2fZ4sHJPrhG8BZqw
dbAr4pz0T5DcpDcdNR21RDpYO4XCn+AEZWe314JQGTkQsV2awnXkMDeQeBi+
ntNopB49e62bz+zQaEDpG+jjzawqOyIGoj1NWFBb4g5MZVkULLxc/C+89x1Q
g1xln8w8

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+nvfweU9wbtSegp454nVuLlKbkeCn8Hp8Uxhznrz1dxa0gPhspblJlf3O7FxEvrtCP+obhY8DIHpr7eGhaIS1IgHHXDaXHEVE1sNM/AbaMLAbHhSxW0En6UXi0a9ao+lmORn/cOEB6s3oJ8JParsg7l6fV+Qw6nabG2DFfLkpKTjTSxVHcpgfMD/P1mf5RIyXsU7VkqXH+5XaQhTbUfbwxVDDZH0PQxoR4zFe7Flh3UNoT3fwX2gSGbHd0kRXv5isJr5dZk81EyL4fywi/o59dHni+8pPV5kEC3ZZDG/z8Z72EPaRP2pzM9nWOlUoXKzQdPO4JvEZSrVdnK/dHskATcfPe6In2F/TlTC8QgJY85CZBVHUIVvDEzKzh5tQaqQIHjM+qErxEquK5fdHu3OiK4W7TPxnlRAEqDQj5ovI/Tg/vzgIIJOHvqDt3b3U3dKWGETAXmSDfg71Q8OUvSjOPMVSLvDWe3DpaGzuqVNsshcMVj8TIO0lhoKX6ZBbWWQLLriArDW/JnMhio0RuqolP+IA3eC55yup230VGiDIKzp8GOSTgO/ILsFlNgylyuIEOl3zAYQVJ4cd5Qg8Tw9VlLBHyZQWj9Cuj8fxULginDv9oDtYxUxJdJQI4MYJv2PzBaQAdu0J625HukWhbflzYExLjaltWde88E0uDxsGqtSqfdCUvdh+xMk8ONALWaJwKUQAO/ZbwiuZ0GMadNn7YTmEuxqP2MFm4cXBV0IGJvbhrCwic6s5sr51AGlCcWQUsVDVvGbBahg/MaV6CzPoo/"
`endif