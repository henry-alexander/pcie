// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cgcEAor6/buT58+FE8k6scxKFl4NJMyhNolaXMl+sk0VtG0RQq0eS2VVc51k
SAvtKvMpnnrcKwHf39TRzjYgKrm7PFq5zD91KZE8jXyD4GZyWu07+zXV1C1m
1B/HhUDVYHialnrfJzeuJSh+Gz16f1Su/YkwNgHevYlmd/yJo408mdUWkweV
ZXGUTaQjb3eT4Vqoc2C/4CrxGtcSbLJbKX/xDZHXXTt5e3L/2j7iFpTT2ja8
4RPh7K/NqrPIP0AQZAnUPjIsWWn5v41Oav1kPBSfakkxJBcWT3CUoZQ/fMmx
cF7R4JfVKcklsDhMNyUdzm6Sh6wjWtpG3hLWzvITVQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IVLYI0j3D0UYVHuVx7XUeXl35Eec7PCYuWFgNrPJY4G7BFDAjmuDvSjDp2KS
BquWo+isj1eabBVeywR7TkJ1E1mKqwhG7IkUTUDHJrvLxsfi8XY6SHkHm2vk
WH7YEEQq48/3W8ieJpNykT3vjKBHJcG1bH2vU9ydqVtF5lB3keTr/0wQcHXN
NYePfopn8zgnVctj0HxFOXdQwqkyQAuLnhS9h8Oilcj1wM6O/1PtaDHKrQ08
WU9Mx8E9VzveQXskQrnMYV+cPyzGTrYkuUNyWUlQ+JysQo6YpJema7AfU4Op
Mnh1mgw00nG6kOj9moY+J79lpRkwo0m8F1ptKOZQcg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
PprM4U/zh7V6T6Q0FtLvZlYyNr8MEidfN/Wfve8mg4Ou+HF9B2ehE4oEKHfO
o0nAYI0GXUMmDjI9bzQFshVWFDuAhbJIYfecbAXx0xvZOJP8JiUIli4bVU/P
u73wazs/CKlAgTGQmDX28Vn9vrtVm7eZK4fDU2aU/IUUmiS8veb9i1dL7u1k
hAVzHpEfznvhDbX/YNmIxIkwaZTpdt5AUcRmWCjmJ1IDhi/ivpcunYGV17N7
wPwEMdSEShdRFD2zPPw8hZoBnO+qP8nHARqtd5qsiTtSYGYpWpJLcK1kNeHJ
f4q3R6rCJEl+440eT0/PFfDeYcUvmPELczgYyJfwlw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
j00C+IFem1K9lNQbYww62QMeI1kAt8+4pyYm3Qt5JU/+XtlYjnNmDisnEigi
5XTnCxsJ9W3KmXuvKbGGDpm8BJJjCAblHplZUKsnR2wt/SD1NFxjre2TPZoq
6k6XtQHSYv6DttSiYm6AlBdm3m8QOxInEVCf8BSueAsjXur/Vos=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eqMb3Rtf3V9/YJLbi8WYe0o+pStBiqu2g6XBLN2DyKudA66l2HC0BToIFUda
YzKk9BaBrmCuNdZKvXgqm3eYEfjqSuiHAhxP55VJI+GT40H7NCNS+RYIuuQT
ql1XirK/9ma2WjiQgCQuTJTKkHBfn8drtvab6hLcvVGAWHyDh1Z/Sqxf+Obc
TDE6QI6GDB3Eb1P+Sc4r7zikfjuHZ+UNZKt6QcIoUn7JDTIZJbbGjfzJX312
bzZ/2xlva8QERlvCeXV/lmMmQBfaw7cVk1fL8IhOCakm/FGvMzUN5CAwbO3J
Ffm8lzcZjwpaJEE/+WNmG9V3hLKjDO4Qkv99/AwgvxNxJFW2jTnOplDuAGr2
lK6hlttxzQgy/XHXVYqaWuqlfQl7TQENZCycZHIcvvRUM1WJ5zQ1j4ttHhOL
annz2n6Leyekz0m0aTmHBCuyyHdeufCH8cxqdvltV4el6LnzaEtBIuXfdmDb
/Sw7ZHbGZrGt/Dr+obIwlpO5D0j+Zp3k


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
D9FsKK1R8Ot4WUEnoQhsIFdnYMK1YHVHkTF71YzQXE62+ozODWybuhuKo8eN
hCfZDHb66jhrx2D4MVllSlWcXAH9qnH9aDE25pXKy8zlK8j/0RLs/EeCJMz+
6OYKK7G/9TeYj7+U7biWrbVS6107lmX7+4a6vO5m6sgy4fnRtUU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
lXFw6NElFaoZpcGUux3fe1qg1Jjfo09xtpTIwP7UDHtV5oKjjLNDPya7gft4
uLhxAj5sH2w3shw3zuXRJrayhzLGjVNCLA9eHyfDINlaCa38oUpl+JXvnNdO
NbnWRtRs1mco2vwXd4X0qOkL5hWGj38RqtRjkMtUHZvRAcYDs10=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8768)
`pragma protect data_block
UB1oh9VRqpZ32z+aevkG+Q9ZNblnD8sMbGAqbojAiEnHOFWcG5AH8TapRytF
IhqdfWrbiSDVKjUUxSqB9MsaF47+a6Kwj8z0LyvTjioO6Ix1tU2LL7khWjNp
PArohCpZLyRZ5x8geAvxFhvDNBQpNoMa7wi0Y4ybbydct2sAJG0+4dx3SLPx
QEyPNANLYKYWzK/WbK2NT/KbAjXxwcmOLF3osZpOSRx0Oqv/6c0ss0E65++8
GUuAfJxRyVkDkzfEZ/Se18u52Mb1wHiBBoN+EdP7RNs2Q2cQI5+oaYxBNPRk
QDThFfO7kkECIFKnIaOVa4bPGKRgDUwIzVRHIbILYZvo4TQwGzIQlqQOEysm
h6uzNC4Sax8MqGLO1VMbW/qLpcSOXyTRNT57xnAePO4wUDbbS49yqloAscYE
4jkg//rQeOfQ94tPrfp5v/Z6EUSD6gg73s6Fa7pJuUHndqBd8yS+H8szTvT1
X+9JgMe032w01zAl/OaH4kc3wStzIwD+iYpRbl33hPOynAzLdm5rZpu8+uLR
kr8IyPJHKLdCbh1nA1rtIltUHlFVOFD71pvHPWcaAUNcD+R8rK/hZXqLXSfb
ciJVI3eQfjCu4SArusnAdC9OIo8s5ABGgiCMOoHNJ5pom9V4JwLTQpX4mg+L
twaf0UWOZhV7X3QsifPEyU5HDb6yB0AcAxIwrNVO7UWN/oNhqATk/wghr/sH
jmOuZC186GSw0H/hqWUi+P3LlvsY6aociUdGStWwYNN4ANq3fPoWZqqKpV0G
YFSsRgMFOXnf707zfqANnKrAtmlUNeazVPa0NXh2k/sLA2z5IDPJRDXuqKs7
F7j3RTIwTCnJEAuUmC4XbnEqhGJPhr2ZaGwANKlk30jiFQXvEB1cn++eF1QD
t3CDvHhXcc6uRWuwnaJe9n1uOaQBy5DEcOWdktOI0fFsJWuqDIxN2yrUEK/d
7qXd76lAMjEPQm7S6h+NUJ3oVgOsfYh3I6iOQfCiT7cEcWnPr7tK4SNBE576
eJb6+d04MoITrQO35DUR+x70aV0yVYEmJF7UJGfBZb2cGNXI1YblaGPtUvV+
e8ecAG+K80wcujilNlAQB5X6g7Axm1EJWbRzpM3jKcBbw9dKqhwV6+qXr/Uj
uxlJ+h00+uM7nBkhyUuKFg2w7VvDLfFI1agBnY270kPCls0gJbA5b2GiPCla
3Rv/zGF4pT/uujFwceQy7Yoy0MfK3rUDBpo4EWKrM7Ju7eA66tFbcb9/yYrW
xj6bvIkHd1wCggK928cxwfTl78B28nVwdJhte5y2HIxcsPsjNy+5/MFiA+nt
MfiVu6F2PUHzZ2P3l+TZM6RkfyxOSBBPIhMqR7nSm8X0wHufaktnMet4tHtc
7VHoIW1nqDPMiw9vOeCB2ECQYRDhJsaIgfw6lk9TujKvpi8N0oz3thEMUEEH
M8Zp/BVIqKAejBJifYjuYUFRvjbRHj2BpIoO0zHiFdpWpbmj83OpJccosY+n
tzgpM0T7jOtn60n9BiqcDG7ZxoEsFnsa6p8Qq9ZpxUEydM2UyiOWx0TwAe4a
yb7ar8rbMd0VBVcUJsMXXzpF+Brd6GtJJaPmCDKfBVGjb9epttPVDDFN10IN
yH7swPe7/d3GVSFIcCYC612P509uJ0lr0vj3vlpcpmD6Y7MbCloXQIgbK46K
tDdAwL2owEH5QQGeS0xioPqeXNJq9QDNZUzLOohdXvKs7y9cqMFTguIoTCSO
h+CQjhjRjxjvICHhzb1fSBNP5k9AFldLLEwrdFJHTOmDzY14/76/s/QNEuJr
OGsfQx8fHP37lnlO/NKRBz+PkNAcYQb4cRDiLgqwxSOGHHFqEZB93rlTnMsl
ue5drUxwLkgVkHZgflbi96UBjYHYYFgUXvKWPMMWb5XzwaNFYGWyhGPn/Aym
4zS0IwOT6TrwIimnQfQyYUI1zkb2uIUFDZqHo+vBZisAif3iqahpY/q28A3y
oZuDowFJ1Pz/wbWx7x87OG3QmEQ8mV9ZwLmIDJW3zosslYHGsa9qucw77b4P
FwiG9adTLh7uoH4VH2C7ELKwli4kbSv54CTk2bjZFuSkTnQI5w2wiP1A+oJp
cYdRz+mQ6gOkG65eCXspXNSzy25zZ4MGbvwZisqKUKxlMI9jrQCslAXgF5QQ
8F9shVwiRJkMcY3lJktqohFWLpFCxrBHJLysbU0tEobK+sTX2Mb85v8Tw5lM
5r45kzwvBUwKMrPR5XFWEp56YoIpLGVxAouwUsCS5c/q1ed79hUlvPBsUucF
tW4LBYINIREq5WQrruk9WooAhm/IlvGjfi+eCBqSDOxYZLpuFf6LkUPjOwM3
xuTnEIT4jooHkeF4Fr5Ocl3Hqi9MZMrnOzMxITgUaA7mjotiVoeihYRV5UZb
pUOs5A1lcqzOD1XZQVNgplJQP4FXGxRnJgh8zqr3Wi3evUjti6t6HzHNS+bj
P6pjv10fb89dbXIttWUJ0oo91rrd8G87KvGmGEChmAGLknuVuaaFCkfdJSX6
IWDW0xLtBnb0Sh3zPKtWf71mgZQxpiq2e46iV1Y1BYoaWYFU2G3dLS9z74pc
Jgu1cIKVa4dL+VdGvABi7HkxYVs2JjNjkota098O1cHSECO/yJdbwRe21SMk
e/xtUtW25c2P+2YyYf0Ch55XCIF/3fulT1jd/upwnPuHtTBgBspQx3zG7Kv4
fiRENVUPaFrjoYQ385/40SF4glO7C6YTbfRa287DJCa0jsYg/+gKvcJREAgp
kL4aO4IYa0x9tb2ckgSsI6PMAGoHFYBY3R2wfcAFL5sPFcA2iB/UAcbh+Y+M
hG2QyxSNAprTYr/QcQEvw4Lui3jei2wV3n6qkBrNiqBZFXrWDF+hMOKqFJob
sUAV5xx2MUZ+X3ip8L9rG7Yu3NmXnxdtbhRtoutVUS88NJjEKYIQZvg27eZG
DH4SHfhca3hc8ACiKHm/47DhnRxN2PsB7oFZ1piCSsM251veNbNdFQWxcNUM
PvW7NeS9T8iJxgVG94A/AB7OLWEBbH+BoVC1UV6bmMvLeBIMTLDjH4PkqrQ9
OPLCeVNF/4AiVptuAz4bqh0vkup4DxnMfpy5dpzLs8y1VMgc/7SscwTD/iPf
fjeQbggmC/2lsR7hiXFe81hPWzCebRpnVEp2QPMQWdEVp46ziGOQJwBgtiMT
NfoaF0N3mhYlQt7nlVjHX+EwSOc1A85QFQGm56odYiM4wIgP7RdqtBupIDg7
F6avrqrXs4ZBSYSE+DySZ8+rWyMzlomr7kw1XhluYckS0sj2a1lNLNhDSWj+
ML6BpIEmEqkn3K3gwk3ZbqzCRG8/OqdWip+mctvcD/7A3PS/GhySSnluRec5
HguIskug4JTfGXjP6tVghZxAtTQuTUxm5JFNFwIfd4nlbiAxD9ovi1Yrz71c
74xww+2vRj7n65dE82Hn60+R5O4B2172ypaavL2lvLoc4P3pTgqsTLVlqfbs
ITdileuuU0DSjI6zSiE6G3YnWi/1yeMUIho5DT1FnRjggSVSZwDkmqD94ssx
aKCke3yWpyh9aIK667ggX0Et1bmurJA6YwPHvwYCn616mmoTNanCNMu/kQBB
/eT2NRH3q7gSsHSTtwEbDXuUBT2H1rw0XjyREJMw1BKuN7DITOTWIqbpAvtM
TX825wLJOP9sbdUy1mUL915QvqvmLPw90HlauvsmSghUGI8CCvrvBiA/wJUY
gvt5Pa0Il2CoCr1jT4KMpCatkLxo1CK6GYJRr7yOxjSS5JwD2dCwAfm0Wijv
M3ALrOXGJSO+x4VMD4/c8ytWeKo7htL6Cpyo9S+MozqLHZvo0j0Bntc1qdPv
7KIxfBXgwv6wUAFHR5r5HEgcvRNbC7da07+yn8cN3JeKdvhkyC3Qs/u64x50
H/Osb4G72YJlECe6p1mA0hYsImAoRIkJoYtW498rEZaIzMEiaN2tfCN8P/f4
AWa+/4UXVywyss0NekH8iE8ytkKLInJX9dP7MAz3CquzwbHEvkhkjnmW/8Bv
SiPCR0nLtA97YOIm5Fzqzhel8hGQHCAPixptXxSrkIwcItuqsd51CHbhKLoa
DuLFSOB5MJp3q0pqUVllTy9rAhxJvwgAgKncGJE0CL2WMWayQtn43RbtctBQ
bGIt0NtoQCZ0RF9LW4YV9qtrdEk6SOcr/baSEN330ZDVtQV6LioXpj9GbMpd
R33RS9WITb9am46nyQ9sG3EAFZZkeZZApASWiVzo8ep8NLG6RQ6vMAwVm1xn
l6tK1dClVJ7r2Co6/DIxFlESzAfPnOiGKGn16/5DE6O/oa7AbMStVOkkTBAl
oyt1DYAjNuohMLYhcq4suB3udC0d+4Y1jp3p5W0VcCKSC+yCLDtCvwVMWNkx
+8YthvRhT1Fj7YZh7J9Kji3nGtjUaO9RtjhmpOiD1OIbw+z/+1CbL+eAB64l
CSVWx9OVSp0d0lYuF7ZueagF+MHqikkiOXV/Df17VmiIl/2ILXp4os2RfQaq
sjruFeS2G+u+pIASaO6agVm4IqQKDMZz36G7mMZdfqEj+sMxz+3jP//Ns8/1
/26Pi7MJx5awkyOFQ9ngw9pweadVrWHU5j6Y+jPdnxwnNn1MOT6WzVQPEZ4G
S1jPPhVA9qOmslJiC54WQZ/kaihtZjLhvF/VgdmEjwxI0aP3ypZHugqOaNB6
K6sBGgPy46E6D6WK4png+PqOuiOfW6LTZsrJ/BIG1HHrs9roo33j2/4q3zVL
1pSN0cp3R3UwhV4I71H5wF33nkArDQWjqHuAWBPSYr5E9W4g+xbk/ikH6fLk
d0yi/vDCi/PpJ9Xcg4Sl19zm0yQEeWNpk8cCfrlydB2mjpaldsNRVe2Y3eqa
2Bng3tQOIqQCF8KIecU5JHbF/JZ7SZUk57UsurA2KwRGu0w6hfcnTMDrj/T8
qMB4JSFOKE/Wa+8CplrnfQfaH8bfmMXE69H1MehZrt3mvCJa38b5sNvefaJ8
ivLTXNnCwkhJqdh2n6Yspwb/8VE+0P4aPmAdwDPakBOIxp1uRml0o0nnO+62
gyIne7FTa7VLDpynbj3/C7pDBqU5sH5DrYKJZhKetUEMtxTQvtPH75YAa1+O
BXE5FMrfCIpWYyczwBQzTTGlG7BaZloXG9bKm06IpSQLNjmbmG0WxCKaE7GA
cRp6xWnAHCCPPmFlwLBoTlH3MLyTprTRChzi0txk+OSwyY6aMKUzpk0hYHML
mBe9ya0/vPWEojPmE888RozYttI+Qu2VtR04ErCa1YimYqKzC4z+N65CXyqC
+hdnHTgxuiq/XfWYiQb8yPBVkxNM7dtcXouqkVvPVOp8vWhOFqnnfSbrEjIh
OtdGw520USFwz7tiX5OQc5/LypMTVHsLHl0nOlH07AK0agoDFa+AGXtaXZjI
osvnynEJ4vNy31RsDU8KoaIW+IsqhvK4QIsKv8pGpfvm2/tBFHN3+WFvVmUD
l43bXAzP6IA+UR285N0haKy1zdtfXOTEdCRfcOn+7RiEkQIMX6HIBcWJuEDm
ffv+4Iuq/DqmcXwrR6XXf5X2q1Uz9MajCfZU7gESPRNMJSciw3No6ZDyldlo
OsK2V/84WvThFzGtrfd6TVjoONU04RRhC4MwX13xiLE90HkQca0RkFEg/X7/
hCfUCCPeS7UyY89DlhYp3x3k9y6sO8v7yQwLjVArlG1K6F8ODeBeVN5uVn11
EGFNv7+oJotbUS5auy96Yeh2SkdnOKr4F4nsa1c76z+n8oq0lOAAvRwMVung
IQ+I+Ih8tSb58GcRmwzl/322787NHEhiHclmNJhCx/AGRbcnpRbLzlOROl2x
0KrPK6cmt1UPt1fdlcrgPZOMma4Usf47AOkOCwineGQclp0bSVfSNZKBzPbk
TOibEPBgqzjww5MSbrMkCgvU4o9Fpkmvb0kw64KEoc1ZpHetsJj0Pfn8qBZ5
2TCTx6SbZMSWP2II2f4ln8vJFy627jelgYZcsO5HKUCR8aKSYXYzRkx2ni28
CnNLc5Bdxiqyibn1HM2VizhmKXv4Ig87Dinf+JgnwmrkdNZHU30l7ubhpeN7
0vNvGRec8bvKUYu8U2Ar97gDbNAn1+eWDVTw6rIG6y/NTAAhrDvEbhjveahf
CLMzvyl0wjj7yupcJUuMVOifwaFcyWr96L9H35NaSTduOKghbplpqTHDF5tk
uIC7CiJvI9hoQfwzkP3gy4RqEdNGmBKmyCp8rB75RbfBf+T6eftpQ6OsNTmE
7ngsrmyjz88WMgM3V4Xp0BSgqZMmhn6rVQ8bA6AW9wrRl4WDOggygLMjRYjS
aFtS2AvY0fmlQKGnz8Cl9vnrykNQGHNHRhQ93isMq9TStSXd60/gPg4EPiCc
Z4TYcNIUiUFU5OwAr1yJSxAXHmtT82Ovhz3IG2st/fUEZZ3JVvlpadVo5Sog
Ag0oN3z+Iy6mEXLiXlmHdhqD7mj2nlYnndSTJ8NHHG8M9IRfWu7TLetqUXuu
kq6w07R2F+8w+AFSPFkWwxFSQGRmBvx6TyjEjsvow5qvnD/5WzFrmMwpdg5l
6Ut4GgfLg/O4asEKIgyMQlYli+escuyjCRA2Cf+YgKYP1hUu0f8H5gwBHfua
NCkfj0VNrGT4xigzB8rU1WHKt1FtN79FW7OVPFhM+nKS9zgblLRH2dQfvm5L
NeESSsGFg6QbNf/hxrWAPGvep1T2/74Y+nenN8HyFZ+cMotz/v7XB6nHWwgX
3r6YRVXbyjp8o2+8qOA50HPVTMfHOzEVcKBNgsPIjKcDGgVrqP2urPhTd3C5
dCnwR59K4B0DvBKZlAn5fgusUFF/rcl7YyKhke6lJigcaoCxVZMMdkH1sAqu
MyISmWOGNT6fyvHjDUFEWiYHaEGCYWp25OsDWm3WWY63eFJyM2cIZznpxbg8
6/2t8CI6RNK/0wlO/m/YeuXlNRPkmGVo/Dgea67rCjKXv/1LuhIU47TNht7s
dUzxjI1iNjwHodVK7thkLc/E8pIeL+EjAXwmJ0XAg9rAJJqr+EEHDToj6Rey
hz7vk/zlervgLwZgsZ48rHfRCxOI6gZ1w39H4dXN0N6qNoYqb7I920akk2Zk
gNMT0l6cUQ6DEQFGkPiV+M+UV0Q/PkJz4xmNBu18csRxR4jZFNbwRGW/GSlE
KUyKln0i4ki2A7Pys576SILUD7PxhjkeCQCgpwcXVbGLC/y7RR53P6/n2nxI
1rzUjKJsyjnJKHXTDE/39gLw/dw453J1GH6oJjjL2EWaRRcFdA0to0cbP9o0
u5InP1Jz8qnh/y45jzczmI7xdpxyg11/fpMXkEjvr2kZbhzW/6C5/UcX5yyo
K8RCuN8BHkCfaniS1SARgmL7esFzW4JbDEW4EHX8F0Ra2FfU6O04mUTBDbNV
m2fZNcmZQqw2oGeUvj0tfCT5+35XMpkPArDKYEiIPyIu3uk2pPdFRxoGVpsc
iWjxPomPEjRxXLQosu3jW7O4k65TyuPIGz5ktcDANIutSQFlq9ta/iAzN72R
8yFqCldOceDEUExmZWGC0UQKXthPjVrjseNufEP7HrtuXPhZpgdDhU69n42T
fZ6Jt4sDkWDku5X9KuaXQTugRhikdTckoZmyDl09MeJBw+NJS6Vpw1D5P4Sw
d4lFFnvRrhjPgpGTDTQCrZMw5XHRVp393QndSe4BdRph218WaZYQoWotQAcZ
UGz+QPg6ad85zWL/cJm3QSeBDMNX8WwbL9fAowarq4Pa3rg3iU6fpJQSkLUK
PCOjgbEImfzY6yOEMeJ2reYf+oA7ilLeW+PRdOnFmvnsyOxErj+k36vELDWR
xwfa3CD6VKqfHnGjv3wGzVfSrDxGE9unJcEIAf3NccgNZTd0ben1zpl9hrlX
VCUPa+JVYOiE1z3nfd10pSHSXdGFpeqk3CEDeSq9qyMYXzYJpVmiLutpe2lx
O2ciTQL2khP+fBm7LaV56T81q/cQPrn0SBL8erSi4T/DgZNORdSErmV841KR
ShzFZBpU9gIYoZia8nzU1gB6BmagQCWxwaVhFengIDbzpn4+DEDDgjWo/Q6j
wk00+YOfk6QlPqYlbjViX+sN6++wtTXqM+V5kLeEqjBAtLYMI/sI2MtjNbWi
4XucetRUCTnSMWze79hymgUWxOLOv/VcuUyR6AwqfBZ8KPMMdebD6KZ0UmJS
c2m1eaO5sDR305QIaXbagnaSf7fXj6QffBOoQ1UWDLsCPJMh15LUxfm7F2EE
R5SSDhOJXrXwDvPj7/3W8DRW0A74QvLVONs06j5NA6jumVlXWTmbNTy41h7P
YHwElh/xBRCra14Jyl389tk35N+x5BpPKfhKPAjIx1w19bLuWB98XDC+K8Wp
rq6lVKi7xzu32qBvhuCgUHqAbhwdR+KFLa6M0WZTD5GUid+dgG1o4W2WiaAw
0KcIXpAcfskGev0nqpsL0teUuynk9SFjRxFX2ngO2baisyEdLtBRlLfY5OKT
dal+Tl3Eruks5Vl4V4HU/B/CDDTco0glffnsysvhU+oGW9POPgiEHSJE3f0z
qeWvLsqRxrYllJe7sv0v9b35aV5zDWWK/+AulOEq/dJxIkCyt2Hwd0iKuVEc
/43hS/gRsOacwaznmXhGafpu1zguHFQNOVQ6yUt+csZXh7kdp2WX2bs5bim0
lcQFcpzo8VadvWCMkhL/Sel4TxViaLf750EVgygdCegHzcq648za/jUOln5F
w4qxepzRuRI6u65pbuWL9hjZngJd0Dj3NZzyZNMSuKtyODYtqylRl0AnoqGu
nQCqqmoLvMltSGzQm7Fn0Uh77JM3xrHHYgPJD4NkRLMPwzSS6VEDlZAxEmvo
s/luQsKq0KVOUCeaXvMPiREXX543CRtaAR+Ol2DWGBcazb6bYWdmY2TCStWf
rYXdW4wa+DwuWX+PlpuqHfrXgkM7ClIj5NdlSF/HUgGSFMxWURRH1+oi2E1d
S1RMdcS76A4Ep5Btr3RpMg6gTF/StgNdskfGCZKq5U8qKHmUoJ0ab3nEtXyr
wo93ZCETJGvxJ3/CQCYDxVMrRmJmbxcFpCtSL6hCC2bopF/JqDIQKv+0GjYY
TaLxMwHedcKAwdjzLMYcOz7uvF0ckxWUXGbxLBmM+1PNPxMo5EIdc6Z+Fl5p
XABo8UnG7OLtIbQh5+4Kxxb1bbD+cUWapFgB0rNd2Q5qx/w0NbexQJKGjys+
YbuztU2hM/yWUS2CTyxGltqWnZiGjzGh6mcmaswo+6ru/sSwy8jK1P/utHaa
yHQ+7kXJFRTq4fLRJOG2Q/KKUt3kNBGPuZhDpb/yXcgNr1Ok+D2s6QAOO+yQ
85J8nFtRk/6+f98XvymECgdUUoL26B7hCpvVkzr1GiZQ2OkyiggGwbcpeYgE
Oq4O8JDH/6VQzBeP/NpfUFUYYV90E6VMvMQmvA6iHVSKu9Cs410SlA7Sdx4Y
vqm+1j0JF71xlTtLpC766tc4iXQ1NHeHJ+txIGCe+zp+GybIxQOi3UP+HYy5
J9sPuau3gpKpIpd3aPkuye8AjzftukW/3BAxTl5tqD41Nara9ZtsklDpYkcb
pISoHxpYgukrhLUYYRjyjmpwkwgDXVMMG+nUZmU3NGGFsfmQ55fUj6ZEbrJX
kyah/h24eq3iTjmBmbhCvz/7PAiq2RjjmjCeB6SJSb8iho7FpvjEF9avr8Hu
qKoe5da3q3Lg5OiRDuUgq55pLOTEK+01iL9X4aZMtzP3gizlPalU8uUp8pHM
rJPZPgtWHpQQiKCD6FCAjpuevsf2PWsiOW0qLvkWbh+jSM38v/cUJvtr3rA0
7dB8I8PuVzzrSoOISGc7PbYEntdeqbY1MciqBqUd1k9Z3suGLNXE1nL0U+w/
ewDDDck9Qq7CJ6RleBR5+hkzyhQw6Z0EQ2dkVdsARGQJ720XlT12/g3Fhphe
UUJkxkaKstEpR6+BOXVWHQnTOys3b6ZkrsSdtFZEgrvvGMOOmKdEByMkj1hS
jBOl0aMQpoNWkypiM16zFW3PN/70HljOf+UN9spUY+yrQlo1XVcsKP7jBjfO
mPPBJdwtjpGxbY15gJ+21iibU698qPhvrH3eBgDRM8mJAlMrSlObGCjqg7ph
D+4C3/5Q+HwWBqat4/RY+WBCe7YcnSBOGozaaE7s3dDHci5FhRoMygAUzGnO
S5tWpuUMOkVfIfX2zQaSRzHIBfciNPMg5ZOqLeggKgkmynAhVht5AlwAVNeQ
Hfp7iOn9UeCRfCTsDprdew29UaMPmfV9p4Mr5XgIKiXn0h1jKccVtgL36Ls8
1orxA94K0nQ5wrj6Y4v+C6FxFuf9Zv4RgZy0OrFPY4vrgUm4Yp2gf2GJU8pz
GPhp37yV8gKTvQFKpWJZZS+d7+V3UtQNUl+Fbrmp9i5sUlY/KKj6FUilIGX1
Iw8uwz5J5RoALDHZ6dkTdw+FGwQEnRDLzRDSwkKEkUh5tRjOvD+pMftyENBt
jvVoxHhVGmBb4uAC1gSvM3g95wrxD9pB8kE28bvFfTRsEBHjYBq77yfPXbqj
JzoqtQXyUs41UCIfbhGRseJuLuVBCx7L+TIZYdHtcwug9vPdv3WwpJUEIXLc
40nbQC52ROSqrmD1graoFgm/1+0aBbmu8DRixUItaRolemaGREIn80F2Q3F5
absrFS65byW3P0V6OII6Pd91xqy4IMnksH8YyCtLOnoM+u/p5HGWqygTwj4G
CYysTc2pRzo7tEpnc5bsYr4Q+W11fpkkJNEqC76KB3JRylt/Sn93VvtWiAJT
g7XW+OPo/jlkg+pYfZ1cNfRkjlf5eG4nH5IlDHpA3cd/QFKSwV+keBSza8GL
o6uTs37leS6OeNCPsTs+fsAeKIYIqOhHCHX41WjaJnhKwa7Gh9lvtLwZbxkh
r454Fkv+p12HWYMmYKJCk9PRp7+gVIA07Wd9/8ZRF+f8SqUesj//dPNY6p2B
bIeG0LCJghJVkuc6BPp1pWJbrnRmZKho1Rrtc8pNUfjTNs7q1QHurS0ojvPA
Q97oTxeQ7flCQA/I6YSPeBBTdN6NVcLyVRpVna3YIt3TlUXr0W4EWiZelGqA
l7Crltx0iUcbXBjw2ThuKH+EnDkKyC9C2htwjNGXmWYrZXzmpSW0OMHPtSbJ
PRW2mbs+tq/hECUCPdyJCkX27rhSvLJXmqP05vGLz/59anCN4xJR+uVQaord
JFghWqXm7LYEAKHKlHeBkGdc60zC63YtiVUwx0cjQk0316Mc/NNia0HoYwL2
cxQwwjWgttd3BnoADf9m8OHZxv1hvUD5qt5sAE80j0bsPqE2XGIM51fdq9Rp
vV+iB7IPj3iwEcWTThN2vAsR7SYWqNKJCmcVBHkQJsHx+rNT+GhhwmRxU7a3
FUeLQb94VI2ZELnrw76dWoMZqPbw+tk9Czr8IUrj/subRv6SXXQgwJnYwPnc
ArlYPf+Z0l6y//cWXor89N0bj8V+uHnGIAdfKlDFNXJ19zJ0AHBjz1ZBswiY
xxmWGnOBAxsqRRf0dXVsXL4riogyFyrl4yb8BqXOGRs2Vz5QRulLg9jcT56b
sbLE/p0n/aaF+QnRHTIphw6+FimZGvlY1fyPl7gHJ/Hv9rewnR9k6ArZxX4Q
3SqDEtizRRn1FqlHjifPQCu5cKEbCMix9bq7XjjfyMBG7R/1v/pU84H9/1Kp
tFbfq87LFQfeATlZ82c1Hu8JQ8JLFR0vI5bpubAagN+Q7AOUb0g=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3G6w5Ekw3Xhyi9j90n/HkkBUIF40pRbJV6+b2yszhEDBQLsti3lZB91gYjkYEq9sK5WfA/RPyBSvvWKqwkjAXBfhW1U70U5uMOMHu0tv95Kyg7mNZ4Lj60tzLO+HF4NvuQypaSp/lcDpu0eOAIStx1gQvaWHeqidCRqu8FeNJYjnf5Ex+K50lg/UmUfj6yz9Ukb1A5OYxrKQEGU3XRQ0LGPCn9qx1dbvsHi6IX7R2WAhXDKAJh6o03xLTsQvr4bau68XEmEZfAc/l/ihP4u7IVsMz6R2kq5dD6fABB8Tns+I/F7YE2kpkS/laKaebmtCQJ0rRA+p+EH6zYP2WTMDdoVLrD4rO4F609p/hlw1n82RMf2rJw4YBtBX534q9Pwl+MBah6lFjUokjP3XqwXQUkBqJ/3jR2f7wTUPzuG+v0FjCFP7612x5vLO81HeN2xCDfsYMdeKA3LCI9duBqNPDBBSk7hh7zPjr8Kd16ghRfIg4WSG7SbD7Vex/TaQO+V2GQi6ThADH4JErVW2QYJlby/YgIW7/Ia/Abowf7TofGpNmsiwG3mq9axbCzkfdvsATQSN4V1OghGjWTxp3X6Mfef1kU6POzoVrLUbwNKUxRzdBB2UFlhwchVwcFlc6UbnSyjf6tbssUtxOzi/4K9QqeNj+D9L/jMA0a98YtICevGzBKOv4rCZr8SWeRaN54ZiSeWcp3Lenc/gWRjQjGKD3dJ7KxiGmq6EY0BDXso4yfLSSe4IwRwwRa2VnwtbNSolJtlzVVyjuYhSXWphH4w7gyi"
`endif