//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VIs2yX17bhTSspT6RcEQSSxPiZd41vih5xVlRxg8uHVwZDOtXDxLVz7U08f+
bASJKCsJcMvnt39BqT71ptB6VDFL9StSWQUfiu9hRDiBfYF1yrC2LS0TbS/g
wLF/X3yt/TXfKhmODnnjXlJL7C0g3T2XMfm9Dek5VMZz2QI5OXG6+7lwiMkl
BRELWNuasAHvWkHu6Pm5pSdPG4qQAQ4FbT/d7VZ1XQj+oZeR9B4k2lWBUGxL
YQiBrbN+xgEpMWvpTDpchySTwTZL9Q/MDnFKIaoHWN0iW95BAn0H3YO6F2L9
Rgk/Oy9quMfvcg+T4rfipAlS2XT0x5vnTOrbZHgjhQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XPJAqtOdjxLVKEvlZEkjTY+LWrapuvC09d7TKaFoQF8uNgx+ZRC17VIr7mN2
I5sMi16EWEyrR1kczgySyHMj0nE7dXF58WW9MxHxM3leKmMS4sET9no7g0Mi
em4nIWGCIi4M2ZkKmxiQE55RssBgP27Pb6XZYHLNuVAO9n+rYS2F3mBeNrcr
FC9DTjQpI4r8sJhzAyj/LI25fg+zbj5Hy78Ru0Arh8SpmHznLb2DK01u09yQ
lB0nSN4Xm5KoJSYxaCoyl9NUfS/pgu0jGZUGBFbWeyK7vTCG6FkTcnCnqPyF
18IzP6eHNBQHo6ZO+a+CK0CO67OScFqvvVFUvKyA3Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
VHKoANMlmtfjnwhXzd1y/9s//j99sFrZLtm1vlZvSLGWvoqKPf+AffKdcKwX
wXtnf9o2tg8kplaqmiXQsGhScO519FiEjSkLXdexHYTNOKkAlHQ06Z/KvQV1
DDDLdjcMbqSI6oLcHyzQCouyOfZpts5k0Cc1jU21IXvdXhjPndv6veDDTGLs
kF+IC3gwB8nSd4qAFV2YAj0P5oHapYpo6TniPMm1Er1ydyQXHaFTGvMnMQVP
JKU3TIw89YXXU2Vl83ZRpQoUtoR4ug+6pqfTRaFLkhaFZQ3zPh4wocXfshlj
572ASlp96GiqC2X8EkFcBgPjTrQA9Y7JvuJDzQyoVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
HYTb0kppddpLDd8TPUJbHiJ9jk1VDbphu8M7HohI/OtG/SnIDJGPAYrnHCnO
CYTuHPXMYV84BteXWyyTILjLbghhIWxiRNMekEgm0hJ60wR+3RBT45x+tS96
0xvnwi4Su8wKiFYhcizVQHs5p0T21GGmIscExpHRej5/8VI6R5I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
G08HVc36j8tPnyWTTuzE9ULdSusxZqgCMvHu/YwvsmS9fhTWfwJqSewkeHbb
3bxDFuXq2N22rsMRnLEzIkHF3XaAyy07A59K+/QAWd4nqikpoEcgEK+fPMSz
BriYrKurwZBDO3DgnxJsN/YB3r1P8mB31ZsJENMQBc9bjt91IwnvzYG0BY0e
zWmtYUnalqfls/nL2PAGQF6xg6ezJC/VQ7EqwaL222yv18SFEWJ4N0giOrYn
C0NnnWdPadqrynFcoK9Y0jy31BqJMY7c/pXGIRuL0ceiyjxIaeZuPZmEYtdM
bRQpgfB/MNsXRkTgGidSp8oRVh1y8Y5l9RtTOPjeqjME2w+6Lt1mAVTRg0US
yxndlBRFKgVH4+8BZCohNq7vZTZAxC3zjVVHTQie9Sn7ElXRDiY/JT8ZVts4
hB5pKgaasjNnxrbKODBJX3TWL3PrAHOBf3sFq7mrallGv2XyXMK+qEUE4MeG
StxP8fQ+nFeTfXXRzrMQxcOnGDsiIw+q


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KYf5Mg9UBoO/j5JmfE67ZN7i2tGRCYlodBwYybQrf7dQvihyS9CZW1UiHFEJ
SzF02CrBuBygfVaG9B/DVoFHOcSC+qM6dm09+ykTygiY0rDtPZj0/a7ZtUI0
JNOzEFOxA6OSqlS+bzA/wGKknAIbjeiI8LNkictaKO/qLSuc1vI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FSo8O2PDZ2wZ+mAUyT1GzsxPyfVYFA5yYylrNhzYnz80B7Fp5Jj+KFoUCm74
nlKQqeOzmwNmsn7BtkjDpAI2o5Ve9RJQSuU2N2Ij2q2D0nM6ofsBSgSrYZgi
JbVmOcibOkHRFX8Qgwetz2lIcjwljNDmqRrZ1v//tDAU2I6rnxk=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 14160)
`pragma protect data_block
fe6Adzu0WFkeId4AL6Mw8ztjIixjl4nPqZeuv9zS4B2rh1gqXQbY3F4vAuuC
VK2E+mjx9OfhYOcxmROtgFCaoHtcESI4X8XNbg8Fwe+8NeczFQ3gN58is1LT
U3wptRPs9YBHHYDTRTJw4xWOIdr0KempRj5j62vqmvq4OkEpoEeqN3LgatgH
q8cd8RKrRbRphYIgJpTwPWefHQXnSUDZOw1uPQQNwAgnBFnd6PwGvk8Y3H9W
XRUfZEo9uHUo9DEXrAZoZhMUXMzhn95TMWf/LPzufxQqWtHzeKquuO+uiFnv
30vFBQd1cA9bdDvhAHWNeArnLRvsqKOC2iUwCMSvalpSpzpxLBg+PfLBD/1D
7Ev2BUUUloGPFnGh02mvHIUs3wVPT5SulsCdJh1ndbmaT/S2Unspvi+GN9hd
VSy1kGJb5W6g/nTVHoCuaUIPJECf0MGB8VA3OYjRB1IuC37aZUj1liF6nXRK
w0gQbdAan1mstDJp1a7nGkk71JPXmeHXNvprBzgNdobX1vdkOzP1pqetgOv5
K0g91/i3BLlxdIXULu/65H5/BfoJ+Vk/vT61llNIOLsMqMGDpS73E9L6nqED
dhCHkliiZNmEmMB4cIuHuax03WmSrwxmcY6JcvVN9VI6dy5XOtsU4xhvHko0
c8YbYRYAzuvBivKlw73aZfUgTXIx015r3fxScnVoTNrhgbanyrezQPORrb6O
+NPgRl5FbJss3ZY1JtBCSMSrOz9x4YIFHisuJk9sAURBoElYxoTfBJUO23i/
APj7Hdti9mmOXyb8MYnDwcWuLnnuA37JAl8bT98U4G6oQoq2yppe+edWYR9Y
XZRgxGZxj0Mqe88bcAAO8YLbvZKJqMoZzYEbX7xzMHZasyUkxJTCmy/3xBTg
l3E87U8TjgKEKfVesEcU73FFN9PWsZQ6HXlkNDO4mWZNdfeiq/0ckfykGMGg
LKbKokWghOWHIcyjsVL2cHRjtUvF5s39rsqr/aK7Kf1CfYUyqkhcIulk8Bp4
RM7Q4nDkQhmEwnAvjwM4AjtwwrjV3M4I2UTTO3miqwvgMo79ZOtlWkqz5C9U
0fwbzhxi1Dkvd7MsoZDvFhaHCGGbzeTH0bvvq3PVUj2QTBFbh3ptsstx7Ebz
s5KTZVkpF56UtTTXszY5vcI53IHAtQoEO7k8fgqvRLCsPx8BtIVBF9vN2MFy
nRQrlUyEgj8y/mLV6Mt9ZU1yJjOy2jWT4m+QWEsoyBzDj1Mb0PL48lekzJI6
Z6otzGznQ3msWz1qC7gDmNHO3pmifX0kMQS/CfM/jMAY1EOS4E4LY/1TzpNu
2PvM3pU4xE5jz2H3AM7ceXNAHUAIHU5k7AWBwiDtsXghjUr9PSmMxI06DYYF
96mya0OmiLpzIpO9EkiVXB6uOfF97n/82uUqLMceyHnUZZX44ybfpHtM2tXj
KwQWb0vAx4wfs63pYomf2YH5QOE0PhxP3gtOMt3H8yhg7cAAurdDU/+/IGee
Ui0kD1wLzeHfLjkMKBAWc0bqyauf11y9COSx5vSuPkwzxBVgsgz1fSNR8kxn
cp5J6RS8T1h3EtYVGSjnk4gBHZOn53MLTM0C6HEDl9m7IZoba66L4hGRq1qQ
jBjV6j3jN6//N4siCEIXjw05ZdMeaNjswkzmxA75NY2orPfNr/ZqJCADrZcD
Wwm/KJWr+g1gjIyfPlOWL63+Jn2G7Kp2D6p5TMHQaoQWPmR0ATwOh9d59OZ6
WJBtEnU5s2TzvMxrcRh0qa1b7n0uN81+NRhAxx2FGwnamyEqXG9iGgOxlPgk
RKQWycYDpvM75nMalV/YuBLdfYjsSF185KU73UQNy5+b1ELXwgw0OnZ6QvGK
r7IoSSBhDUnhTFGO1VfcrFdJE2woS0sEahAuEIndtt+Jifh9/cn27xpXqNkR
rfL0Ov3dYDYv6u1xPTeTAYpRdBU22h2O0PILpOGdDjGPfZrOpmjE/J8kYTj4
+2/2CqZvSS6oSzvN7sdbhuZxzp1cvBbBvJxRA2sgZ9v9+XxOl7uUjH0B3y2y
lACPj5XfGOzIe0rL+i0a7WaCC+hmQ3uni7GmzKI9bikPfxmAhyKhEfe6yfSr
Gl2X0RVLrSa5VvLxUySXBaFAJSgNMwRB/nCTD4huM6THNOskkBOrzJdFP1xM
DOoHYN8KmX36sNjcdZGM/PSJPmzhco+kNq8Svh1I+awlKPEOSlpZ7FNaPLB1
9HYiSMDOsAyaHYXMmiw+zGRP2aPV1e7nor5C3iVDcVmNXJRKCs++PU9D1b/X
93Oclrhh47qWJOtU3LXLkRQyiyZhHbK75u5Yc6rIArXOxyqanDoxP+5KaQaf
hu5EUQlHneK3zZXzfX/o8485xc84osZVkYBnIpdAWbCVNC7xVarYFYlkIqPz
NdJ2jeUG0NzccWXk78DjLMmKTjzvQ/mbrf7ZGXiiPTp8RyX009wjBi3e23BZ
6bviMG+2FcH94RqUX6GgI+whTz09J/E7Sif+nQhZZP168ErSL/H73OIJ0ZN+
5v7EcBmoDK/jOKlUrm+SV1/2JuDb0XMFnVCOvKfYa8ZiL41hGok8Ak3uZZc2
rj5BHMOejSwDsoCU3qowQNX+dMf9VAnNRGzp/VwC8/Nlm0ubHWWuDsYQdzSF
sEl0q7iUDgniiOQ0+vqd+OA6ZIoj7yCfLljLWLoCSwpT2gXjc0mKLnM4fmgo
ZidrjEzDCaCJs+Kn+gxEajKh9teB+WKM259UJNzqdLorJ3XGkmnZoHtmqUbV
Qw5okgEpbDbtIoCL74AdYU4Pe0z+Sob0lSLsIqDe2ROB7u1/IK9PvOZ9SbO7
OcyK/lMianTeHJ50KWbdmYi1GPZ9DrKJTy5hxX8tq2HMuSiT4Eex8FP4JoTb
KB6CNEzAuma6c37SypQgiFrc6tllEABr/673e00WNMhhMYoGFORjvK66zvV/
WA4+EAIGkMqN6TDMQ88NDJARWxNgFMJstixUtL6HZ/d9L7DlXxANuqmXDdxD
G26ZWX/xgK095Ggc4Dz0Ao0arPmySQWXqZBQdD25U+ivT94O2iUPF25d0i6M
zlVIY/10vh9IbcyBdZ4EeuAsoIHovfJQfk+T9LSk456G5fgHGn6sb2nvI/tX
59mTNQwoTsIRDjPzGkyR529qdjAGLbzWDqsuKHgaYnrW2NkhiP0sE37elGGV
gz1fDWj/I+Ok+k4E/VBiSVb06NWcOxlCIS2By3yqlemGy5sT7bQIeHv7LqI2
q3QcNcKvwQkS09c6UUJe9W8XwhGUhuytM92+tZRWLS0P0mYx4FUSqTivh1+t
a49oxJ/eUPzQ+C1pXlHfo5V20RbibjvGnWZB2dhPIFk0OpfXB961S5kxBGuF
OZY4C27JAFjNiNGREMWlq3e8kMYLuKEOm5eG5nW4I0ZLm9dAC3VgPZidR9Pr
bW4Zr1KOi/2AwhNWc6BpPk5MdESHHyat7OrtQNFeTkF/i8MN7pakqjoiv5h7
8TJg0YPSafZFzhwK9IW2feddHxARo+CibkYKdVkZ+UYCTtPKg4Du11Xt6uzu
0sfuO2LMY0tMs8u40zIlGs9FBoIXwZBxqHLWSoNtuLaDta0jt07L62PK8r2b
y4OFkVueIecOtzKXoZoV3EBkSSgT57xypiYqzaw2FLrzdtVdHJ+6Su+oMdku
1D/AN6JnssxIxlekBoWjAjlAZV/Z2ELb9wBU/+i+bzm4vf2E4RRKNcJqoKMR
mfNTZ4FQ+LcmQ2zoCHyyq+KhjBXa1bvUJX0f5zeO+OjRG2oFfHhahd8OBPJw
gZ3PcJztbbu7U9NiKnVpKkNUKnR/x0NJSrl2XilNYn8QSmS1wjhGLiHGo5Q1
TsxOLh6bpMq+RS800JI80S5+u0630HUrnakXgbpcEknrBYAGrL6V9CsSncvJ
+qUYGt46xWI4HmxG5Fva94L1AJ5oPkAY4kwHG/PGRbUBvhBQpeMwW+7yvPj/
257HVmwdQes7FfUSU/aknjKLSMBPvB5USGtavjZWid4iJ5z3jDaPStZ8i595
r+nzOfaCNVYvO9rd0UR72HRx+1nnuSp63XGF6aACwoqG5yU3RAWToLiX+Irj
LrA2rjuPk4Mnjy6fD34tezjsMCi72fm2nQPOTYfwaLgVy6MMjOYJ1sGncWge
E1hsKWelwZSLB0wks6vGME0sIxZAMfzK1Jsas/gx/Aq87I+TB1G27fctrBZz
2ndt8G+Xpp5a0R4o87m+Hgz9+Aowm7TBzlwrWGHvnjFd9O9aa90vXevh2KBG
zFLKb7oyI+bHyr3iGss5H396kLICq4QVMDaGib/gnm94AUPN9krc1Ju1s4mT
VxaNz9NFXYKduksKl2bRB6/Ya6hPPi2G1z2oteCAaY7prz/yqs2KYhYD3s/j
OBzhl9ePv6EgZ9bqqwzAti/j7GY3gf9MIjcmb9/LAzPRiU1IfKSiKjOfTiGH
+Pl3ALJDTg6mCrWX/kOsnTqzWBy2GIqN0GM4TgAx16DFffAVUD0A40EdMxzH
J2G+CaBa8XDG8T51e4L0XKF/IUYfTgk0wGYgvRxnDbHM5DUC+v9k4BTzGs5b
Cfg0Kg0qvyj6unOD6W2svyt6VZcyK+R3nhhNYbNVL1yzbIaKO2IneLBqq/Jb
A9zp8tHrBPKv+BSUrVRJfkPUZNii5x7o7y9BB4b87fkUnGF9qxWbSXQFvnHD
AifAniHLrYCFmNVuH2PWevz68t8in+krPEmtc24Y8Up0blOv8UVNoQmAg5Ej
ShQa9tjn2awb8jC/7Ba8KuVkvUxK5E7AVpoYvMSlGIe7f1jXIUcP+rCk05yF
MliIkpPrr2cZ78EDe0Yai9mxmkREGQnQyTpCWu5csQ0WgTCz752GoilMcHey
WFXyddyWRk1+CQbhIKhhE0I5CfRlSbqicHndSN6nodYsfBJckJTxPm+Go1Dr
mzYai02n5xAz87zYHPpvbI4q6dFh9729mjDXJvUuQp2UjIEvxtYx0EYS3nGt
B9xOH2dU1oSfB/8wqrRs+l70KR1R2HErVhsH/4O3Sl3icD9MyUvxmcmg7Qls
aOtdxALDTyHG9oJpshs6ERJmdQuvhuHEvgSBCqiMtfL72aRsJygmNdjdfEQz
pXv1SiGwXhNNsGhvN8cZHVhN678PHOcaHPJmAL9GFQ0Enz4U4DwtJ3777Toq
8IsvXUYguTxEyKyk9hP/Enlnt1OCs/g96sWZ5pXDzWOgI09xzKaQYaqx8QBn
gxIQHUOslP1IOuK1zA6lq/FgHZkQbySshKs1hscYOsVDZ8/2CV4FUw85cJGs
QgWyxBEJHqMiyP8SYOpBmNl6GhIXhtmGo4C10yYP5TIuUCqGXe4Dgf72vl4Y
GxzltbkD8dI7StN9VkvIPZsqgP7IVMUFAkqa67ioaMEPjX2/muSi2IT1AB+H
Hi5u/CJE4/r9WkygTpJ/ZFqRMX5ez56qrthVjE99GY6M3S4+0T2j6iHGgqCY
OHiSxfOqfqXyOVmAVoN4ZVee+fuhJmok10I/npGWzuJqiUmjzE9ZKH7LB7/3
4mlGEsiH9B47Xt2Atk/TK6arq8P3H8s7peZMxNy9YzVOYmh6AeI1x1RvXvBK
/luOOKwXGLJYi/02mk5PDRokXOEj3HrifVSNJ0OcbmMS7wZX14Uk9MYOlD4y
idkthPw/A8pcp2hsqzWr96pHVic/5VYmR9zvvN5UyoRdKfZSrWre7dA0lBp2
o7GRwBPjuDlbnuuPxlfMx2GB7TTh84bOt2TioG8k9loZNsjbtmNWISvHjAqK
8AggpMHzJTJmh0J4cfzjOKfXROA87xtDa63CNDdPOxojgT28zNmu2WCzuepi
y9vNHDg/XXUfqgDZEdNF2sZSrhC5VsUy190j3xRrUX62pJvvH9UDMIfrpGgf
IPRQix5NMCTxRZZAvOcHpbZliSDF4qWqeScZHfqky/cKv2OJn+T1VcrGhXV4
LdP76f9Y+DS94QfS13J/eIFylVn4mGdgJbl4pbZw/MAtbh28RDDZbSgEzGlM
FWsxI65KCArlWeVf0oIR0SwddH5t+KhE1lPyJyol3y4gvfftlXCXzt4HanSZ
x6AaKb4h37Vuc4CJFkwmU6TxnFAHsBznijbA2U6BoXN1iS5/7RMtuCym2Ql6
VUC841F3odXwRQR4kxPN8d4KA+hfTMQ7OIks10fQ9Y0O4E/hyCW5Hq8icbRw
s3k+DGFrVYGwFRU3p/Oh37ERuzCG/HipPJlRfqpYtS+NnL79KEAF1yfuPsNs
gTDnfEe5aRBKPrzGDHPZOXFs2prbqm37m5JeZUHvmsHretcKxjNeopNrWUZF
BAyfUWjux8WKqtc4KOECUnwgHlx6kX0j3Fcj9M2FjaWBoXG30f4DmxaGmyJ3
Y9hEzZFYWdVlYze2oinbPe4K7CwuuB18MCw2HZ4poQp23NWDoCBL8AgBj3vi
fRyNptYaV6dvmVR9e8zVIaTwReSMueQC+ItxM50YMQYAnHjTRgsDvRYDKVjY
gqK9JdX+Jh8IyAEhhxw7F9iqF1ehDC5HHmHIgsCD6oCYHPsUhJ9c/JDJ46dG
noOwOdKOQ5H4KT2dYtIQAAm62DY8MmjXU0nVuxOKvqylzWW6rYHr+FrVGbhm
ARAc7fVX3HxbaENzOVVR8zuKm9RRzKhCa5MdnKYJcAiv3/0eAFnD6iOTnyXE
j1zv29Mdt6tu7nzTxkjzG8gQHPwaSoDHBnef7EJzR5q1KJtAdRj1yDBcUTNY
6/kr81e3n6vwCF7kb2/KJLtG+WKcMrF6+ve7PO5UO3ZLRWjSFb67EO8HtiTx
tACBzDtvJw76+tNoknuqw++tgRbsjwLoYRKYoYQvfgxD7u2VyfkmVXNIqONo
YccrAgN7LkRR40XKk7UmPOknaO2hb8LbsXNmlXU9upa7rDQR1dXuDAV14VEE
S2vKCFpbm6QMlY+qP/sXid9R9PULNxrtA2d8emF9bdvvRBpWCHmVLCexLKBW
xaSpwaNNE5AVs05ekpNgZhr/qgz8Zx6ALBWMtf/d+HEwi7MNCJo9nFPKlNRY
xVYC3epuXyMStlchHXh7DCKEvKbHkYUSfUzR5JNku/w8IEuntra4OVZFggN3
GqXbgWpPp/U6tg2YOHf7+f5AwtI7a10f+6S0H/THAAUnNiSoVkUpbIxa0M6o
s/+0PwED2fYGF8aLdX/Wtd8n95g1rcZgS+GOKK7dUyabFTXoSy0itm4F9Y+9
S4m2XM1tQY3Zs1+Q+4LQm/dHk2sF0gl1lZyW+I0Oicf45HZylLSLu5MLyL77
dKKpXbW4MHh5qLPMIkm6Fb4ov71oJ6U3rj8VmtaSXw7HuCAd3jTxT7mKYuyu
n6l3p+5jInKqOWSOzsKWDgUYj9n5oL7hEF/UA8kRpJcP1bgxfCBmK7gvLlWB
sMkTnzbZGz5G8gK7UQA1daMS7fAWI9GEbnq948gt0xUa8//pqamtLa1/Zm3S
SW5ySPKx7mg0U4IV1KRqA5poZ2a95M7SqZBjO3bjm7P18txO6zS181ljv1a+
uXG3RhFzEClLdmqLCWqViyBcvm7aZBqfAvtPKH0JMaZj8hLmF0+IGm5CBCIq
b6KaH2bFD4TglcQw0MT1cj1JZIAxfNKqbLb+V/njoO43olhMJFxb0Du8Bpgc
yDtYAjETZ6bng8N9ilY2Vn8c8WrgAeRdzjiBF+n0/+bTdt5fvjxVdverBwJq
nWTqaIL3+zBBKTFF5UI24c0EnN1dm4KjMzuGSICu7zD7bxs9qFOag4dKLIJy
MPJJH0odxxiNqaeduryoRZrjy2rMc83biNFEIbHXEkX369YVXLaZUrzec6iA
ReG6s/9wEGiPp6GBxj/FtmIRurKO/M/DcV3PVIHuOl9PlnT9Kqpr3P/0X2id
v5jnEzM1Qdu/VpwX5PjnbOPaV2IOT4UJprM4glo7P9t7U2E2E1Tog/xNQfgw
b4ylDau6VoNxI7cImAiZN9bU+8X8SVd6Wa5LwPZk38RzA8Vmql/8uSHn8ogy
mgjKqZwmVTsRPeuDT2Lxwp0QCD+COEoJoi84ZHzufSzegWhQaAa/UrWdb7sX
1jnOQtyz3zn14kOrpq3tW7SEbFnwkcQjTPXxiWfiKeeS9QDK5ocsxmdcEbWI
K3Knj4AqmGFaoL9rZzC9hzMWE/aouzlJK0mwjWvS69TqTRsf9H+eZphcXVzd
pOcbDgoQRC0fsqdNhx2oDlh+vZUTFdbrqySv4HY8Fv6hwHAw61bWOi8U41Ux
etn7iunIejK72dU6ObW1cEsd4kMfw0MCENz2lRzKaWaUGYP2fYgiEkFUO94O
LL/TPwx9w+qmBTmAIE2MGTMtJ4sSQ0WTh19shwqyhYL5p356xTfZihbBdju9
V22ruLZ5XoiA+Edtoq4QSqHTY/nP30kIIGCblU6dSDhhoc9yuD4SnX18vmKK
rlIOMZ3qB88n66PTOfGmmWXCjWEFNuB4IgXosUMQMnBjXGEryLwhE8D5onOj
ynykRdF1sfGh35FGjaTYbuxyOuDHsZaYUTD3IompXWNFdyWoMh1Twn1t0W+P
//r7PRcfz98fK45E4drFwWQO10odNV8J8Q4UPT2Kbt1UA2TvkWkYsac7KyQz
uu2EPmLIKgDlRZel4z69VMO9GzBLfEy9QFqQIz5Kks1ScJx6E8+ztqb+50Wr
7ZbMfPbqXVDKqDq12kaat10nO1gLJb8y0kRMyrCvvL5THDs7DtdYAzv69p7/
xgl1RKwXvZiSuEoDYKkk/MMYhtxnJNNm1TGydUUmnXWda7jayyK07rkyqf2b
zZALqi3ZEGIVCFC+bQV7vnPEaBEGvEgAE19c51Munhxnbv04ho+SSpOC3S2G
8NJgcoY14zBfNY+wmcGPnumXn8dU04kyQyuTxLPwY11OD56NixnHK95rml/I
YOAtkkU3h3JkqL/tBz+jfvnvNY0bpqYSctkDv2iUz7a6EzdRExyygoJJrCfl
khf63ThLh50uZHouI/8Z88TzFFM6s3jHoyyiMqlDCr9k94gtpUDuR+JLq4Lc
+tZyxGkDBvU5YvnnAmw1pLmPQjUuSJsnJ+HtGU5guGO5dMzefHt/8fHjaJol
noY1xRomVNk4hRHtySirEu9tHV+W0+Ye67ycXz3J2iptinLRNPjdu+IW0IDK
e6QIKSiy1IR9Vdg7weThGUGbFGEHrimXkFY8uv2l3CnMRpridTtyBIINIcQ/
CjwPCI6id2tmHhkOMC48RY7StFVNYKqT56AAJJgcA4BXjUwU/Tm07YPrrFHI
6EEBffH1GSKedD1yYAkVnS1gPBOJD1+1ywo1dVXi4EyZMO4PskSXEauaRahb
J2v6CGKuH183hsBT8B+TSRohXmjowmxfXtN0rFAqyL4JsQL3VdCigBQYvtys
wCH6RIqgX1i+GnKznmm3ISBRt1F0XLT7V13toD77rlBr0Y756gvl5n4z2dfD
6716CgQ1cB24h26FHoq6x/rght6e2HFGQRQDT9+liD3WM8r2M/yC25hvMjLI
+NLNk4R6OEM/dwDbEraOE5Owe9jKs0o7C2RjffK4xb8Wh0Udo8PWLJXIjv2g
+BhQHGVFgL5Yk4Frg5kCpeoluxddoEF1F/d8oEYBVbvZASfvqe3PwLc/O1Hi
eDVL7Vk34rRDgCWvvn07eO3U8e4Zaoyuvwwyf+HgEdZ5PsJ+0icevgCmmiuS
CxwrYo+FXDTcAy6JPMhZe729mWdZUn1RxxEUpPTTxP/B8Oxj41NM1o9MR0Kx
7AMaQz6mafm4fhy4vNpvDDFcIJ860wgIGzaAbckTQj0v9ItJc0FL+T2qHg5r
MXmODGoM/Fmi+EFBHhPTFOuZ37ooOVosMMDoD3SMlZxNOJ7g3d7bSBD7Rs4C
ChifSti4EYcUuJ67YkLGldeKr6e5RS1VM1juDP8yXilDJdGnGvDO/WoiU8aq
3qYLDEMHNiFhJXBb4TkPbrMH1v4meVNw9d5CMO1c8cztr+Oqr1TZHQ64xLy1
gz+ccbp5Vd5KTxvXsG1f00hVOSImTKh+MjzmBPUv7mKNf8tRhOMphTOeRb8z
xf+XeXnL2ZvMyhk2GGtnrVvYJwXvG3jT73ZshfhE33W7wsa4WS3drY7N9cTn
I0JJrp8Pm0yEzKN9L2rrL2NNgDOLiesTWY6vO3ZF/gKkkJVAkJV27Ap8a0Ge
GQRN1/xErIJ2TkchXsD+67NRAZ5yr/TSGQt5vsWnpMsuxf0CDAHMo/QWeFdj
Oc1F1srFWjroBkBPvc47v454aRC9POv390dQ4YcXzWyMeYtrOep346MZPiSH
gW4B6cRotbuDWS2zslenIRx4NoJdlYZfuiV9NUuoEtefvJw3U15pj0wg6hnY
NoqygS31+CMouhOPd5+mqv5QJSwZxDqPLGaf7Y45RKzNt7gAfitjnpD+fqe8
ihTJCNLA4EJzwp7hcjitET040xTNpFyGA9DmkW/MHqB98Vi/CYU5JhoC4fF1
TUbzaKu/s5uzDLORgYy/uQWUZJE2HOoh/qPCU1HHIH4OhD3uaGjL7l1AEMSv
wTp4Di4EYFrk0oGpCB6pH9NTCqDIoED5NKufGns/wlmJ1hM50L4IoG8E8WQh
UuruGIAckmWX2WoCvaEk9WvfVyZNbVagc6++VYUTZcTIavz2H5TUS4wjyOkV
cpdDg4nqak05ACC/kzSXh90shJiRjN/liambysLRiBBO6KrzmNr53vLN1RAF
b6jtE0eCQSKw+ChudxCKhjDNzGFWQ3ptvSjT29a8qSWPKwFARPwZjZ3GC/F8
JGxScejlCsAhOo6SMmZVuDhtk0RZnna6Iz2hU+z50Z8PwbUhwfvHc9ygV7WM
WF7XaQ5uV8RwuXt1ZoOinKIiRNezInu46ZWUYS4FJ5Y6nafmzYPBVK44Vzv6
7/JLKbRlkIni7As4ss1+EsSegJYxtAHSjJT54DlN7Ugf+zbiJb1Aegw/NRp2
m2SJh5yrZN9sRbuArLa8pAW0JYc1wKzHCj/mZtLa3VGYQBDFth3cCenTFj2H
ELhaXssH2aB4svF4I2/wSTOUN5QtYiqn1j7SwrFdnQuFmbzPxsg/ndESNRWQ
BWSwmpsTauMC+dmwn593KEDGrrQxUFjALKLoF4eZsPDjZiNDQQX52kSriFT1
0DmtHkb603jWdRKM3Ux4DEtvZ9NYSUKWaRlKigwXbUSXzrSlthvFpOIr/IuU
T7N3wZzWk3vWUNEbZ+3o1adCXxlnucl9rVid/duxvoCniqNUksC1moX0ebJC
9qsAqEdc6bJqp5WFXZqKM8nx7Uq8dc6Kn7Kz2j9hWOF0cleecS9aMqNQwpaH
4fI4DWAhuSNV0o2q1dh+VMCa7kcEK3H89J68lF+CI6B+QALWU2JNPzfeA2QU
86Mm1SHu/s1hMBoA4hwiCeMFQALb0nblobfZ4FVK34SBRuRe9BCTJZ41Psm0
mGc1djKn8A05VpbgwmgupYgEXue667CEIm76ob0lteVE3SUmzVkWuizJZY1m
jqsDHftIlQW05ieV+tE6bLpBPmNGD2nijXwPwUFVqka3yUhc+BdVTx3FkoB7
NU0eIj+EpkEG2D4yR+Jo7bgEIKjM9rgP3Q0uxN5dFFoHXIuh+k8VJTLD8YgR
OkeXFP3eIHN9NhQY2Cqf7qz+/guVVig3NGH325+oU/+mCuH9Hphy1MjPhkn6
B88pMeTVU6+qnYfCu2Q1SikBLSTreyyM/PUFct0AAbeWcSyfoLvlFbIfUnEu
KusNzKcC4aY/IBYhodT+6pezU0MaNZBhR83PnhpzC8zAsew/uu9UqiJK4u+d
kChfOMQ5aIljopWiBYCbXm6UXZiKHXZFv+lm++ufAPykiuaTGOhdLaGftdXD
nCg3P4OaG0jD4f0TFn1SDifPzbHIYY3s1aWtYggEyQV57YWXyCWbJdM+YfvD
pl2ncSwLZGW6baXFiwj28KYRJfDkVyTS+supa+ZNctpyOL9pQ/wsgZKUZHQp
fjOdgYmhpcRRF9mK96mFAbTbzH++YlazcZFyfJIRUNsS9JkaHjb4/HttYvJ7
zXwTRo+4c3WDuWn1iiaWOaRKqsRXR1CWg6w+r5BFm4U0juwH1aLWgEvisPKI
NXUZfHTVJwcTVzpD+ENWm6G9j1WkcMBWWGZ2otVdJ1c+rtGXdHEfoGcgmGY6
FGtcy5wPjEgWh0n35TRy2/s5Ik6sBJ3YgkIAfI/lErfhfHBoc+kFQQIZQl9f
m0TSrNzMp7+MqvFi91EsDnySucKwG5xwJ2vVyZUw9iYX0dKDieqifidraRZU
QQbXIIFTLDblUAB1u8dFRI9AwV/x3eC+uIThsGaVKHocchIvjiz7AlwWPzDt
IcUfNA9WVOfXVUICt+3eX7ySD2wLtZUXC9MVy7rxBVhK72SL4oEemPnuRS1N
8xer7eSKKWH1MrCPbfWE58OOdcEb+VDTywac0q40aQHobzl2SC8T+OgZhXAi
bdQSJjXn9ybQA5AV5ut7CaFZb0BqV3FYRHEWDaQUbZ4NnUDtHW9OOGkStvij
uW58NYc9DKO7M7GXgz/3cYwoWs/UD72+iLFIXk4bB3wi3FE4YCpZ8PvJK3cb
v/rqrx3+2n41XSirlc1l0zH9N8ptiFhklLKm9c93diUkrLkADbGNSqRm+GR6
kH4/f+JR548jDd1obmRGeuI5pIqY3rmLgP9pfihtKsjAKBG5P60SrUNVqt0f
Q4KM50y+8f/iNhZMgv7rQt4FkHAivAmhEWTqvwc15FyCuwy/VLmiPigKhBqT
SRZRxsyxOrVp3qlYNLNOBThJ9HxLDlj9372NcHyRWuuG7kNHWi56CeztfO4G
WZiPaIt2kHkyT/BJHN4oR5Ia053+HydrOZGkq+u+OURqN/vE63Egn96h+TAs
bVkC4wpBhM35HCkh7v0aWjNYrVSpVtOjituVGYoHrYbJbjTSbRVnaSPocefX
uG/mrlTRhgvO+IZaJSmv9P9b17U20NRj5HsAyEeetSMOCXMPjHRRS8v9uQ49
BByh3jk6gax5sd7rFTz2SE/SeFt6s3Nh/mtJthTsF4lS/Z1tb8uoeTdhuDB3
G/N4Xd1Tyy+BEuH2mq9UTEcwYZnnsaasTUd+MPAyrloMgWvqIOa2SZ09hOKX
262UkDb54HPGgAa1F0Wx/ImNcDfW13lKGvAC9ZzN5USK2ocMFTXuYi3udpAb
x0wI+fWvanBgGwt7nWoyoKOwiH5PMs6N4lI0Uzs6keNv8FgARIj/I2byNcO3
zaAzrPYFcHH0BEagy+SrSQjjmHFaUdTJeUSHptJHzdyQvY5bVxzG13EX06Yb
Wasc9O5fkcJcaFACJR/Xj9sNkbOKEZEh9YlTzIgXRjScO6LvFqrZHwu69XJs
YIO4imXf60n74OoS/b8bUp9dISr5QH39uUmtvnXssI4lcFeqKlP8UdVlY9NM
fwYpGS4FmXopdGd7MbzKmf/HLRuLNzQCCORTA1uJD3PsSjUmT9p3J3riG76j
51Y/mQp5fPRRBxZOSNDi2E9nfuYfHqmwMhHYFBiWDq65jgfeI7qVIIUaC11y
NpmXk9pOfpISN+Ypa9q6KVLHrk/dRYDrnEDZFrz6MhHIBjuo6tK4A4a157uC
OAf4cTdH5SUiD89mXA259vrV1rrkfEIfsvPsCQt14qlANIU8nzLclazhb3y9
uPZTcMKguoBbm9dHuNOL0dZrDuEpEvTqJxhqjDRx0FOo5WcNjlMZm5J16kE3
adf1Ehi0OWzB1/WMOUtgh813HZsPls4YkFsAYHRYJgTUlgZhTzhOPsqN1k79
kHdQG8dHgF17qQj8irekl9pfAuwATL1vwIeeaUkIYW588HA+mDT8Gv8UTG/s
0Jt55JQT1tqDGZIES3N27Gr7zsz/QrEiGGpmNrRmzBhpktR9O/J183nTw7c0
Lc40k0Et0PYPoi6NH8OjkhlMOvP0deaFgQaPsov++WZYVo8Iumd+Zm7ixG+Z
V9rYJpzxyS3OR0Znw+YvT0uaIE5tpv3rkGMwIZncge060ifacyLfM8LfWflw
OwJY7CW9w9sK2yfB0ZhBKsde4M7lUGESgCoFgqi1K8dbhbgHPGRvOuB9phs6
cggPfcTs6Y2hNcRrxnNo59tGqLEjJQKLUKMoko6cUFe2GPsiy68sKWw+zjIc
ISEEgjdSbZdvsdv/EgTrcvCDJeSz/fNAsyKQa4uc0qF6yrtKpg4+zhDE+d1c
le0OJ11CvsIJ70kej9z+hhtVxBlyDLJzrHFUsO9mkX4rwVBqqFVacFMLjQRF
jqrleps4Rp7eY7GkjozQhHKy/vGAcnKWhp0yUfKjOaM/7Jr9kV4tS+G0aXJC
Ob/oSM8HixItWnCgSKcGsgLvRlnMWVD26WWtnx85rWNya3SSSLh4M+9jVZWp
SovZ/Akt78Jlhr2HzLl9hbnQAz8fJozzg2AzotAU2LO7mseIgIUKs2JGut5i
uDBZAtQiy+w65GxE1Lv7G8DYwjwyjg6q2m/SIuqIGv6Wr8bk/RPNo1rx5z3z
vwXAMjsTTU5FLWOVmHI6Cey3LxwncUa50pYSUZqZzXObqeWVyKDDPlRsVbK4
Y6m8lDUu2JIecipA0R7VFps0thihvSSqnYved4OFBmQkEoK1NiKWSkmqXG+U
fe0PV51OUOfeRh9iV6qZ6g031H3qrPSYcJ33ePf+KXGDoUCF7XsxmGmgBoPW
ctGcW6JaZ6kVBKGuYMezBhb4hAaXCUtPWX54D8i3FJEJ9M/e/xyhKC3B7/3C
BOK4scypFjiVb9G0WIjVLZFD5bNJxtaSPYgsCJyhIy6zsd/ZQYeQO+2osUXq
Noq2yH1MBaUdK4U/r9cjCECL08Sd1uM/nCd7ZMYhYlJXpTvhMLnphBa3l3dT
yGXAEbf9HCwR9zIv3J5Div7BvLyN6lPNVZNtUNE/IWpExzzAy85A4mHidU3c
ZzrG8k5568BBA7BVCeAPYj/WR2c1q+kIyDOOGOaNEAIi26aycRH8DH5lShRT
K/HPo7nHLa8FMdXnnxLPQ8mbeWlu4xP1NS6ldylaYqe34VZJFg2VCXCVjzlo
u626ArnC9t2A3kKIMDDKHgdkGgXlL2MIoApVYp47Hcp1Qo1JY0BhPzhNVGj/
/xYqo6ShvVO3JR1JrwEOwU1xruGotzD+lXgBSe1HLvbp6Cc2u9SzKlT5WhCF
zxqu2bVWNJKcLWUdVs7thFa0LUhS1qDAlZgmB8kDQIR+5+A2ZwnhJ2I/us4b
LsPuTWy+UcmQRcs/9CTk7cattS+k0yxVbxTyBoThcosAm5eckuzeBirYRobR
VNYko+YkD1fZHivO0xxU8tEvTGSS6srbFE9ShbyT2RP+UQ/6ciWaaweF0TUK
ZNzrTKnRuEJGpOKJhw5lLuXRwXmE8VLIca9xjMUG/LDbEpHl93yiSQ+JCXMY
09VZ2bD4aRwVZL9/JlvQTOWeHWYjcd+Ff3nYMWqSvzzFMbHrSFkeX5qlRmN1
1quOrO/vyR27kNkRCMa3/X81RfrMVm5OfihWnAd50L9RxzrHi4nCvjuMhHLM
NKmJX1humA6bKK456u5J4V90v4CyUcqChq9Mp98SbsANvkDsi396+ISUOnnu
W/92SgTvL9097Rg6Nm8n94vVvJvm/QluxVknlovahykO4ZX/5v/khD+HJOSY
tQlgujD43VWJFEYaFljP39ogQcXb6vWrMoT1v8tnqnJMVKZSbHT4vbI6GRZB
KfZdRs8juGi9BZGVwbM1X9PhqA4FVSgIhXHcADmIzPniV27rBZaboIhwJdaq
aYTWnK86yeH/WlQEOgNPbaCojv6oBab5XJd4+pjglPuXvprASDYYSr8kD/Wy
x5tgmXxAyFZCIdLQQaYIsPFxyO6coUA73nVXAWQs3K6/r++PPwK1xVjzFutR
J8eiEwhrHFTwVkvNxXtU3onFjkpbN6OhCfskpu+X/clDXdMNHyXXKHyVJ8Eg
TAEPNWEdp23c87BbdVOiSZAuwz2DLJtUm2liVE+jQacwrIlG/C0wWUAd6CMS
6Z0y6cWctNR2/OBsEykZW0Ekvdzs4WL7k7TDQBC1bl0Xoqe2F19UBDqOALOH
O0f6HUOafB4ONOW6gARoNBqfNaNZgkMQo9dOQkBbm1Ek92RjJdWbgusN0zC/
MA4p6+bq9U4AZElcB1iKjdX7/RUaxJfLzAaE3BhmxPx6nkQyReCxyPrb3iAf
NafUvtIuJTUjAoFRTtN5dvqphgNfo6x9GaETl+zbAICP6YoKYc8l47igVWWs
07REmrhI0fIq8VERwjZG3Y+X2F71PQ6CIdkzAKmWB4GV5mYPhGhcoK2hbIVh
sW5vAULBHOyh1XhKdcYDqClBOSCatIZZ0c0bBX76HJ0IaDXDbWjo1vdwe387
/DhHlRNqO4vRe6sq8FG24xMl8sEYDUC+OTrJjfycRAEQ1e/ftw2rPeqzEr23
TfqotRXVeeHTrJty0DaM+3nl4el2hW6YTZTaPexjdvrBTvvp8pAGTw8cRnHV
kusgzlrGagGj5abIZ88ynBftmxw95U/66fjfHUealQX0h8QD/mxAXAvBpH57
nadQCsr09RzwNhx185LJim2oRPXdfYyyiCgPOgTfnZ0zhgcYYpssW2mAmmIY
2sRDrmxlUl8Af7pedKRuLFhDT134OMgGUWB7COj4FgsqNmqCB+LARCDGTMSN
23yl/VqUiZU9hc7hBjbkpgrGNSKoJVX2S0Y0zjqgdYmRZ4ZV7Q3feo5LWzEm
HTO1aBVGYxbPi+jO4YXv1YNHc8Nk+2nXw+I1Bk4lZJ27JgLMutGGzfHGxpT2
lfF76ATaIJp/jWWCqc4e/hjmtJo/Y5hRkjugmwP+ryi/NsaL9Mk97OGhgLNx
P3zjVVpZwjlSDypgZEGTVTB+mP1kSvbBVkszxGYz8bw0Gi9won97RomnhLxT
g1PlTlzTq1LTyIQv9Abi3Cnt7RmEYitaOnOPAxst7ZTIK7RsqRmWrT28+0na
NYBP9yVLnUBhQw/yR8n8bDAzOoELnyZtAucpQnpxAIt/vvI4u9lzkqNk7bte
77o+0gNo6bs2En3EoY8mCw5EyOLZ6SKayq8e7i0SBsXvG+8oMgbwof6DAbpg
vQexyJ+ujcjl/FcMhpXkz67g4qkCrpnYa9P6c2b14bTvnFv9OQWF0R3OzOX1
dQ9E44kkXOLO4cGL2msaVnZdCCSZbcKTUMW+8QnQNNJs5972chaz9Q4wKo/E
K362s9euDEwRcOom/dPzpuqTqXk9u/kayuFiuGlrYqtlnXVsZm+4QrcWrH6c
TwMKtvLt0B64xbYD4lP3pcu8Mw073i9tLxH/QmxES+IHWi0SOVyxLw3YImbH
QJ8z+pn0O52kFtNsBWcPesZF1MA5yZpac9A2h38cU+CmDdW+jCaM/GitQe+p
Cz3Pzw+QjOi8h9IbVu29LNK4SYiOxrLP2kkq0uRMQBanNO9rPxfNIlh0kS7P
wQN3RnX8sprMF6O691E+552tmI5fXUT8AUROHeaAmN7C5PAi8MkXG1HEOtmA
X1El5x1scFIJC9lfQJpGCTLGvJwDfRZd09LXkfmTzjxwNv45+OeyLrnQSlsE
yoKch+MuDKQkrFY6udS1020xfc3qwcqVwgFI1P1UysL/cp0QXjWmzjobpC93
/t0bSLUzbkzO5W/BKMQBPskl79giH0r2zxXHNAG6yh0or9KXsqMIewittSAn
YyTsZ9he85AkgtHFBRKvVl3jQkSpNx2hid1NB//1rbAsLAsz7yMztXeBHLqH
e7J0HMhAKzAdSNmzxeo9g3NnNWUT3SM26/d+CJQajy2JMBVxDxu+/9c5GUZb
aX8tpmKTSO4/oWjRIUvQlwULAhfR5KIYzkkQjvZklviFJqxZPeZCXvQobxUs
8CndLdxKM8k5ofxImK3YKx4mEelJSn82ONxjmvx1VF4MXAx6G+EdFjGBFN6q
IkHtrw8/pMBkv7fX3UzvtaFzF07+lVjN+vYDCs5JcbkoONrcFnT4+W/GkfPH
93lfn022sxswl34CvzR+yN9qHDy3dPE1568eKelH503StZg2utPM4BZRTR6H
Y5grqi+MDvOPNuGS/Xf/yHazHueBRD8r3rJp+fvXzm0G2YjSYeSpfRwv/HXT
eO00GtJ+zkBZnUzcuw2/nIU410qw47PhWtSX0nHUIglshlG5+iSCpNfG6V7k
Aknj8aLycgPHVXtwzKZVeAzRmV06++yNKU1FKKlzlmHw8C/EyXtD49xDlMSi
Kr5/DQciIduksLjQKx82dFA+765dMUupe2byT0HoTYpTUY6rvJNbFHU3Zg1O
pQ0YGtuGIBww7TWJ+hqBG+JTz8WzO4VPkHydcTbS10rwlMreEo4Yh/OuClm3
Eq9w4l+TJ5K/5FpT3EBVVFeLUd2cKWHcb+wEzLfimfOt1K63g7xp4MThhm8v
f3tYiqolRZWWpVqCwGHWPVGUwlNuJC7ksyld2r4TWWq7jfL7l9Z0NR6PlLe3
1HVuqnXwJtY+BCb+4exqs7oDGOWz1bC28Rqtwf4QYsJE4PhPp4dAF36YM8ca
z4BSrRZrQ/dYba4gATeSlbgmDwFPuqt2y62byZOxwYwqWGEAC67mh/sDP3rw
nTC7VssiapuM9DngeA4sHofFCDuzRAuJ11IDqZFeDj3nnD4HJQj+aPx3fFE0
WxVVOIo4IlWK51KBj09z1U+U6oJaQJfHDO00gs3OasCJ/GbfknvIQiuTBpVY
ypzp/+zQr5WObN4QLDLd32JPgFPxjUvyCHKiNKvz97YAoPE9nivqzoVEdHoR
tN5DniXfMts94VgkAi6F2rsnM9K0Yw+Q+c58Ww7U27JxF5/TknkVHbAAbmqW
+yBbvnB4MFTijGeMz+dTCRcW8fC6m2V0wJrAnEr1f8TB3dPCJ2c9fZoVeZsi
nCpbYSx0Hg6d+VYcd+xQkHx6nA8uI9IDY+Kj/f9Z

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG0YV2cgZqo3+6rZ38TiQaXdO4dTThwzePrkRU0R4Uapy3fPvhPAJ1QmZkBdxMSC7UTNSnR6wFSNqvBsSsRp1RbEDXWEAlAs/UzCXNLaIt0MksG/YnwaZJq3jbxMjKgbm1f6/poWBCZOQCDcpf+hA6FmCFCKkdRW6rdkC/xB8ckWOKMhMOU4f1W9CoH6u5DVoIJPg5qv0IoDF9GW11akAbzk493tVfgFfIM0tV6QW9BfD2zLZ26rHCqQLmIV3d+8YEhEz5XcVK6c5NWdvxREsxJjKAfejxXe0/qMWAmleB7Md8AGL498jRPkw9/+wWko0DIuI2UlQCVDnGqTe4gwJgfZymwm9//qWHcj+kG08ZecLqO+IJCS/34pUW0So0CJkjculeW89h9833BzUH3stAxsu9kAxuFTpdFu97tF5jUZMXpxPiZXcHUdskLhYKLFh39IlOG+HQy4K+ndGjjyU2VbhD/Z9lcDPC0izcKWZQSHxvCCo8jZ5zPrYWT9BcroTrguDpGat4N6PCB4mvL+jpsC+Q2CxMiF5G6l9UwRKrXH5+b1QBS8jP7YC3l808iQxDLoyU0aLGUMle7ZpMVdBC2KxT/2g+ETup7RpisawbRX0w4M5JL0WH4lqzo7oXg9hXsLFgIHXva3nFluPxhMO+7O6cH8CU2YrKwkSrDuyITQKhZvnM0RzjF0vszguoZVla8Fy6SpL/1JDpdJmIUqce8Wy7wN4DCBsJ0iXgJYJcOPU5+cKtPFGuLudDEPKJF3NTRSfHhsCEJSsusrBEw8YRXK"
`endif