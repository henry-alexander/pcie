//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
JGzoWOabKopeDtOTp/brgJYk29xtHhrKpfSxCwdDhWu+DCfhMTHuRa/8AFkt
j+zRKX6XFZdbHtgyaa6/vxzioCq8JqNKLUZYHfIHVDSmTjj9V56H+yTQs6vV
xPloOy6/J2sFi+m014tc3z+KgSfQkSlL/TNJRUPg0nNRBRJKBk82k1Cn516v
GcUfda5efdxHcXaCPB5T0xotR7a71HW/CeamKZ0JdwTVu7kDw2OQzB5A1EPr
yrbRSPHh1lfYQ5l+XoMgF5IIvzUqVizA366aBPXYladddCESBG8yi6TMetMN
rMZ6gKilPABeDmxOuFRVGQIP+b8c523zufzNhEZc0w==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jwh/I8UNNoALKrq9ZNI4DqVlHmVDWXh+mBNTbnW7ugzdK8Kevu3LKiHr+miJ
yfplDFYgN0iWV77fJrV3HoDvsq55Ko0FRBfcE9moB4Xh1/aDqnsSEX5Cd0at
yVCUUoMm6v098zFUocnQB5I3MmZqCSJmGMyv8rNL29Wr6YlFGg5iKd3E746J
KmoV1pyV/MzLpL/O6UtJvlT6kqEsVSpiv29KwBak8vQynu45oOtJ67wz5lV+
HKxJFwxEq3LeGihDqVDHQ6EcO18d2IIbzFTXwJ1qupMe0hdefUegg05+9eaq
r1NMoyVWHJ8H5ECynbaIf6Lnt6CtRUlvTt3H+omIyg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
QS9FSLg2KZgCFjwg3p6dZ9YpRUFasXJuuDefzrBKd556s9s1hYz4mGLmxzqi
U3jCSGQW+FEqlXOvPZpIdwT0w3SMU+FqdCMkbP5ngPcc5M1/aFwcs7T2R6EM
g4b8maZzteUJxPq+dRzm5P44X1TPBsgfAQE79hpngSVOR2Y7UGcFsCAVcPgh
CvblzbWVGEbSwytJp3qbpe/Qr5BNPKtwE9q7Rfa9O7KK0d2vTpOsj4G2yXpX
lWe6Yj70E1J19awrEavzXxzX7R6NjKDZSvUviTPd2z5Lz8NKzIV7Srcxkewt
28WpoTAyNBC022NsJSLTZ4V28FY0lqDTFjtEGSZwBw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L0fKyMCWYgx+Ozkjl5ujRFyMouNc3yuOhdjhvuHgK+XBREFtT+UqVpkgbtel
8tES361Z1/MpT6900NxrWLhw3wPjnyNlEQzT+522tjAjjIpnoE/Y4Zw8ktza
MW7Wagm+6KZ4lDpH6WelsGOuY2267+xEddAHYFRNemoSqdcasbQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
HpLrlZZPg4UxdAZCVd3AfTDA2Qp5z7OgGEGN3LSw3j7ZyOxAPnP56v4ow1wx
D2rQq1zSE9Uf2I8YW53/Yf4WbVpeg2x3/ufZmhxdoqWrVMyCGtBTd9nKq07C
SoSLgnchpIgHcvcB1AT/VQnVJcrACNFJ890DpKiLXrm83XjI59RK4HpFPOoV
MQlbDsFFZOiJ/8nO6mJLViDhDa8Fcjwiz/m4fsjlTl/Q29gDHXZj94NR6rhv
Ue81MlZqJSYpz3bVT0d4nLhJQYZjYgTXxviMG0pNIk36QRrJGBBuBxNUh1wo
S4ARsfpp+Ui7BdFsfSJKt8sMQbi6yYdNc0VGigze/raUPEK/4J2mVf7IIIZO
M7rffu2D+X+SiQ3ub+yNTccsNLXSwBZpZFMIeLIRr7GHW5HUTerC4E7Mt2WK
Ew8JjE2Mlr+BHcdJrBh1uo7eXPMIA5KoShfclmmbc4XiE9pTxII8z+zmYPeH
x9KaOXHAaQnjX2+gBoMlgPC7UV11NgE9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CNdlh1KWbNBQMRyygDTbiv0tvT2MK9m62AAVKUo/jRCugThkwTTasrCD7Cds
z+l1+Ue5N36JFAbGRpJVLmoDDh6iabw/YUbXds4JiAJ5cHdlBCjOPtI1yKIy
UbZGvelY5Uo+d5XvA2+pgUcXtyod8c1QhdAGoFlGBWNNgcBoNPM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QHAq04BwxOzanZeLbXExtYmUpkkG6sv8J9l9WRZNPilyekltIN5/azjRRQtO
6qhTGTPNp62KcqZ6TTqHvrVLLLR7E84/ev87JHdRcmdAdjU2FefYRy9uK6v+
etOyPA73ZOv5hj+b+VeWHc1eOQqG6QiTbMxPthfcV5nHktD5hno=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2064)
`pragma protect data_block
Yap1cuMwNcjttS9YeTb54FAkxf0EzHdPMDj4UaoZNtdkWStb/dTWo1+JW3jU
XaBVaREhGm9HgfeW0j2fiUBcSdBLTptr9HB2UyKzFA31F4QwT1SSPAkQ2G9V
WKlzmWJOhXcixDrkEvhTQtwbacZOKD9Kan57pF8iRAxjJZmjLggBJWYzO5l3
YEK1GbPWbCBMM/82Id4i5l9lDoIWp1yMCbh7GyycfjurK9CRsyZ4gcMvL0I1
uALIs+CF37P01hd3Ow8rVYK2OL2kRfzYt6b3JM1jkzy6DdtP9vxAYIDUt7L+
qhkzUBiYLnUwrsUz33WeBiRRsOnRlYQBtNdTSDGx26LVQWQ+k7hgMuF+dAxe
UlfMNqx1iqPgS7nY/mRkzMER0cZFEglsWUYpwrBXTnisfJ5dJptBLR1K7bYy
ddn2W3PvLlR0piTUryFhzlWdKXEjH8/llszkFRriMrTp17YSGI9kcli7z7bB
9d+DBiqvsfuCKb5ld+RixhSAibcaqBpA1WUoYcRZMkAX7YAi3qAMbRAr4Iwd
miWK4Yr3bsZ//TUKHofwTdSGhO7l6eIOOrQJgSscZ7HqhtXDIV6FSyUAoWm4
e/QS2HTwz+hDmzGjbHjVSxO2YBEZORC0/RHlIOYjz6CLLq7IWK40MFLGEkdH
WT2VpF19hz6gp44Y4McPtDNt+bCfnaX8MXFZmrMEAjJPE1rx0vRv7JOzQn1H
Twg+50eAisupsjePb1JGIYpXr3vdrsMwgCcbIptjx6ubQWpVqcogbD/OpXxE
PCmNe0eaRlUIjUevmZ/N+wcH43V4STnIl/VSj6sDE/qWXMmK0QnCjn83/TI9
NPIAxoI4/gqrKAQw8npUL2A7J+wmiUZ0Ki5JW8b9Gizw0RSpqAlVSRd9pgqu
y/k9qHFTvSp/0z+bM4EPvPOiwW/7dxTgtnSaw9ry6aIAfWZc5hBlRXOKiKwb
iFoTuEdtHwdufIsz3KKgt5ft8R3ZOngSL12tZiOHJInw/IvQ50kkSRX7d6oX
NFO/AHuHe+zUI08sVdzOFDM6KWm9XDbfN32zuqxu9GvuJcJndo0aYKXxBRiw
VLFuxEplzngKaDCnmTJDX0NTe68JDWmu2iUnjLdO7A99PKufS0vFa1MSmTs+
MRKMpJMYJKSa8JgYVQO3mMJDEgTzNodpByAd8V4xvKQJGblfrWE1UQ2SFXiU
D6GKPHIBxlLrsQd92vyyTr3BIPgMPD2ZzDOXG42TEPwNyoZp0cUjAnWUZbXf
r3vf5rfmm+Qmsnm8Kw2q2dsRlnjxxeTPCAP+p2BIFwYc1BGAJye4vcKDc2Hh
SXYsa48aS2SyEzgAflXwWH3agHl01uyslmVUIHj6BcMucoyfai/I1Qc4ayib
8aKTu4MBoAPp/D/OcoDZG6eKkgjPQhUh6s+4sr5dPfTtLZD/KxP7UBOwhpNL
0Cko1sZnJtF5uDQh+xUQG9hE9lPK7OVm4LNx9bnNJezeTZpAwu7DSMXjfOHl
w/FYyBENjC9DrNVSiROd1pCPdXjDqzvvPPOIXgZQYhJ/dmR3GMnEuf5sIgal
/tBICED68hy9CnHowxgYiBxXulPvstlLm9Ccy0sA9+6w879G4jTCgOBRjK4j
73asVQvQrHk18xAYBYs8cXedhsLUSiVEd93kPKUZA/IASfwgVBs5N2jMS2iw
xUU7krJqee7ZIN4GqFJkpKF7FEOpCpo93a+5EaB23sB+/YMLokuqvucx0keY
hoyPQGiNbE+bSaEB173sOLCzoXISRbIKUvrbbERidORi7O6ONxYHRxE+vzUu
RaYR/IuKUbk1pOhySXFo0mpKL9oAkpUTrlYeUGmat0VxnnuRmlHfreTHIoIw
dtkLlIjjP5PWJzHvC9kaUNIIIzZwtrkLQ+4PVbE7mU6FnMwokBrOsMN9f8If
9Aivy5HH7F0q8vTsnhoZBUzTBacMht7UCc+Ny9eKbJd0SyF656LstThe1FEm
pXH080TeKM20LN2W/c5gx7NLRy+sy73Z++v0d48NmFwNykLGH7CXgJezIrD0
c2jOPSBl04QPu8xMwsvLY3oFyeVlaKog0KN/6YTVc7YgDXYQ+tfZJ4RXf2hN
U/eBejMdFj/sC9Xxa43TZKFB5e505T+CgIGnsjem2VBKVsatu/dgWlTmJc4u
h4JiEFDYEqzmlsJ/KpfKSEfwclt/EGpnfgEc03A/cGyzStjhD98BrZTDF9Sk
t+RKf4FzL5kV4Lfv1K5naL764h+YOPTNcewykgEhEuVtJEAdP1Bosa3YBIfj
c2VxxaFt/qPnF13r0CkupCqqF7WD0zqcpRHAHA+hcQoT1KphF/iNsot5YMbu
9TCNlBFbPw95qrW61mZDOcG+LENQ0uoWvvizjkYcftpn6kHSG6CQe4aiN6jg
/XB5o4CTya0A79WYrwe+L28uuECduRq2zDR/ON04yGJzbrA+qDQ/VYDHVMJn
SL7BJKkuaS/hxi3GbJBjx9uUKXZlFRV+LQVGau5xsriXCg7k8Da19pSm8ZJy
OZWc+6hbZiZOk/5DTk0FWX4FxUTeS3C/3Sf0MWzNSoYpSMypS+YC2kCQDhww
an7CbAYsjiGKDVWFlXuLnDcyghyCa0qy47djyn4AaGhDXwHPky+Ufr6+JwmW
WXzRzfwg6Ktjv410eq7gWfsKh2ImfWsHYa08gB9WJJTgbQw53aUpjPYmcbUh
o0gHXmkWoLJd5Z9Wm8B1icQZue7zKkWNkZIedSssNzopQM+tdPZl

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+lT5m4intNXZ5yGbdfZgo8UZH1mJQzlgNnmaHYOl1qijn8xoT4XogsUwElRfmKdbxK1LESp/9ftFuS05PuTPJhwutfRuvNXVmvwAsxbVB+zWSqEorHCG7nfjhZp7HXzzc+JN0K3qRuG01LXETKXRU+WevnJFQfq+eiHDbD9xLvwknBP26O1YHx8sCBM8sTXS7n5anhoC65BXElJAA0KK6RMlQ24Hd17UyUD8fBRcOHpXEvo/FYdurHEeSJd5kbZb/WBcSZDZXHlhBNcN1oWSIOTiEgwGj69exFKl6So9u0cAA5skNjG/jDKF+rkEh1te/Ku1s9FMrWhs2qZjdEoZPNXODY9cO+AsXJtpk6PHPDWj8T/hyKBJ3PATJQZd+8PoU4pQCnwXeHfAIMrP9/Ud5F5W4QLlMNJwAA2WvzOTAhLrQEws6ss1bk80vqzxCm3Irz95Ct8WRW93XCGKJea8lkkCYcDra0/bFmmK1kqEu2e0UmTAp4fHGdz087Pj5fAkkX3AQADgOf8c3m9m695BzMJqZ7/4pj+LBQxNMvgJyBUX3iOZ/Y9sU/7ALQKW2UwvGBYmlBFbh8VJE7I/W26wizlb73e2HvkAhm8E6jCBX0n7NKjMMlxRFC1eNio5Ifdhl16MAOe5BGlQCJYt4RJfpFB/EVAlTIsC/cZ1Qhjv+FsaYnOrYObpBqUpwHZXv3fzFbPDdQJirLekAFNF833jIK+ety5RhtZyfC/A1cc/zX502QTT9vvEQ0dgzJTqNH0RBhczq8z7qva1wF7YenFKoi/"
`endif