// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
paKqzH4hbORdaXSICokLR7okk8a3o2GsEvnRG3Nije3RaOGDwL09uvrZzfqu
KCaMCxfUPcDqJI3U7txtzNiO7A2NRIt1MiP9F4ARali/C+Vpt8GVcVsQMgnV
UUElE8aaiKa8Qj+fYwVT97ZCTyG0ew7Kr9Hp9E+JYw3aUFUGQ3Eq9uhkQzMN
uLFsg0H1xUgJeyhnLB7Rt2RuRtm8napwsj9sBt9BwRW7E37VOAU2xJ1IiTLK
0Ez6rek9AitMgtPJ8zx2FC0LS+OzbXBi53oh4wCBYO0xgfRsIGNzJ/uRJcKF
DfQU2MqJAtrGTu6XLT4b2dB0SKLuMfUcssDjJNuqRQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gxdyI1C/SiFVuOD/H8F2iDUOSaRIyJcCtUUTGOQCvQcC0fPnCVDNCCYfV7S3
gY/EngE7kaAD7qt7/tM8kXtGnboPGtmnGrj6QXiVf6psDm418TjfB54YWmgn
fD2hHt/3YYbsNYovYkuN7bpuLQTsHb6DH1Cg24LEVE6VwNabcWh7X8Lc8gc6
L90dwWjLzs8c6dfzJo6hVG+EBJvv6cPuAx2IiyYU/KCVEK853shuxCZX+2p8
/ZYRdgGOIAQL058hpOyC3yXfZS86OIEpFxlqLpr68+4HK/M/2elEpGM+FSuE
8xqD2EMMgN+bsKxOklC1jC7cwGowL/6v5dHxEXGQaQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Jj/xWKq1kAGFam4gDjpLjT6bE0LaZmZyY3sON49LJTn84/EoL5Jl/q3vDGt/
5hf1R2ZXKoBCAD2aiDDIr9V3DKigLomR6MMCaCH2qEe8N3Rwc0pnw8RR+2/r
CrrW5mXBsnavqIRgatdBdaa6SRkSY0XbmZeNBWfCn+7PLb0Yafzz+GkB5yiC
2asR9Mr+mf4GGvbqXd6m2zBY6DHX5x1AcO4luJbX1wyBxkU26Nv4oAat8V6I
hslcPTLNrkbNeVJRGpO49V4l0C0TYtupU0xga3pw7rTr+sNawiK+hTOu+036
GqdM6qFz7Lu04fjj89QJcCjtfEF6ygk/Z9UtSPD/9w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
GZ9mTMuVQzfjeN7ViSm7JWqa5vVhvhvOfmxPlR/bPp7UCYohwLvzQL7foXvr
+zo/nyYWkfeWWyHr+KWPkJDWUHvxkae+2YjT/9JriuFhIdBzCaB5ZkCrVJZw
yXBNLbehCyYjuUwadZEeodgyt3XW+4BU6WJ3jO6rpQGp0EmFUMA=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
r4QkGSOyNOnn9mYdWvQye9xDvtZbEagHK0ZocfEHk5ZMwv9xTIoZ426LJrgf
OvgCBHzaq1TL15iLLPhwIK2Tg06A4LleKhE8ZQoxoFTrj7FhCDY7xuMvE6DK
6LHBsqZ6QJFkHEEw47lqs4y3cTz0aA02TOdf0M2dVxZklA7C4fcY2UykK2hd
vnFvlE3AcZLCzSEA46e0LSp/8U+QqGQhBkX/sXEUHSGWlA2SeGF/HQnMhB+V
ZGzQBYXwLmBUq+HAjn2WGOCRD+A4AlYtHUSHNH4tJapBZLcVcPg5a4saX9Rz
nA7d3mJOusA4g8peuNOzG60lrb4WDM5Xf4Bn7FJ1WUp8TxCG2+0Y5ImKCgSl
khx/PFiHvafkwN7EuerJnjpcDbgLUYp7Sy7ATYs4tDnI4qtqZ8/PPcFUH4zy
v0zCXgdrg5ebSyXt3H4B9SSHwny4uf9Pul3hd8/s4K6RtQH6yiXSSJek7FZk
ioP71BPupQlHKbPiscYlHctmReuX8oal


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qyrbTWZqFMUGeGdQAl1M6xrA7EMCr2AWz+IskulIeTlc3d3Mkr3y2Prj1pcI
CqSpEjmzMYOQo7OdlPTJVlAaPd59NuBHGK+rV0HkNatlAj0WZScvCMwC/Ia7
UPe1/x4NZsGOh37MS5DCIZhR7DcteiSrmFUvCSEi/gBQYKgeAi0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qMh+thCB4CZVkx4/NOCIwjsv8t2c7DCqKZ/xBweRfXX5v0mKo5DAqo/zvygY
u3M74FuABrTEZ86M5uYtSx901WLboevJH7aOZgHolnFctbkUwr3lnmzznhi5
XEEQ+XHBQhcEp6lLP03J1TOCsVBH0to4JNY6Dtl62+zuhJBmdkM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8288)
`pragma protect data_block
dD4giXseSsbuIWAuar3NkHkAuM3/tTaeAEggyWDsNjFBDcHBcNfWb+5XAYx3
Q4IKirZ7KG1L/8ZRdvSItvmGH8qSRa+Wm/6r+0J8NaFzIAzZ6/bEUzgnvrwn
VJ5gSIIaYmPQB9xJBURBbjUFMnRvPRzwF8SQMrE04jD8uTjmqzL41DIgpW5J
VdMqtgxYmrtjsVTbaTUQXeMMkSbbtN5mYNUa/YIKysfkFKaTh3axpB7/zH2B
W3AkxoSaqOUuB1gDaoRfIwemarKNBzwtMuALc7nww7O/Y/BYbExRuld3R0jq
QiJrnpLi881zzUbTzzeNmoeQrob8UcRkGxJRgLVNC7ULSfcdznP7dL+NbWM9
Bv05aIeHL1Bn42WSnLnWYhCRHHFNo92dLs0fC4v6Mo/2ZGdFoF12bgRLzZ4W
eMo4HKHiw3/HdVGh9wf4eOuEld2xEFwrVBAK8efvAr5jDETm5kXv5DKFq2XF
VPNMSPpRN67VuD7h0/Mu0cWGv5H9nKxG5clXacwUDv8WDuZ2U2Wv+TWipn4j
3Z5I1ywZBsM8yPmDPdmYb4Lp3dxiQ0xdWOlwQXmUYbw01Yb/yzXn9YsTlnYr
csUX0tJ8so/wuImz2k6oklCBPJzFhfdYOjwZNqBrbssheZiAOnPb218euOBV
x6UbBK9iVG2tqeFk0Z0MwRblEb3yx7IKikNx2nXulAaTcwlGbBFGk5v55hMk
gtTxOT+nulmlB3mxq9DAP/0I2yZTEyoOW2UB1VduE8Kh9Ud3yHkIpAGaErl8
Lie5LOKxRvzRgA/QJxyewqqoLFLFQQCVk6pV20UtvlFueVlVLdfxkMzmH2cx
97X5CxzbEfdJ/sWy5alXQfOaY6gZTlo8fX3xOqp5JrwDpawje1+ONDCSmjWW
DVENUn0I2O6kb4d+aslWxVuXJp3iCEnvUj2SKRR8USyFnZuP6j/j0ghFg7ot
4UwOSruMeuSz2vWDPorPWMbGEjlgrNU5TsFu8YZowLAFMa/TydrCgTisfbGP
I2Wxh327s4W166JMSuP4j8ZdYL2o8z7gfc7G/Ois6cJvgmqabZbKEBgiEMVi
cgozN3C5r/VPvd/cyh/S0DjfcT//bVTrPsxuD6HBsBanGQmEP++mJsye1x8Y
rzSDJhwuQD+DP/MROP4AV7pwROeQxvRNJRvCQeoe7JOaf1S5iSRcgbA8Hptd
4NvIari7h94wwCp4J9wSRcMl9A2DeJmSeKIxZ0fUGM/UN8OoC/TKxUODptoC
AJcUOpZPrTrgFLoUnJbDHkIjGF+9RSFoHPExSP7vYcdWsK0+QGXZ3W7dR89H
ugJqWcsCw1xtrrgMLQPukmYsI9f8NQ+wneUzlIV+8k5Q93Bjs5bTafXTART7
X3USPXvaeAmOmrKoimMTvLy9WO4pqUsj1TU7j1iAY7HqurA4r/pTXGXPUB/3
zd4MCoWvduppI9TQpAWd9Ls6u+C2vK1//N0VenRUbJWu85ULyXMptSyov0UR
yAFwmHHxeU2/mQssFfQRloX7SlUB7WkrKNWsKb5lhoSEa5KmJmztdA1jf82d
rIXYbrkWwntzGN9GkwXF3rzOrHnGg0WHXprYbbDSlkxZ333VTy+0OU3nzxja
LtIJh7+d6VQPxGqDm28SAGSCrTCxJGvRjHA2Inl/lTyaD8K4aWc5YLh2VlG4
evK1Rp23LjW0726RccZUajcZsipjFgxlDC1q0JnKEZ+fSXnTDm8FhLNNKGkY
u/V2RDh6tVfXr/j5mk89Q3HjNqRCETsUrzq7pdNbBSo6+hwpqm6TCccdpo7T
WX2P6DF2u5HD2JL9I7vLQQWivwsr/e4qe3tnvXm8fF2eODCn2Spai1y2UwiC
ojR5wQGYxGOQWC0gK3e58PRW8AO0eAApUKJGEOAzqYSeAX8IYPl1fcPv1nRm
l3OUsBTVShrfLGF1dsYcR3h3j23QtdcWrob3OBPBtG8/EwhtrqRa/lSTdsMP
WWAVYMXzb6aT+6rZQkRUXcJMrzALSA1FwJyGsYNgdJfO3DQQ9avr9+ZJeVpK
bsKjJ1P9T7Y1E39uA9uK4Im/ZZrS4nkSqM8Vf2HjebH+/4cR+jjL+Vz/rw9g
wDfOH5xqi/GO/Z5FbvrVqfE7+ZwTblmThyDSbbvg2Yl9LERpqyk5oKhoGr/A
fFFs6qDlgoj1nVQDaLknMOkgxEbWO+k4hUWKRHbpPKcfPr3WA6rjkr4oYLUB
UMnwyR08rdPb7GIi7ugtuUd4phMzweLuDPSp7PubiilmMH55RWkLbN0LX6RD
wMjaFp3DE4x2VYszrooiT283jrSra5nC61UGLvA15Jlv4BPf7f5YDkDNyLoZ
Kr9pq29x2CfGWP6H5J5LB0g5qdqAws/ctP4CnzozVei6ysVpEspRPf901NNZ
vFTpWJLx/BF7kuqNUZbJO4TZFqvR7UBhj0FyXXdYOq1TiUIZ3XSeB/Foj9xX
Zo4s0tIzbEtvnHxYjMleYihgwQVKGFwQc5ZuV6OsybACb6ZPAIesx0KTuKHk
ULnx4tLNG88t9+0jTYCFyGaKujlGbnaugmFZgMWbW2lG/kkkz/n73HEB7F2r
3FO/8jYiBs9JOFZ3V44aJ34USakl9huPtvzhrUwD7alGw9/QxRBgqVQno1SI
dJLB+ITLL87DE5gcBa2KQeSrcfSozbP8pDzufy6QHOX1OatAhOyZ+TcQ75St
9pJYsj6KoBwH32lC6JzBDDtAtT2S8XApoBZ2MbgL+Uu3qucwNA6E6J3uACu6
WcsimKe1TKttc1QJdF/J5biQBSua2rVjJVInKdjYtyxTVpqOaA+cEh2MJI/A
2phPf4zIvWvTX3wlRrFFqDaNt+u80QTIFr31wPqM99AvkJK2ggatHaRMiXYB
8SPLbOK7JrbdC8RVgt/DxtuQTfGbKxNumtT1ZqXb0VVMuVJI8v8JbgVfk0w3
0V1go6vyIqCP5kz06ztoMBagLQxBDNVHijlkkXfQxbRmTB9WoJ1EtSCRuDBc
G9TgWdtZybtcNiVP/Zmy0NHwSknO7tCsYv8dPtdq36wCCXhJQn3Qjdwvo28m
GTmFc2X9KJUXbDsIDDVMHTTZ9wj7WusflBVHIi5CShYc1/+BceN+Gb/UCGRl
bfOVnz7LtwpSwSEbmfA5pnomVx5lnz50ZoNAZrciG2r8z653cfiIw7TfDnb2
HuUclO38vdWRd4E7vn6uYxX8SstYY6Q8E/WpztZ/yFHGIoeyjJmgb9rRg1GX
3SS5vWSNKLv70ovsGkJxKfg5Gbvue0qUclKS+MYe/aHxZfSTlmAUJAh2TF1a
cDLdjXLVO0vjOnAkDTyOVGpYvuv7ely/r2o35V9thYpDNYP97c9C4fwM+6m4
JFGkcDWIFeD9fcXUhDSHmXQR0hAkKXYFhoFe1Wv+xkPRmA7ih1aO4qAFYeTp
yY5sKNY9LNvHz5PNydCpnPt6yVwGlpagpsUr9lLX9G1e9VriKG/Z8a9KQwmi
8T1cz60DUR16hyZ8FrNAwGozVhpPFwo9t9F6H5bpDSu3XdM6OQKHpQBaRXWh
ZJqhYIQah5kIOdmJrR/K7zTHM/tMt7MBMR9TwG8oAjgM0e/Ckap/khjyGZ9x
9VUtRw05jyRsgqPJV9lRobxk694OSeC/NOuKzxLm2T2Z5gXq4XW1SZXUsE/5
7JlATmMVUvzYDR4iguUieB69oG7sdu2wOCC8jkiruQ/T8FapTY6OJCqGIs64
u351TUX1PCKjE2tlXI9cO866fM5MIH1mJESMfwuyMwrGdmtFoz3NP6yaQsYz
63BeUoK+Yr2IsrbyeIAUf24cPL8BSPlc2hg0aiKnpMv1H8IcBVCrQwkOs/K6
rISnYE4Ft4RNUPAZnZkpaGfCYYhQaozX5RUD0a8kDRSFiODhF07KtbAQPQzZ
UUM303O4dzXwW+OepQPkNCQriALhHIA4Lyhkkbk3cm4fjYMH/45vkqdAuieC
2/cC2Kbqkm54EgtRL9vQ8DpvL+dvRcNzqiYvTIo9dNYb1n+Dbt0YmWHyZ4VD
il1WS3et2DH/8D9EnaknWm9ZfEpri+fJKn4TY/QPNCtEvBRMWsTS+BFV0Kvl
YOikKaMwAxMLX/2dSj7QnokoPJXrlmEkHdQKKOYDC1QpkwE0VeJah7lhzIWg
ZpfefhxWCXlEIDD2PTMzC5tVO68R7BrEWXIkxj4Rwbu+BtEe8MiyyCDrqGwb
L3uPkSYTGuH8lqGy2tXGQhNh8iDTSvM309wiZnYU1HK3cZEsi7yBjzSGJd4E
sm6S4/7SqWcAWbH1LGw8nX+1TS9X8pXmpPHiyeImY7GU0Pg8O1lLYN+BTDd5
35LKiPVwDHgtQNllawRzkCfibamTxxgVvRnzfSTNDtry0rjMxKOZU4rKHVVJ
zs1XUJqlhP/6gtKOdkmZ+kvBJJCkKcMesspSfrneTioxWm5RA9zv6D+U/RrI
5UynWvoBzUqMrmlSGgDCi2HoZSZJAAsY+8XlMaMnlfBwtlLZ3zRUk4Cj6oO9
1GbnJYpPOcfXBMIKTpTWeaXsQqhfflLNgsgurnIoXAfb+elVH121AMDQq2Wh
I/697gehhrTEG9wO3k/Ov04/LsN5kxeveo7e6CToBxU83KyINL1EVKUt4t9F
IhEPuH46XEfNFMGfrlGWtZd/3oMbUrKsV7yQ1uvshUOrHM6KkfHEpSMbx6PV
zbIm6hvaC00CqbgIZtywe4kMu2be0YXSaZwjVCPpb2aDlVnl8I+wb2MnGgss
N6ULwru9InzUiZGOd6ELg9hGj80RfaXtr4EjuCshuAXbx7JkYjZt2mEplWQb
dcfylY7y68iH1B7se6BWo6hnBCnzof8wDnW20DVkKlupBcRXhjIBuhEC9NP9
NkaAt/PVPPfCFs+/k/Yz09J2dO8ZO9i7lOtShKB/XRXnvDXuDdYhBYHydXLV
yMQcJaDRay7s9S6GqEaDyMKI4LGFutPJLCc9oL9+c8HMnZc/RNNYDedjmkva
0GcDXUqTxb8bhCNbBtfOPMmjGszTKYEbjZk6wyiucha7z2HN/NBWsJ+4fQeh
EXLsq6eB5Mkb2ReUH7MXps3d7jBZJqRZCNeH7e4wgmspGgeiXOiWT8mw/JiS
N5h4F6sYHtBUPAW1u4Pcpne6vUY1gFWoqpc7UvnqE2OVpZqK1927V7t/d4Uz
pSr8jkhM8XDN7qzg/AS2akEW8Cx2eXWBpMoe/9xsIgAdkMQWfGIxo+5xX4lR
h0VgUhqP1QxGBmo3BrXStIui2RQFgz0Z3AMGrqxwfRN+VjYaAmmdE84cRp1W
vZ+/VFBkR8IfJ1YDiFj8b9mXxvzWTP5dLiTxWWbpbVbzye/FkLHsrYsOApUE
1dETugtTqgKJRJO9aW5x4CvZZ+ulhJfWKc3C/vqKRhu/HLJoOUK9eA7rYzyq
3mOW0owcepPFRUSpErAfrw/89Z7ex9Crz0+cd213RrJ2PweCXrERt/G7td4Z
cddzc3cmViQ4E5pAz3nJTQHhls5Zuh2torfVszac+lm4BKE48dxT9euVdjT+
oiDoBBxVvMCm4oyxObPyVptwGfQ57yRazZyVECvtWskf5eRCV+R/ooOSRyqx
j0IqDKe6GAL5pW+6AOhsH3mjNsO0riwKhxWmTlWbSDFI0dixxVk0Ybro2RGM
xp3WJFLfEZz02w4w6rZVW2TNwvOGj2ePnp0a2LZw7l1+uW+bxvuk/ty8JpZx
UTpJuhxbspQ938M5f/uEdopEFfPRw7+1J9iAzgBaIBouSM6XF5mtjcAOUgiw
41k5b2zTqrSi2lUphL80RbpBKlIVIKsxu7JlP4KnFqGjc8RMZRP037HPSL+z
PYMSW9GaJyHuiQrd2fJocRVUoK65MzkubEEDtlDqaOwqBP0zqCipGmmG8i0X
/J91c4VgrERsYfTX4gQ8gw4zWnM+wOJMrvnQkJFY3aaOaOF4RKlS9Mup0KUa
n7NBj6GFRDuUWZp6KV5sA5HMmdbY79VilCQZwgNWnvd1jO3ItU15gJ7p+GIT
iGtLEuRqWq5doOuOYuMqTWIq0XpI6l9XcQgBrt9/VZ58AX4hNlh2y3pEPysd
sbFLWTQRC7fN/RQbKVm73bJ7IUpembS7phhcx4VYqtxLDCo9Zn1bPQFDAWZQ
9FhZlJ26v/e4K/nYdVV2Y0rdINkDQIBEBUGAz3ZDE280Bg/s6476uFcO6ulo
sR1fNZirn4f24Sh2ICQTfvlb5Nw49ECI678XTJsO0HnppzH8buvLz3FGGL+l
V1WP78hV/ohPCEPtMyNgm27YBUKuIfPSldC333n6h5qT+GTs4NI5SgXbqxNl
+Ikn31XXiW5Ym7ixQ9Ap36625SMOKmaJknH5lmqstvZJ5ZgCZLbcu/0aYgFB
iOYkjBcv8FHnkiyYh4EKi6OYQQv6y++xtNTHlNtYyF14phNdqY9+kU3ehCYZ
pz7Ddqcl99HnVPh7uHyiSHsGYy3slnG2I+aUjRZrRJ99mJweskGQBDaTGUIm
TtAjzGsng6jRBnujs43jZouex2oMSUD1wEpakaprW26ZbR9OIvd+9DG2O8mT
XDLZi1XAXMkrF8OzLCQIGf1dE53KhqAY0yUpRj8F0NZcGQXfvRTcEIy3DGAq
B2kIxcVKIDx4FTEvBHwxe4RYsgis9rQemWjP5VEjlBoxZcZjWZA0P0LqKEv/
h/W447CTFUUDTm7CTAqSIbxWv0Rj1iWBU3hwn9+gN86SIoXBTs8n+Hiv4NAP
rX90JF2rT42rKR4ZIPnkt52R4vIPY5cf4Y2f3ouocitQfv4+qQLB3JAJsM39
PBtsco85aCXkX7GPWk0rzsrLHR6CVaaZDvBGuORgXEVz+VdfIUWku5W4TBHr
P/nwxWiKTD7PChbpSQo6+rIkfQEbGxJKZcvx3OdoCsqm11tMA+Kx643xKbs5
JQ4VwbSjlLeeIsdKYIckYFFUXSODjDRAzC9PsbtHbwzW0cmAHrXqvCzTmk4a
UeR73LFWeG+nye+DDRqt5dd2pzJS7lgrV6dy9wb78CZVsFxj82kUNEjJgWD4
kyMZNs7tJ2uxbHAni1HaeEKlMh/ZVApN02aepk08mUA7Fn+/pqjRJro5+3ts
zu3l42ty0xusPGM0MPgLGOkVm9pw13rmsp7TTtwKuUE2dXMh4BG0/PMlF7Jx
nQ8oNr/11M9qOkfigyUIaksD6elEui0ddvFr4/ZEbphAOJajZdTlQyG3jxwN
5ik1ByAvCmVbbBloR11b2TP4/P4mDXsgqBLanWYv7Tw3Oodf5ruxg/rY9DXz
yp1ci457TknVV9UmYvdbT/wM/WDP6jQ7zU+PDc7NEfOgX+wCMVGijK9LDeoX
RKeFMWKnWZEj96HdCjU9urNNyAGpWRfXQAaTy0ZJU7lObsfCX7QV+eXBMuLE
qVCBOnwjeS/7jdFt2E87r0IeafE0iohRGmYl0m93PBuf3RRR20hH5qMdAK5t
gXChuAL5yFPNL1HoY/bQJSUw4VOZZwsYlnDXOrjxHgzklIvtlRZf9bqZoCzV
IPA435DCMeh7V8a0wUdFKiIBquiyNY5EAD+E7vJGW3W+bRRpYTfREzIgE2cM
9R8MUaoQyxlSKKYEy3qwSH9GHOlDyUW1V6H1k/dk5RDSKt0eNIjKhOLWsnMo
icZOpBVrdCiieqw4hHYrXq15jYdlXXX7kIlqn1XMjJCpKqkWVBpcKtLfypNN
iL83N88H3UodKz8QU2KK5YIkKP9FrCnLKJMsXvHIl9cxlknQaIYAdeXfFWm9
NCzrKzEEID6JuSURCBNlOv7a1CWdz8M/BDoGPuhhxBI062HJgozdfY7lPUcy
HswxXu08H+bEzvNnQ74Y6i7fZIfbXERk7YjEYCQUdvnOLNYaJItsz9G7l6tn
NyS4bNeU2oMQq08wBlK4sh+mLMpMqYfIdLAeVHUOnbbkftcX/B8UwDUyGvwO
VAu8nwqAxiWFogzNYdQuSIwCttg0Y27rALi1kLdJtoL+UY27twBHOwFh/6rk
jdTG5KHsixt4DcDwAyj6ZHLl0dqiEEVPXH/O6Mo3OsynaUsQ7kkdHpzCxn+z
+eb9opI37Sl/ApohHFfAgRFl3+xOGRBQU5Rs7FLjEiG2DCvY75LeIGSx/rsk
rKcA+2vOmSY3430GWpVenICe6mcUfhvEFGaJQU4GZBkAw8woetcaLwzUXUzk
scDeUgt+dxc5osWQYVMwVa1Ffh7a1STZa6ufp3FAumaCP329F7+oBkf/wivU
9Kpmml6FHVRGR6NDQY+LPFKDVNAKvUg+IBW+kMyJNLk83TJ5/dbd4aJrnsCc
nCbqUEmKkvcKETnXJA3qN9fMPiOLAO8OO8aYxZaXYtzXgpQgzo1ctxauTZF4
WWeGbTCmx6iovx3w22H6JQvPh+WHapJXNp1qh66G5N6suofSty9f5emL//AL
sG8TWCm9yoggbxK64KJHA0NfBYXXFm33FcuwzMnFb1MQH9uoe3JkeYDSdJqc
5q4tUh8F/3YFexEIGChsdN10X5VUVjwAvP5I1v8W+YwTuAo82Bh1uS7XtJgM
VqANj6JaxdbTTrHXrU8WnDq0P/s5g+6Z3Wklmj4YU/9jg16uVpX1ZB4z8cR8
CLCBpCiXJFQw4xxiNxT9U4HJh+g4F8MXK21pGeWSCM5pDEtHPzoyNANZO+S+
dTrUa16Er7F00jnsm9xQMov1xODNK3DjhMqey6Qjg5GBEHZPbG0XTSYlHMrZ
xzkqo/d6kFsu4G8KbqRog1AaLQmkprkbnIhbJ4ukPsmcGSjJEP1XkCKEfwoz
X5ls0J6Kd7xfhakN6CJm+JfLC7NQri9fpE5w2wmKS9TaMGz8hDqo18+GSgKh
kaQNiVCk2p+9zwRjpzTdHOIVe/pnsqv9qnTjMQo0mi9wh6F4eQQPnuCohAT3
T8XzcM8E4HO/syKuzYk6/Z8KxMdAp9Xa1PefW5xO4avxBUDp557eXKGcN2hA
tpdmxLsPaIP0OmwIS9WnD/GNA2VBeqDEg5JxuqoQHbBcFYluYeTEoh20nE9x
wiIopnO57f5myyoJjtf6qgGVV1VBsdntyB9Fl4CrpJI7FkcApl4qd0iomNAj
Qf1iIwUm+X7wjqQCglD5g8Cu72ysikez7oAIdBkMaurv/ACsL/V7kNSOH6cN
v66ld53MvxzXEg7Pz4eQTVbPUmjA9xxts1MOJ0x25awPYgZzT6d8R47UYOuh
PHaYC7rIRsDTXi3WEq813Fxqz2i8x+1xYX0mvj+qtlBBQxu3JIz192+RKzsJ
sSCpSwVJvXU/aReMjsZ/9Cf7rR2MVohMFzTO23GF6vxw3ewJdAnon98y1UVd
t7zAHYrmUcKhUWrNNJ2bsGfceca2kBKZqNW3H2Cj9I96Lgy+32kfVSBtDWa6
EqvNoHw+HRWzx+8qMisPeYC+QzWfrDbZVLzoqa5vMdQu4dfSe/pgaRA9MJlX
NH6nAxtUQjLhPXa4H8xGo9sabUxX4sV8xZw/FA4l4hugpH7cUnVY8wi5yES0
hGGRmw2tL1TvkCs9ZB8DqFOiL73MXPm3I8+3TB0PoUjdj1Sl9+uD10LAXUUk
tMj+4UlnaqDQe9FWdY+FgoRKUSA6ovbSmIaHzodZMZJDDITIGwg0Z1lvYKZ6
VxunSlhz23BzVPX/UvY52t3E2LIA3SFj5YqkCnT87dSpRakno5dLDMjX4MGB
TYL/VtmUktd3Hs48+bDua1lGS1n98CttNacR+m53b+pDGX0XRphGraj+IFhc
xezNw3D3a+tQwldJPfC2fOP7s2PT+mQGAGJXLSONgtwEQFA1gds8OtEltzoh
k7cuzwBrlYfp6Oyk+75Jg4wTqEeh2iZzJEAy+SPkBpFSm5u2eLCKskGzePe8
og5JaePaN1bh3qynPL3k+wuXiIT8EAfvf4nU/sf990k+xt4LTZ9PEaf3BM6Z
QxCeCLvb8jnbSAJszVxmsCYgsHN+yogSl1PmyLU/uA2p9u6t6QCZ1r7kyw5C
42ssR9bT8n6APuovYAXDvfqj6mgq5GdcYvxsZzwmtkZ1NeGhBPktjVp3ixNy
yCZu9I+TQNPYLl9vXxVUtFi6b180wXn6buYXbVkPXtQxH1KYCfZND+zWuntA
79n7YwrKcac+slFR9jISR1IMOF48QczH0RESlvXHs59/e8vneSvCX2uwGSd3
8/1bhI7yu4lm4Fgdm5BiFaeHONTsRmMaQ+r3fFp9imqLYrmmOtJS8Z7jh6uN
0QOWx1A9VlQx/2Eu296GKhi71dlHKOnSbSZp5CyMR0TF/JnCzvw0a5RpBMsP
D6I11G6EiL+wSgOnMX9FEiaZPiPaXK0XbvQhSgIlrJvlGkqKswbfkxNdZDMg
1YbWAR0ZlJzRLGDqxK7AkrN26v05OkwgGQKp4kuBgODOP8OxLjGjvb24Foa9
7de/spI+/rxHO58XV/ZHKRoPucRazxR/oyLWaax10CBXHZfFWjgZEdMCJkCU
4OXpE3z9UeTCuc6BlIf7ozpTqF5zAU1vhrP402Em3SV6R2192xqVLnLD7Lov
ipDYYUBFLKevoj8kgSbjyRiCX0F/9E+VIFnGZyrtWC+PvtyiyDCAWEmE4xBp
1BsKFC/m190JN0lXn4TaEqn4B39Vfk/TsQFsQg/Etx9CL/GcoVaoc7pJntHm
Kxt3eLsD/G1wxe6dDAOpZNcPMPHMijG6wAl2XoBuj36ahccDLnt3b7KmmjB2
yYHl6eXrYpXybyhG6ggTwjqK3ehfLcVEmmM4tCvU0vxGvV7+aU8x8W42YAZ5
Ob7mIJrYAgpqYcGS9WjsObZCJ9gnwmNShDhDxs5m3Uot+G5gA92dbZABGQ0W
IX2VQmMhWQTtGHFmG1TODJMZAVMT1HgOblkWUPTCaLR8S9FJX4wr08iquDV6
M3U3hHhqkOhvJWWbrZ49PlpQQwgsUtAuNw1KaLaswt6vLXWH/yZ9UGPwcIVN
H8xMjvh29501gzv5V5SsKhvt2BVaKGsgohKm6rlFcXUvOHJzhvcTBvJhjQDj
/FL+OAxpYHE9+79eEY9wHfZ09CjlERiQPlhKAz1snqFilrx6oiXm62ReL320
E+a+vcJrWQ0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q5NymhoUOQYn90+m+60p1pBJ4mO/qUEr9LeXzlfFVIlO1BMpfNXTddA/yM+YTZnbgy+6OY9TaeB2Wn1nAnThuOP/gfTDXydkoPLT81Jm1zBlJvsNCD8N9uNNqD26IC5PVHaHGjAuIAS+rt0bOmzay4rYE1Ptncq/1R28s0wa1Pbdh6X5F/UzxiIIFOMNBhv1BQ+NIMDI/bhPgAYIHVMygDZXWB/7Q8b7fb5DVQH8oAPR/UXsOE6vJj/QHUp23qSW9RrdRV6Xm10nphlu27Wil7yJisMT8F+EQ0NmewRl3hQXFZBS6v2WfnUVVNQdP7E+glE01TtcZ4mg+S+tPJzmX00/uwFExl6dVuz0QsCRVJu5T2Rzthxs8mo7VwfXZfprOpy91qbidoNzwQ5+1pLZ9LNFdtVW9qbtPWB9hUvZSEPk1/Zmeuv6pYQVgSGjFuEhX/zv6JysM8T/UYb82BtAYmkAK3c67OvYmjtjwenFYc5zWd/G0c3q1N9619Cai3chcSTV0mVOav4jG40UPAYVOun/saBHS+QwXz1UvLF0MPGMGhcN7KUBf/rKI1qyYRIlLlBJhpl/yGiUIr0H/pLa6h4RtfOL1w7tvmGl5mtMlPVLASu+Nws4wFJLX3NrRA2gCWz+xVGyIad3QZSjc9auxksEfR6uHnDtzREkSwFfWLDpv0UgSWhvLv5qWdKFZtYeFjGl33cEUOpk9Yvai/RcTf1LHJoYrgBxNyLtb3YrSyEMvUTSQ5WpQbelmRZpK3vEdjjowmw3N6dhH0CeI9wkab8"
`endif