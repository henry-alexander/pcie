// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AoRDFZHEWAu3P8u/2AFZ9ZN0u9mZRMjt3qANqy7ZLuJWNT/pOs+qpSUN0/G7
mSOfdgqV34YxcsJ9hH0g5veqQqMZEU0rhaOtMiLGPKOponlEdv2ssnuv1WjN
R4NedaLqWYa9OehNN68vmiT7N6ztm+/Xnd74dO77CeHuUO/IWdKh4jvgoMnU
YE3zFtSyz1Jhnp2DTOiRIHXI9xdp+FrvzFCu5IS5jjowQzaCiNc6Nv2wn7xg
gReHqBQ9OJI87EDdNdH0uoGN1RFylDj/n7rxdKWY3psWin0Wy4sZAWJCRyQg
X46xuu8UxOwAtjlH88i7lCPmKDgw1k536Q7QXSjCXg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cegVYeZrEvDxq1etR/TpB0U6ydg77AiaGLoYxCcrhEaiosiyiW98vxDH9dIp
7CDCzPHqbz5SudDWSlK7mnZoW6R2KHkuNxb4Xq5U+kgw15ezC1NZt+r5jJuc
H8DAvBqwlN5wv+xc2BL/urNkS05V9cTAdyIlF9eWf1hmFWnqtxHqxq4+3ONq
rLwEqVYuZRgtnwsx7FuYlGbGpBg2mm2hIJ2HVG/8gt0VaKoK1HTrcZ9+eh8e
1YHeluOJoKNU6S5uer+sIIssAqul+iVZjuz1cDaJ/M8wWlm0nbxEadx1+6zS
0Qagpas4iNotavsN+/zXBkfeGO2UG6WXgzmUUWQCpw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
NmMSySXbMgOueklSZrLqEAR8e+C2CQe/QNrgyoemhISkvtxoakOCOxvFLcc+
NZzsfpgqXgs8H7Tvqj1M1KWeXh1xxcSOOXLkISfJklkKH36LcS/QxZ1lHZyy
x93Ablp/lpRFv9Pdik9AEJarz6NWT9TAaUydM03Z6u1+Xn39BqNs/Nnh5uB2
QzYak031LVTbV7ankuKO8X+pX5WEka5hzUdE87kmfFbzSMJf58wr3XGJO6jp
4ti8ba4WmiEPSbu6huxjW2YlDBkJgHjs+oEIU2WNANa0jIGvAePwi6ltDewG
ZJLORsStD39UP6k0fzc34Jl5Aw4wmR56ASgtST6mkw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
a6T+pX/Igj+W9lVdX8n9u5ppUunCgCmN8IpFwDOtc8uRs/7jgeNngumtoaXO
Nnp2rdZEpEBr+Ka7VQDwJsGkRwnrnmyR3jPgH8amwfwmVFfa2Ns0gvUIg00f
3yAx5Ty7R7CVZS5YrTTWHMFmQzTvsUgzYLciGEA6jTExapz0uW4=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
K9/V/v7qayXC3Z0BxP9w61Kcbe1Nh2YPc98wVyX3rTa5K+Y/JHUiUavf1zwb
cf6Nb7q9JBBp/L61t6cntTFrNw+LIw4gs77jLQ2lWPkiSuS02P/Ipak+Opc8
W5tEiuRKm8XDckm6ccCRLyXTdsvl5MrEycXjtii5cEPy3I9YbFr676ILqbNf
rAIT27048BAi2FO4rPY7THCodOGpOU3o86uuDZv6f7ceLSh90l1kl9MMJBKB
NupXedwT+J45STPnon8dffdNoZjuR4ZkTXePM4o6rsJNvq3yY61azL0QdMBW
Vf0OQ1d9s4izF44pqNgRYwMVzhu/of7T1Sl2C1/NzFvCIGNRuWhFh9lMteXO
4q3aTdkjZp8/8Mgrb6LA/mTsy/VPACkgLgg5iUaoKFyQd1RoAzUPB1xGg9W/
I/rGENNTtWHIv/AXostcnP08q6aL8lAaDNET5PH3raWSx0+lyznqflgYAn47
vVyZLuvuGsvGjkPaf9+gW45LBrbrH46G


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aRW0hl9kfcskFFAwAt6cn2D4IJJ4YvCuQMGxqo3/xWeGvETqcM9q1Cph/sL5
7/FD3wBlSznYzz4wtdaIMYPWzWDe5RfQfF5YExoY9xrhmbQAvv6uVUaiyDJA
m2yvYyo59SLA5sOQwgH7GpbnJBw8RDqTjwVP9ZR3z4SwfjK8LPM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QGa9norYQjaZrmlF/2Yp7bAbWocD6nSxwK5rKRpGuX6e75sxGE0W4Hk+WyLR
kiq8ZE67sJ52NrSuGKYIgk1uz8qw/Spts15ffYQBh+heLKE35lkIwBmi4pTD
t9NXezLX/fUry4B1MF5b+B2fu+4UlVfj24amLgw6Jzyz95nZHQg=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 50256)
`pragma protect data_block
C5Wk8Jm7t/SES3mynq91ZUEhl57F/ldkd4+0fZXq+zmC8SXhqrakyQ7PUD+T
UcpoXaPg+5mDosy84qxu8P/K0ecUOphOJxUwB6hIQSRWflA7UzpA0Fk/70VO
F5OxyBbK6IlhQUzs0Xh9AZ4ootlqs6a+rj9jo95kUpJWS4lRbQ2PJ/B9sDKD
b0pbXvDPLo8BoTHafPe2Oa0Hv1ZM/UTE6J5kJbczKvjTOwVfJCB4PTzWq2IJ
nDC2vdmDyUzHLpXQ4MyXPK0Yc3VrnscOl101jzRBKI3G9iTfe354guLnevpQ
XlWyasdSRYMgcZm5/U43n61yGvAG43CgSGkJ/+jPyXeErE5rKhzha/Q2fsFd
K80I62jnWxvOYeh8z8hVGF+DUTN8NiaR6UZk1IXhD3q3iKbzKI8OJ4XzJtpE
Ta8Rmnhi89qC30MsN/wQGxJn4sR64m+WkVsmzeg0McXJA5Kxm21iDVFrlLtB
Mvl+qTCskreX12C0jGfI037ejeP3EQrzjFkzBhxahpUGVS/sK9sfoe9xlCWv
bPwDpuOw/cHfwJojDwzGENZs2yBC8keDaVtgX48fh1DL8tNI+UqLP9jY4d00
R0jJjGGNG0F+7fAPkjbrD3itn47oWHW+VvxqyRxlu0MxkMUCG8JfrQP8b3JT
QuvHkGl7AB+pVYkm7z1/dVsrKL8niS2y40MZ2/9ArEzmVbJD6BN/2OuriOfb
7+M3tya0a20iKtfR97CAMcnetFsqilmB+PAuI/zLtRZtbfn3VqWdrj56EB3a
Js13Wokt3wBfxDrkF2BKf+oqkd3wCc7emR9Bii7b2IHWajatDULnPBIcvL6Q
9Yl1W95AGcDk38bSHoC2uu/hO4zcLDs6HXPOR3unZNt5M1qZDLkTRZ+ktyFk
ZBLrl7i1GLioVEppNtX2/GoiODMTdDcf/XsxSuZVxQc8jME3vl0OxR6jQ2XQ
B6BZyIEipOdXKCOFg8IXj41cMYRSeuBlGYs3wV5fMGzXlVuQ4FM9OA1tL/zl
oSnZ8y/qxKLt00HKo7x2dxx18Bksiv+3mOgUybuGLznkzJnlXkGOpLJcU81w
filD2pZDt8fwnQcFNROeGljjpQjarG1rSTb3awXfz6Z1OyI+An4PverXtVHo
Y14goTi9E0V/Pwbd4f3O/3IxEOCj7VzJDnLEcrs1B1BfDAWYmMlz+iHRSQl8
YZkLt/mAiIcmflCo80inrywekXczqsVh1RWSSNQvMnA9HbYA0sx/LSVVd9D5
Aa/sP0sYZoznn89oov1js8t0Q1kT/oWJP3dL9LTwaWQsXcr4i5HGLQH2XOwt
Xfx+MMU4XR6oCd8vKyAFcQ2affN71nH4be0WBS0o++VhrbkpQaEW7/vI4Zs0
Id9LWDyoYNFcW9wUe5LCYK6/pdioiKrAd3WzzYiOZRXigqZ9MVQ2/RLx6AEs
jRcgtjtbBGVntznChAD5rinI4yaCGfIcWtuxyr0k/sshsbd0ObA5IMTnKccy
YhIjY942bRoMKiubzVOj7VZD0gOlqoQ0ntCYeWeb+ciuycL9fDlDTBkzLZPb
UHTq6lpp6vSdzA3WgxJ7Ev4hmsIOqQvU+JccqSgt77atas8YXldV99djEbfv
OP3w5iFtEMUeosXLjt3Tp+eWQ+Y1XTyoZsm0HjMZFi9E0+THMtOs8vOgt0lk
HxNqCkLVgKhnZnt/WTG9sCMoEGUHsMhisZehoMweNedpBNhUGO5DixdwS8ll
XS3MZwPt/clJ2SPjG6nnd5z/sncZZhGn6ALqKMQlQx8yMyq3e5uJISzarlkQ
ZdxtIgOlGr+a0h7yaqcrGZXeo/XWhxPJi9NJJ0aUmMciZ6Lctan+96INANUS
9RVtZodASepy2pZOGWNCGHaJRvgAgFMV0591k52nA0+ZPs0Smr+ULLystxPT
0mJktfpS3sv/XxFyqu6eSt5kOwwjuV8phfTQa6WeVVCnt+d81D1+bOcRzHy+
zUlgSz5EiKPhPcI6Qf8bs287VpSH8Cwc7yzR5shzEy7SDPgFMepaM4WhYwPD
ucVhLGmVsZV8L1FKxGCQhFy3mp6KOp8dO+U1IMAmqnRLtUDfwz9HQmjwE0MP
sOWTVRtnv7DSdRif+Rd94wvQ/uQEteKRmSO9oZl1nd9/4gjAmYo/kxKfIckK
pzT18FKUmURZK9heGl7aBZsI/pV5A7NHlcgf+dpmkS9klW/KYUbGeKlaPPQb
bv88BxfkYbgEq6wcPwUXaZ9dbw3RgixrH4gtw3Uuj+7mM5O6iH+4te9IviBh
oZmeAvLFQn6q6Bh2Wr9KuKJfmRhAM/6qu0Bmkl1lhcB8uDemHZCBbDZRGH42
BB5vld//ZOvtyMUY2jVx7WZKkfe2UDvHs0OIeObpzUbJdQ/dpMfpy159c10G
eOYotbXWC23e8C3gORn9koj+Odn6yh8qZKtd7c7c04cO2GNj+5x8datRuwEp
jTLDwXaLMP7W2ELt/t2jTI8t+9HZSGPms8F2Uzk25ctd8s8UFMUf/ODQnnGU
O7SQL6/dVQnhfYlzBfDf7pnPSaKi6rg8eDim04zcZ/C2AqGnUws/bOnaHIlm
smEJryrqf5yr9zfS5QaDC0iOmbW2te6VMWXWubfxxA4BpBZ/AnwElcDY3ybj
e+TU9BcwioiUjPexqJeHH+OmABA06PqxRvKKe/Q4tOfyVsK4r9bi6GoqUXYa
PFgFRYF1Rfedc+VucPwKnSK0Z6CWMrwPkxO+y63xSU5MgowvigF1Ya7s4aik
kLb4mMPJ4dvGawGE+Dlh7nOsOoG6iSd2Epj+RL2ot/auwOcVCJO2CrIY4lR8
L81EDBe17w5DfSuVWMb/7vXgneGAPT+dlvHxtaJ19REr9smf+YFTgY8HCL4Y
as0gIebkv8TWeA48oxrSninLov0v3E5XaIZYq99b8fMUZv05nn47g+yjEnO8
AhU/jkDpgM4saJ3qWLQJgJviS7in2IlvjGdEXblhlclJPta7vC8PHrVAsaq1
dhVdNmoGfl/IfCNqlDphpYtFz4Cm9s/XewvljTyRO/OYYy1TGDs59gncxTDs
RTeZwJgc4bclUufR3KWwo1S5McR9Jv3V2RMmZD6Vg2mcZ/PjhHuJKp4s4wO+
z4Di7Pcb+XFG1A8mPU2jfUBlo1n8E94SSoDQ+VdF99alcVK4jXmsjNrtQJ7T
0SyyuBodMAmLSbs/GhXXusNTmMLwg70k/xn+Q51Svg83W/TUFesiCubwrNJc
45GLOCvI7r7MWP2st0XN9+dXk+zIvH3hn5stqAJYcCQYL4/84azbP/+Esxvn
BBTXZewvaXieHOBqieiD5C8TZIxDduV2yJSl8sFdkJY/Q3iDZg46M9HFWQ2e
tcLrXVP7r9WBKvcY/EF9u/R3XggtQWogSYr8/Ah3EwX8hr7yU8y1aFzy9HA+
+4pR/Yp5BHaA2rS9L9qaYkp+ydjsv+5E1sZnHIRoznSRQ44H6v4oQauvxTqC
DcL24PMEIW6KoPWtXMNjNthNvZrfvuuxTJXSYfp98II4bYUFEenDdUx7fp0R
AMHqAzAMdqE/+EW6AhwwFzhaNenowSLCx6gleBBRxjTdOq2vkGs6btXJw5ca
PNOIxMgB+wYREIDLWTFZDWcd6TF4SDq2TdFmA43ig8EkBztXzUs/W+lR7o2D
76X5baCYaoXSQhtEoYSkUa2eWtwHo8fBrBXxX1VZ1+XZsjUO32yXWFkMIOdH
TbeTN22LAkHqGpyMKGyY3X0fXiImq0d+hCkCGnxnanAgKUfHJl+CX6Mwo5m0
p3ewl46135370fw2cLT4HKylQL2mQHMEpKTaNlxsLq4mvXncjh9Cr5Qntjch
udcyG3nJG7Ag+4L3LRL+5g+vnFyblefLytjcnEqDcZw2mbiWsv5nKSDJEk05
hQPzlthQOjSj6ysIY8OQLBbSunrQygPxerul3dOtEDAXvkbTQ2vl2fSTin0l
b3WhdtL9EDLlzMEp9euhSMe94aY0xmgtOUbulBE9+2L6eLL9/vcWaPo1G9n3
hqbAvtBnfwoZdY7DYgPBG/uMKlUI0aHZ7qxSgpu1QiqCNsEWUGZ2pd0RrF04
gd23x7o0I3jkrlpu3Li12DPxspai4ijZdI4dKp45xEPdymO3efs4nGZD0waU
ypq6Jqp29d7veDKrYthHJuUvOaPLeZONje/NDxATZvEl1Ukaen124O46m++G
1uTZdEtYRNZfcLge8xF+agAlvIaKxJOYnLbJ/iGU0lyQWF66dPfkrA6P/Svb
2Q9WiVUFYTR+568dg7tK71qB9imNk/9RS1jKEX9fXB52p7QFI9qc/sNVeVI0
53vxVa3mUJNG7p/4woih1fRvPyApr2n6Gw6NAJYk2LbifnGNmvW6LJVenfZf
L/oOEPAspceOZzrt3aFJ61+j2VX70iTNjmmDPspfjmxLwZySxTuh2gm68tX2
rNGHQZQA/JmUBsTfmS1CFh7VDQz9M03BCK01jDjsYaQmqJxwzMZi76lXt8YD
PY46V7i3f2BZfrmXqmakp+TrFZipxukOMmAD5GUCKTdBMVWJGyDeXB3VqMLu
1gOZiXISt94tqSsfTvjxhJDdvW/QS1b7ojNCWzO9FwcDHBwMXqRYcK3S2OFg
niFJMRrBNU1fhtLZYc4nMyEmdd2sw5iZbplW8Qffu9kj2PPQkSSBEwO8Q6Xo
sVX0aMKWme1RgsQlQd6Q05f+WeD6MFmWWnqpojMXpphMAsZU47VeZqXlnnik
GzG9nFDc66bJMTttnnjpWryeghHB9lAcGZ6CItDWDmfXyeuORC/3+Irhq8S2
wrNETqPQ9V6mRlDZSFmyjJkCcGDiAUG7tKcywAVRtFVNFNrn/GiKlz6eqxLt
2ZaHKJwDaQ7xbjxI+Z9czPLHsQEad+f/rnBnbVaM6YKG1ydi5KI+HFUNYvCc
A8dwM7OZw8jb6g20sMLJZlGBt36IuQw2CLGVjzxV/Q/L877NpgzO3ZHCEdQx
7+69m32AvJB92Js/STlEQt2PoCU2ibi3OGQv/s3FmAubNlTyk8pa+odcEVn1
gVKAKH6/0Qw0T6HvBKqd7RXqKgM1069ibp2TG7GewwZZxheufs25l2yYcyce
cHSg9F5QgDJEH3ZxnP4BniVQl4apj3YCQuADzHuhr/jeevfqOMANZTe+INkX
IigtjOXTpD2jI+fX6S+Ox1f6cnN+yOmWpOWEaIRY7z33UMzFkDkaK7L4E6Hw
88qtOrNQw3WgUGqNPErHkN2oIcyWtiBm5WFyivila8r0/AUnf7IQg1ymQf3F
Z43A+Mq9RNqVRVwpC9jJWDiseRwP22hyGWDacXee+mBEPBmUfo8wI5y0IlNo
L+j0r/xPG0L7u5wGeXBz/w1DDMxFaO/OmL1Nyl2AF01d2DKmCSpohWf8sT0b
4TGHs/4IzVrvh8nn3CRjcHC2/dSFmO152zKA8OthOWLzxI5KK3jlbbs2Hyz+
W/D+VQmuHiH2/A2ag1crsjEO3EMK8zEEy9/UVq2W5LyOkLUhdMc/JIPYX56a
zbNHdK9z53QSW6kIaPhDK7lggwEP+yQcryEEZ7GLdFkVowGZ5CXJqCHiO1Su
fI2ELuGGuvqX0kZ01nkXt/MNupdH99Q4+BXkZrCjidUE3uPmCoENYn1sko22
XziGzqzm7lfmI2XBgnGPvlCZG2Y2TJ8m0Wtl5WtRU0QPWM6GAFHi1grlw87p
OAvkQ7Tm9lNzediEjS96QnFQHmFBJjI5CJgtB7TTnvfkHuqv5W4GbqirFnX0
DhKAekDxXAiLbULLTasbSJ1hzGg1ohifhFjoBH5/F12yD84kFWQavHlarBx9
l+/Dwl+MOB/Zo0oVSytlwuHvOuQ9GMZjZfpm8Tdh4MpEpQdRTby3rY2PB2wj
HTpe11m8Vs60HpGjGcAtBzQjZTuQH4jPqw8HmN82p/O9xRQ/NZeEV3LCZqM+
YnQsZJ7/kpqUMMBSdyknb2QRUw0bhoeA2+qFP98sK/PK9iIZmYIXdbsu+rZi
txwFp3V6afKxtmsgkRxK3af32Gf2gpN1XvoEVF2AMyZli/nIdeI4qSS/EOLh
Ww+pL6mblpmXokM+NNWMVawwKqzUZSDStZ5RMK9tmdZ49uE1ijkCZTbYWiJ+
nQaCIvDTzX6Dc9Si0y2PBMmecYy9if0+DHnGOrKmGvmJU1EMDD+sknyqldM0
fq4SnVx2h/MDCtAotL5PuY/i/zAJZuTVGDInKda1yFruo/I6XkXbcZgTnwOI
xsTTc+KuYOWTlPIy5NRnUSv7sllBhOWkod4SX1ZzfdKN1g3Fmihr/WcYMK8c
KgbKm4Ejm4t2VYrOg8rDYdp7XGg5tcfOenn+j6r4NHeXMwf8NCvtPgSsQY2x
0nWo2QvfFlljCJ+ppl1f+UbOdBms4YYzpD681hOIDQysTsBukskzDVsK9Ei8
SZSyaT+X6HO9KJKMeV6G34m6XgJcmB8FF/DGlmi+/YTfNsMpiOl6fGj5fKd2
wUbKwYzxloq0S62EAqkjkc48n37BUbn5y42BXBMfqxX9hr3lf9HBsZD4PU9S
ajlkS5o9LzV60n0F5AYScsDVWJO6dl8oEvePhXPcITk5eXHvci937PTYTWLA
Nv0ezxa97VOEf9O+9sE/FEt6zt6VXB7kvm3tgn1ieEo79Wo1Mhpdi0F3LgJV
eYC4JRxmLnZRiTWwytXQt5hthFryoNxaO6TehCnak9nHZzKNNq4qTmynSSQF
+YqKKQtmXbPLG2w0989xkISGysIzgPQlRnXccPtlDFCFrRfpwFQxaVhx3r0q
DAhnfRTLXwlWdfwn57vPikYm9AxBwbr6M/tZEV8FmgaxP2fRjUJiP2tRyqk0
VQn4EkJR8lzAOKAUhXDMmX31O2tPnj8grO8RSblrAUhiNHvnW18AzwDcd4m9
4u/XvvqxH6AT3d0RgAtvzLUA2a+U1yRK0ciGZAh6zG/ivGBxFZ0c8zm4+TSh
BfnWi8eJIBz44XgmA1yW16kVCogH2FuSoCEmQqf3BbsiRx7uLGWv0+v/1MnQ
bqeSX1gaX5XR8fkyhDEnrLU3lNtcYWPY/LfX/w6ZvByeHKOGGLp/NkFpLe/8
1YqnCK3MIeNMBN6McAbjZw5pzj14qVWEklri9LGi/PdA7G2Uxo934Yn0TMBa
WW6qRHWjSWKBgon2X13xwb3P2Xqz5iSmu12AI4Pn6p5Z14L74BfdoHQiDEiZ
RLQFKWXj4qMN0AYJdzby96GsBOviO1/iTdOHZ4KzFvKG/WJ6avTy8YMUJwSh
Ky0OlpZh/E6wRXKE6E4QjuuB2t9f4fjynSAhx26oQcpWrLutNmxcmSdOy3cm
YdIG79J0vdj1+IFT7PndK1+t+XTOu4MRp+sHzNwP9uo5YLqzB7lPL190cOjN
VdK6JltXfiHSXez3xqn8sV+1Rkd4ANVHUOtZt4/tP2tQa7jzCQr4JmbfaFML
D0lfKGPm6y6lDAQhuBsolwreurM8wUq3DWFGZiJtWduWQygIMtcB2cI0VlJn
N2obwIZCMC2UEY6Ei37LeZijYO3mi7ns2YJjw9us7p2r0Jh1Xj9P62baeTrX
f4FerM7WDOJzRFs/U147Vm8m97czJq6r3Abyqqi6hPSvfeKxQbVDxBrEo2mN
320LKb1DrtI3sYPybDKuMFeLvn9F7bI3Wue9dhG9wKNScGdiArrOBfoY7GFQ
hUUaGp+2Uu17mkKQwduu1oRQfIRDJ2CXRxZCdgy6TIUi9WQt5tyQip1fz1sy
uEHCdiGUiBYEPKMfRFjBowCtfcZ+DVCMpGr17kZn9//XSElk6H6BJ36YlA32
U9wQmq2jp6HFjJYuqXuDm/FFeU1XP4eHZAB4GLDcDB1qyN6JGWEX57FnPkR8
r0z03vdeSBBkQyJXVeNejZPRCQ4emXVo3CBBnpeDV29As2WM0tpxQ2nhoU4L
XiqiRz2zBU1gyTSazkgX4rgOUQKYvkiOXfGZ/LZFRMA0alXEDPzcPgj9gbgt
CODEyExnX29WKpBoWwzA5Kq+eA08L5bRE+KXhu3VWpy/lHP78L5GH6XhKbJm
K4K1rw3rVMYLKuz05Drjx55uPrjkXbILbWoh+qnxE+21xby3lVTri61jViWC
q0eAIU7WeOwXoYq9zgUB8FR1OlQqwOFH4o93nlCwhPNKxy+SL4Rj+bVy3r5k
oHS34o41iIhYBNiYw+Fqn0vcQNyWnJaiVvpMKmNFkW0aXWJQNFP4K8sSkJFl
gf7Q6whtqaQLC1PUgBNm/XJBb/0jzLMzAJH9IQ2salW0dHCy2hCI1cuCLEfq
usUtzWsYoq/VihQ6lgMpC23A6Vi02y1HhziRWK5ysZ/1gW9UFTJ2sRk5yk2X
x7c8F3sA5KT3O1Jn7ULU7sV7v6qkFOWn1eXrA8N/7k+4XS0Xru590ujOFEGJ
PT/zNKTcUrJTq5oq1lVSY4Gfh1odDYhKCCe+UenExsc0pbHQMsmPTc4kAC6i
TteGH6O0MTkVjk8jkk19lAw/wYI50yTXgmOJGF3sux5tPlF06+M6rfev6Lx0
/Ls6GZ+FVI6zRiiWVCTHcpaDNa70sTFWeCbJrOClGFYBxaAXeanb+7AbCkV0
zLekfQFGWMoHfh5plB3fT+6+ACQF8xtoBATttaKNNjmMKTTit2+w0q7SgQ37
xE22XB6y5DOMRIKLn9/XxV6Zcunk+kaDjO+nr5A8/nCfPX1Fq6IyMy0ZVi3j
sVcT8+fafz2ZpEE4/NwuSNjhI0IW0IbmCi6CcU3YpY4Twps7acTOd83fsZ7O
JIs4KXUEPz2Niz2vkfRtMUd0CkJlclLGoXtFsa8gVbuLCmnq11D1HrNnO0aP
eYjYrXuHZHvR9fvPfvqCXkYGPiCSCDmsOJTD7HJHRf5iDdVKg9QMDsL+u9rq
PEovOpkM8eUURCGsTktXvbr4zSQkhL2yU/hQVNMQm683WWjY9A9SbMKBK4BD
Hn1+YyGrGI05ugbmST2Hblel6hhFvBaRT2RkJ2teUbw9kkWY9u+PkMfS59+l
j4dAzqiSMVqanJEyDEEspqOPzlbFcfQQk84rvsOaZVDIHd07FK/AvhU9JOBl
6eZdVPrUOebRk9gNds/u03S3V/bpVjUuOM/7cn7euMc/r73WwwqIKU4BUTbH
oHcMJVTHEu7y3pCYmOpnbANC1NYjHI0aS7I/iOUK4haO93pmcn1PhVeQf56d
9OPgSG1NEObUC8DpUkpsVIjyfDCZv0R07Ar3oV4g79tVhp+yDL+OjR/5JoS1
aQXbUOltd+f3zPrXWvFtV5PZhopBgGzFO3BjCiKFFDBoTRF1X9UQ8yZGF5nt
C8i/npFoxTE0/2y7Tt43cxU8tyjpnAfsOLQjDSM1Hla1+VzDTH4J+bmCmgXc
zxFP9FCAO9+hl2QYqUbIwsbSHmJnc4P1k6o+3t+UbB2m7j11G5bB+JF0MnvX
IwEcyuB62WWpeK5LXtfuf+YOb3VKPvyOeZlhUP0Wt07FATYivNRRW4hEspZ/
iXkVyS3v9LjkjZSGzPhaRzStfXNHnM68QvNpMm+14GaqHWlAVVxY5D+MB4eD
ZndAwH29t4XcogrTVn7M37dDztxpEupF+031vC6ukDjQZL3mjhAnpaRcuo/P
660hffzv0dbDU2r71AD86s6X1GhOD5T/CoT6f+b7WQWcrOaFv7xYXgUuUYoW
AAib7aaoPaorRtAZ8KjDLTW/6DTOhXz2JJnbzq3WCjVOv+/m65GrMs6eKwbm
W83SU8TNYrkWRnCn/4/4FEivwkzz1+U5inuWKLkQRFUIpuwtDKix1tc+0AUl
p+YMana4t3J3h1iaFsCDigGcikRs10E0lm3u0GP9OtYQn7uZz+lCtMX9t5nJ
/g/v33cmJG+lPGxccL1q9Cf3WWZdvPQgPoFAX+G+OHzH4p/2lK98pP+9swam
Y0gbwmQbDGMUeGr7NvMJROOI/0x6VO1Y0TxUT7SCIzIuvAeiDyW9MJNFq1hI
0BCD5zrjRSHpu2NmAM1YU7jBiblyQI9MpR1SFMauQBuo5waedHCovfqOW0jr
Il8wJGyirQI5v7ujX104P9vOiUQKIhZBdInoEMJZKNc4pNtfwaxXdX44Pesb
nOo90DYyYaPAqBYJB6NtiNBg+I+NOQHAHtHdmJ5jBLacy6LxyYkaPkHzC6MJ
wXlxZBH2Taxd8RpHOy+AvLNfTNt3parkb02VFDG7RzC9GVqoIwi2md6LRTtE
Lmo5LfunyzYF/QJ6AnvJrYQ9QlbN+l9be8sPWcmj8ERSrpmQRkwrV8Jjd6Xt
MrEJlt5gtVkJhzZ3ntoD+iUIp1Vodys5DWj6ynCB8YI7nGdXjSOuLyC4Fwq1
xHj7BYlAfiPcZwPGD0DaSvPypO1qWQkhvvYvODXgBV82TvKxB/CGuWHhSaIK
oytKRjdQFSHRS7Mdgdoead7rjLdmYhCb4sxb9VH+GbrEBm8ArhS/jfkosm6r
RrSD9lL5DbZFeNzPY+mhn9zjeIVJnTctTsC3ydMuIh6Jb1Djlsl4H/+EctEL
4hAhoxUmhxnqo12TWnAyHSaPDVkvm2LEPnEj92K5mycFp0SOWJZBVz1oYwmR
p5Aym+7Wg+ki2qeMFLQYcg0FEo0tyWXIVNh5XQCNPgrhX3byenSyyAUBNRE4
2CrSHGju6nKbCEWyAELPO2Zp06VhTwM5zQkzrsVO8wUMP5EeCKHWQBWMviNC
XOKJnHLLTKBgPgOETVQSU/EM2spZ1IUSKIwUxLG6hZBKQjNd4LjjArgc9Rsb
Ouuqr0EcVkiigv6fup7BQ6R4rVdJ9ns46Iey0F8tS7yzzJTJI5Z9qtDgCyV1
LUHbEVzsHpalEU+lfqbvhPZECMLGesbZ3aqsWx4mm3swn4PqHJgTTXYqFKri
9nX40EexUzTpIsqZUSN4wdDKu94fIm4ERue4v2XzBx2GbcZBkC+QCBoxh/K1
Rwnu+DNdH+UqcDoYDsP9Xq+i0Zvn1MxpeCqP+8TEh/cGUoWFXtlCDfWJav3F
FRj18Cev9+jaK1FVYGvFzQcMyb8Wbfbr3KL5JbxVJ+jWe4hpuINjTHffJWTW
4ogJRcLC1BBFtzKGpkQ7S542/FnNHPYm3sJnVNjKbA5vJARhDpzQ+ejEasHl
eeaQPrvGWaUq5vZOaYtYi6/hKHVWSfZIdWkh593wqA6IO7VXARKbi7Ea1ODx
IZTl7sdASg2qSFU2d34qX+RNRct6VwShtua9NySL9BarNFh9WG3m0Hc31qeb
8n4OHT4ZzKb4MvY24ygxahSfQvvvtD3Tf37AnZrUIN4T4TsI4/SFe/IG6ZG+
YRq9/z0UsIkb9udIdDNE3K7cgwPnRLPgyD8lLsu2AG3qxmAJEHr3hBLuVCb7
8hCmkKoAtGTcV5SngJ0uQZ4qprJtYSepy4Ooc8lZcl9aulLrnc4DXXaw4tM2
f7TouNNihFSwj3JiKAo0KQ7yMRL55qtF7PZYtLM3EyOTayB+jVPLtJQAOLqz
xneczNyDyE7K/MAQ62cA6NUjQ6nbc7W3Ic0gG3hIkt+NHlH4SLBZmKlsFjFr
qSRuQIAAht3N7ETNMcbGl61FRzPwMtdpQSEtIxwJ4ahSTzhhMuCKuA4Z0npx
KvFw3Y8Ph7Poz8BRsUHJgCgUA4Vxw/qKbWTmiMaHwE8/7q/Tmvc9YiqNXQZq
H2ZdUhkJ8cVM8yd64k+8GWVaIhlLX7feNDrLh0gEU6TjODRSg97JJ/iIjE0J
WMBcPJz6Gfg1VLLMrixs3385MoJrDKSPoaTTYmVCo0BlUkbOggtoY03Izqz8
6BXYdqArizpc7TiQTyl0g0kvNnK0BOBvEKhJ1jkDUYi4O8I7uOvxlVVZcpAq
pNJa3+hf9seRkJ8ORanE1WljJOJ7vHqXqDJXbeAVM/QKgo9KXp+Bqs+X8scF
/izcQo2MPVYJtMMzFdl2N/VsB0Zs9ZvJ+BtPZ3/LNfopByI1Y/H27TowmXis
FRdAEh6uM/EY74ppinH+LqvzGqt+2A6YkPhO0UIN/U4T7wDU6TKKZJNPzETu
jawpoyT2D0t4yvVTrBoPZjjWc8MrGtdXjOuPDJCRqcUOMdTsBoucoaEixa5u
1jEejMIYG5tEjQnhAvLyfrjE6Qigy0UV2wQSJ0LoWmMBCy+sUtrKSgd3J2d4
uCRQXnCC0Uu7c9hHmScHbZta5Jwj3FsUCZxM2LOCUXEO5Ad6MzByaD8TxDPn
MZUqnkSCUcz0aILPR2OfYAjlLaj1X/o6jl7L1s6msPTVppsMrjqE9um3BEe0
RrMYR6yONCcu1b283b1GSBPHWP9GilGka3gPcuqOOnQGnmeBe5J+OlRz4xVz
CQaOgkHiny8yxptqOCi/O4IeKd7peSA89LMhYb44qf1MKQGcCdWfjJKIkJv4
ncF1whiqpauJ4izqFbtJ17pX1/K0Ud9kKRnSGGMJoN3wNuknk4ZNADB0inlY
WhtoRdK6tIBbWlhpZp8GXHANak2Ysia9rQuNu4qTed+mIAxxKptQDUW0fA56
TdBVD7MJpsQsTUQ/cSJT4GYIHIW9RizN4ucKNGtZXp6luqNcyrw19dXHwu1T
tAIbYIMHAkBU+Urgu6VL3qGUfl0a9E08Y7erdwD981w5ls9XOIyxzw9lMK1N
uqrQD5EKvuof26hnjwhZWhMvT6Mr0lV0xIgvKm8poaE0zs8EnimdjzUm2ZcO
4B9gxEi+Qw71YAHzZd1W/ZLHy+WekV6ClC5SqQbvSpBRbwXanm0rnBxW1IYZ
rQs8w7TkLHs16JQEZeqbBGrvJvNY2YGzWdM4cpBI25i/MKB3coS9DUtCA23Y
uCtYxcc4NjyV95xB5xQnOBW1oQitcsmL7pr0Z3RiLR8aeHBudxi89uirzeo2
Ztk97U0xqivLRbO9xoHx+LEMY9niiMP//ygTVuDf3A65Ny7hLSBq2FxQVWYO
232L/TL3hpTy6ld3BaLdMUHlxeHiH4aDM8G/apYe2yhPLDurTwOJkFStM+K4
gEgzTs7qRY7nhsYanHNpY8Hss2LNQ1I9pP3w52gJnhdNunK/XzXJpOig3//u
qU7yT6VP2mHtv9JD3lZNcpRu1jY96cZg2ID6fLYCw1q546nmgDNdhEBla5kY
/bCzyiZNGlOUDEBzAdjvp4ke0YT5tRK10n4HpQQ6dtIxPpNHsY4VhGf35dVv
QvEeOErRkjb2fA7CG7twZIMAqVg7MNIUT9Bkj9j/4z03rPFo/P0Rktvt6EuG
8+7/JHhIUyOfzUYzKK5P203aE2cHuJDdNOu17+qiGKYvhlU9EfOSMRwtt3jS
Ow3iIbtrc6Ki6YlzxHp64RUj8qZ583Ft4QJAZ4X9vhQyp6kRsBE9v95r18V3
D8AE7BKgMh2QyResPNvw20nsPwRUq9P2xXOhU3JdRhmd+92YptwZsXbquPow
eaFr3/Nf58m/qdv2fAcxzLeWbVM3tlJLSzt7h5t4gtAsGsKu7lifIHkFJ1xg
0GFL60JH/Yz5k2a3eOluGjYoC1fv9EPt2twZ7Tb/xEJ1+1xdB/rNnHSkTTPJ
yGOi+xB/BTVdtU0aZNMnmnykeOTCvtPz06jMHqPfrDx9pakVdFHnceL/iI4c
0/z9FPgAPoXvl4/ISEAD6Fsp4YvhaNrgQ65gwpZmcm2spvGtdNrdF2q7RSj2
XqCGysm/n0EstYgq1s0L6rPBHnsEDsUITTH2lfcWszvlnfclyA2d9Isp3UB0
x6SyEhIICi4dG/dnGlERywhUgvXD7NhooQ/SX/RBm8M52qxti6HL4kdXzYl3
kTn0mWIPpVEMhlQm+QEbnMrspUa0SnIzpMW6zCXrEaAhudMlnyLfIYmoeeMc
x6ysLpa42sAsDb1Yig18/HQEHvJayESd6axwf7DSDsVODFfb9b94IG0MTGrl
B7A1xTI2baE69js8lmj1e2N71W7yLa1b40bM8PU+k1+rrr0kcnjVdjl0lhPD
8WAv6TJs8fhG8yAuefS1iC92tNarz++fPIYiXxSa3Ne3mWOikpUblhuMYj7b
43otVKs6UUj3V2d/kKImwWIzPm3LyCq3V9xic26qFh1Ex/a6H0tpZqAMjExp
D3DP/NBEbT2rXLPchVoBWzRP9fO0ExJuAwNCcPOF5Jp/ZWjTpmevKpvWi1Ox
DfF4gAZZVoqidAjSLIpJ8rxKd5sAsPHIqUu31qTcmkU5ReaxlcD65gjoxGB9
XTz02E5Qp9Jl4mBo53QQIDBjBHXYtubmKf4Zi3Rj75XEeMseDPuLhmgXxMIP
7MhDGImOcvXhPw/Np4lHKaJNx1uPSWDlm2fm3xSGgkNqWzHI9eYt8i0o+uvI
KFeOmsxd5ohqgAXO/bP8rg2h9a2e9gnn6/jur5bpvlALqUhO6R4h5zlnSNNP
BqvFavBfN9zuyeLCwkM7SmDGL5QM2A8hzhDrsqesWSsxzBrg4NG4h31uRvze
wY4e6dqHWq7H/VgTnpvyZhfZUNAhKFncCZ4CWiJ6Qx0VsGOj69zRjG6s/TEQ
y+GUXKz3cqxl3ZZ+Xhz9CNsvBSduaXG22r67jDvpxLjGyqM2dsISXnATIL1W
cDoDB5xD5/e511nmL7m194MWWq6EeqGuXken07zBSB59b4hdxr+FMh57lCCc
jS8N9LTSSDfutgFH0QGYNER0Y+/LD6s1rRVwy8EWZpyZtY5fVEazaJ/+8/vY
j2D24WzQ3B2KWfDV3g1G6/owVPHQxnltz1gGcMrywXnQ9d81y6/a4rF0PNN2
C+JYVOjsso2/nkSUALP3Sr6JG3eiAZEhzTXSQkZ2bvUaqfjc4L8A5Gr0/co7
WHYCzqDJMLWrlh27OOaNZsMrboFPyC/C0xGeSg7I32DtO6PfKkMKWqoZyB84
ply0wBDJ5VV/7DR4WUWVxiTluYq0hIaK5TOiScyFK2kOjoO9lmVpVKNOOLNp
ZggImEkurFSgbraaqJpcIoPEUPfRwWISxjJv/zzT94yKlU1Y7S8S7vhmD7Si
cYR1WT2DjQZqIpCB9UaCXAeyCPD5Xq8k5vJ8Uvj1cZp2PCltS98Ojh7v0uuR
4Wke6xUSiK2EROmK20VsPeMr5vpc8nxfTO1plRyrSKBG6hMjndxCq9sUcbq5
lyukFD41ahOK4TFL5hmJLgPYd9OrwYYfP/2d1J4R1PAZIqRvE6lf0lv4VBIh
K4qzWhmwqsT6125YezsjBoYPn44++JjHVH0xwUi2Q+nM48otUuOo3Ez7LVbv
k8muJNGWpNTYpiEosnMeeZG1AylJgf+6iu3rWdtKgXFHPpuWG+pbYXBQ50bR
RnXW5A487jomlWCKp9IDqMo/I3DVLPLA9sHTJ/kwG9+5yIvtItnomrWPP7Zx
dyvGDxEzAOHZFrvpBT6arfHFT0KXSmKBwxuMCMlX2S/AVv+6UtqtiQUf0N/r
xxYwLHxmim7C4aw49QzGMolC5YgsQvdU+WPHpPkCbgYBq9R9on8dCAm3NHg2
jGHp502TjH7c8ShpVe3sNNcT0APQtCV7tpgJeYocv1KjsVeQJc9i4HZ9VZh7
ps5Jjh24f9lM0TJXzBdKaRP/KpiU9kclb7dbmLTqA56b6olxGNSkrFBWBK6p
gkgJmWN0ZbX7JxsYHOPyGvf5Pr2bnO7rLnOHjXWDf7t377ZlQsfQoCsWSISl
pDBsO3fT/CFggEqIdViFLPgMBKGqb80mid2jOaoh6YJUYa4MjwZl5vgmtiT/
IuNWhaVX50owpdK03SkalEpVYx+s+nH0GW+qLVVv8FIMde7y5+cD8U8Wo7SR
mWOuRMWyM+BZXFwFb8ojAaM2pMI3i3u/E4eT80vGhgJZUknlXshYY+SWk1cL
IDvvUCn7fxr5gRtPwAdWe3Q65aRrNEA+aI5af8p866N6y67/qNIno/pAkwEk
mYec/UJQZ+EtfkdfofIR2Z3aFZFwDu6NaqFQiKS81ABZloo8rZAJEDlkALgz
eEbnAuVaeEuJJseqQ//woZC6QUCMoYja+nhFMhEdYsAEYKyT8R4V1JgHB8lh
D17UvmYen2vD8zLwTLySeYkRu7UysyZ587RRwrJieNorupxX2vB53kue0gVY
LmkwkrK1Wxl7ev5M2ZlfjJr1URlWbiybouRx9LSFoWZRAuyHg2zXfUFfypPe
RwnHEAi5YhMU0CaQWr8+sN/0672cv+f0RsyEJeBON3orCzCoId0UvquQTymI
6dt3jyOqOR9jN/vPyFEWMuyWUnrbHOJ/W1yholYod6J98I6rmZYqNTl4SvB9
gCLdG97aJ8qZhKWiSpQu4fm/WvZ+OZf2FNe6Z9RE+gq2hKP/fXI8LiRF/B0Y
g8sH8Db1bYOKTdI47Xl7SYxgW3APzgARaQi62YomzCDkD23k7ruJAeNz2wot
JJfIcoSIcogo99b6+/w5kMa+8oXVA+URcv5nFKUxotjLOoTlUnYCP7Vi6I3P
ksURY+SMRnm8PA4D7pSQzli+pk7VthDCxw+ZUOyNTzSNvS7ah4h9ChZECetz
v+9yTsFS+RIX8zebJeOwJ05axq4Juab1sOrosSZpZ3RyzvqdO4xCKT4secpD
fpuOCMotPAohPdbuN85qYUPvEZKMRaw9unAsQGSQQBWnL/QleKwWOvmJSorY
vmKDkjYIl/GkrYVCfCPqKsd2pkTScn/hVZ8Zn530nuujUbbxGe0oBVWuE3fX
bFuPzVLyxoGIGrQcvzu3AWetnz0fL1XkoMArXq7ZIIbhBM0kibBFQr2yXU8Y
W9QVssemaIjc6Yr/XMUPDB7GBEZHbYXbURjANiFXh9Z/hcwMI2AQe0bWbRnU
7RpXF5WJlzcQwa5kSEHFikqiPEQKFXbcfU/C37FDreEg4WgKJ+sgVT3vQiCl
mVmhD9rSLDwZ8XIBrj/mKk27X+5GPJrRpVoRJoCEm/qTmcGxrh4e3UaUBKgo
nhH2kIfwXwT66jpAuJG2BjWyfDDnuifQOS27PHNHuJO8BQFlpgUQxWsuhAvC
KHQy2ZVCn+R+qZtynyLHSKbYPG4F90tyaL+o6SVM86WDdzVUmHIzP2ExBNsl
acsZhL7UsVaESxd8nsYMYNKLhCKy0C+ojwHOfU1Y4uZlbM+a80m1nvll7ds2
jQD/ANkyEqDh+IzyelfDa9upbBnkppzl4Lojj2SBG7+zhohLcm3+O6Za6SRI
DyhBl3do8zwSH9H5kNQN5WIU60Ng9tCM1LWtP0DF994tgWJ0ULD9pob1j88u
T3nv+L6cnh9k7Kc/BTQdVOXCetGIG4C2Aa5Drm+UgFRk5xu1EnElzMwkQV1g
9pvSQHuHD2ecKHGbqnmYenx5MyKKZywAxPzErD9lB+W/Q+5tUI7p3x56brox
EEX0+aIKJwWg/kr/bGIYKIGIfLtxSlTocDq0Rlit+WnKWbPLcRVxAKmSR5mG
z3PVzBVUCGdZ8O8fAlkk3fkb8ZvYRKxJdMZHMoEnl7nJ1rNI26sHe8/Crk7J
6OR4q1EdkQMYEtN/pnMuR3yJ2b3j1UUiionT5mUhBG+GNpJZXHRQzx8Jbfsw
pWRSZEJoo9SNJqlZOuFQQenx28uJSMzTXESuWnkhMxhiUCvj1noP49LOSlxX
yU/yTxsv+DLTflq7TQtJaRvnxUHYxHrsOAqGOEBboM8BzbJf2z6gTba9AoEb
i7uAwAM2yeoPt6V6p3OcV5A2WEQTuPqEvWQ9GimhbEqLIaqQ0798Dq9zwTdC
EQGUqpPoWheMADssqcmoAMVppl7tB1wjGpJXMML94/t00By1wNq/nw0hMBlY
5ndC162uqu5c3YhU8fzt08KaRKqMjUoyasJsH0tHbJjuBW0eJCjCN8bG5Ufd
cfXyH2eHWdNux4GxVjFMRPCHryR/qa8kNoUrdQ17S2e3n9rbOBK/IHgNwiPa
8qHq9QWUJo1WESdRudb3+Ff76Jgo9N99QqOB4wIzcrmljVx6thAakLDrlkJa
Y5vD23G39ih9UWMc70+erQ00EZHb4JI+zmmDRHXvXSLHjDdxU3MXgiM28/yU
Y80CTcv2/tqMW2gVtlhUTgx5SuzndB7OPYWa+ws6dKg+MqzXcJzLgVwF1e72
QcaBDLafaFRznVdDJrBn0fYyga42P6iJfkkWuI39giP8qhZ3saXJUe8BHYve
C0u1WxB5T/cqW6QZtwP3lnv2zxR4hSLRgn2R4ZBN7NV6+DfV+wDOBqfco4BR
7cVBqjTB61p4fV5RH08mp9czUYqk+T6E4asPRjOHQR5i6MaT5KJNx2wyKlaV
EQQ3Wggd9pUliIpH/fNx+V8pfmuoN5lRkwNakSh36AzXTTQmHnxOSScofqT1
nM1N+Le3q9ZSK3Embqfh+z5wOytgfnzxNQug5r5lxGn8fPT49anOliaLVd6r
SqD36yoOduuvIXhgzN5gKri2cyAEAGrrsMpAkjZkaqNLef1bMJe5sPh2pCuG
e8Q3QFAo5KJOWaBHh+7AB+VBcd8zsycSJ/sLVbneEQJ/a8WCWs81paxIWNgf
2OjizpQUW0SBVl8m8IsWsPzO+ixff5i9cvQamI7gN7nIy/c28UA/4IeBRaHq
5/eU4LEcdt0S3ZlJLIvA8YeZuW68Na5x3+Dk47x04x/73vLwzy5TpxvsaOkz
NAYxHiEEfqPB7cRfLOnotvpdpdPJuLdm5qb6cD3pcJLRh7PwAnDI1M2idjZa
SCKiez52Vr8hROyJvCNiXIfFaxdM507O6uPsAtSA4B1MJX9mtbwV8jK1daVf
oB3MX3wvFydZA/UdvaZj4cMdY1EwOYloTNm7l46hRrwioyKcPHpsLeYDODFb
HKl1s/BLIxyRTgfi6Hb3G84gHpLxvD7QL9zKLLXhKUEBa7c9bDBAy+L/VJYQ
+FeNLw3rVQeNTZS3lWIljWJ079IXupCXHf+7evLh7fGVadkClBRE2w/ZLNP7
SFEdUdZLRe89Jub9tfptTmdraeP04QkbQd39CDUGbW6C7/CMe+1E7iHk4jGV
2IyWhAW3sDuDIiDcn9cAYgKSI7sbhaSx1e8L0627UdwN9xVYrpCaZ4moz4D1
Voqg1IzrZ0ToQIvCLUfr/DAT5ojA4xgq/ljis5NSb101N7hif4zUERLXXUbL
NVpRZNZGb68S+2rVdUrgVObkNLESOYT282FSTln0G9UAuMHV1WiIyp/BOsLg
8cvFMvjktku6G0w79R7ITVBHEvTI1C4d5ephwTqp/pXxebiNJ49HbVA0fKJ7
Agh43sb2mxNVIxQmzR5w5i1RIeO70nbhtdbcRWHw+fFFaIpV//tp607KMhDq
fyRrCpVgGg5DcdAFPwcEhx+ts6jFlHF+wh6WpFOCH25RxZhVWij8ILnC7drQ
i3sAUbgA10zdimAoHCmNi7kJozeJNSA1MfUl7iK7UULGV++olTL5gdwveN5F
mYZGn2LyhRihVOQPyQZ9LREgY52uSdyIkWKxwYfc7CKgKGMrwrHc8EC+mYNg
HMXiate0XPMwX4+WZ7r5cNV9kdduTu/pK8eJwB+MC5rU2U4KP41+trh3kFH9
i1GqsphoM/GskZbjJq1JNxetyeEmnCEuZFc4UGXM1ya4rvx0jt2CHKExSjNM
zwl0hoRBbjTOC75nyCihCJ3HqAth88mLGebOm4F12fEMit+VYjlpZ4IDipHY
HisxtpZ0muOAxT5h/K4yXJnrvAmp1fUGydCU5kEk21Kg7dkUtcAvicsIazaz
Br8WF4y58yhJvE6wH5ZFvIYHG707MVjtDNJAy99j3lFRmkll13h126YRA3vM
B/nCFg/8TWjzvvjc9tdCzDmzIVBP6IHbH7r1veDDhEoRuM1kjNrQLFEoEI66
seMEzVkqx1XTa+ONenzaVkjjEQC59FYLXq7+1B4MG3rCgtkVHHNK+SvM9LZA
zDwMfp1GIGInwHHmQk/Jm7GiCR+XYsC6I0nsQe10LZcybWGEiMJ50jO+G8QF
0/j9aAJX0kI6C6kGZOdASIQu7milUo8V/C9h4thU1OFfd7G4XRu2YZRvKDmL
Zpo1uXVXFT0VGMB2iOKByGXzNNWDnCWEfHWwpl/5Sw936VzH7JkwEDvvCl+P
oI5GowPjtZq4elk5kF3JwcCyCwPYr326lcI4CnBgsAQ2BXTKAg/9a4HAYBHF
bropbdRubqKUhweiI9a9Yc9COm9WySAL6AEJkF8zl4Oefi8/5xmV2HtMvAn9
N6vMOQEuOEeC3NBHLz6MyNYkMLz3p3L+3z+BifRRc91d5QvjHfNkBQRH4Zqs
rHwskAbDwGNnoV8wnw6ZnO++Zgwjgi0LBaEa2uEP2ICEl4EJAjPqlNkW3tZg
CZUNLgeHGMx62I5mgOHS0h8MycCrkxaPc4ocrGMxgQQ4Z/wqsoxCf7KB58su
WJvSMfYmm0f+jLqmsG969beXdYu2uYnNrIUOAEyAqrshvIj4kZbZsJRByI3E
QsZAqb7Rkh+D5a8yIA8XqbdZyCIBKutDdfFR99arsGo9dRZyiVIz14/oYf9B
S9hvhD9xnRom9CagZKmt5A9opsBcOJp6mZFgidoYLCZWnweWQPEaMFlcKf5k
AiGnboitT7XJ9Aod3KGVD568xQCjmv/MpQvjjLZrYseu9uK0SPzzKjqDe9tz
G1svzDFYgH849Y4fcerz7zBRqG9uIBWhkix9INy+ocKngH/M1oEj+hT8dPA9
inwkGm0UlaH5x9dj1afR2HpnopTm0Qt2r/uX8KvJZdt7PhABFkwDmNdFkykz
jWmqzFzUNyAWDXlDMnKESrgl5u8LXU8nuBZu2ElOdXmXyECjhAzff83HdzDt
SpecsUaiAnGsG0SrnL3TuXDOu8c48pGsH0H48auPriurxVgHHQmeLvO1w+XX
8MAWeZldy803EOD2fGoDlZAdKd5Egp65NjgAec/6SittDHMdI5qh51SavHaM
/HZ87hKLfwzL4BPba5qodLJiO2smJpjX/Gp4yF9H28dW0Tlv6xevqy6SZ2uP
WE8iXVtSgS53GKSl6RFWjRWIlxxkSij4AKOuxpT68bigjsE+t0TfrD/mxOcb
W+gWK7GxalLDbkHBcTGgOUF43NEQW3AZFOdXAL5ne2yPW535diW0IQhHMciw
LCmaCJ+6BTK6NgPBCQzhtCvk7enJdE+mpC7f86o6uejGtxFdcrpLakSWrtPW
Ahw/jPYzockKTShYLnLOwfUnExE1MQrKw+4djJpp1rjISpm5ZLOYf4NElgnl
p7QmESuZBBsWn+3T4fYeESeLAfOfBJPXqkND1/vtJh1TWv9icS+8FFbiCuv3
ZjEjNmAIl6aXSRTB+7GCgMnN353RnIGkULpqT4kmvnw/bfsyLE/W1L/4dNf6
gzYL4iZcvDILGUPZCZWdD1km8WcEB3J7EcP7DghG1zK9uQbMhm5UJJCQETXb
EuXT/pe/7o9N2ZwZWjLgDPnW7FL8uXdYbmxQ/RmBxQWkHcjjiC9O1Tk5IVR4
MyATylqFA/uTu/FD6rP7jNfAU30GrSQHTYge198uXAB9b22QuA9lzc+2VaQb
t0qs7ot6LqE16j2mXB5EBNSHfsemZHMFt3ekzMaESGJmdtr16WEnfz4TRM0t
x1Tyep5rj/ZUdZxVJbObxY0C5yLDJCIggIOGyGnjs7UIlCXty7J1G9FVTy4Z
prVDPrtk9McrhDjmgXMqlw14t5gI6BqpbkKa+Dn4NY/itZmPbpZcaFcTeJZS
vZ5qde+YUsQCOJi6sQlISxlt8DdNseI95EQYIeQY+nU8SE4I9Mfaw0IiWsAR
voL6wl2J0BUHjIZNDrTS5avetlMLfCCOzu3us8mPHnE2rHAWc4ljKFJ4tvE4
wbKN11OhJwvZDT4ygUL09yKkodA1kc/ZH4xKl36jdqBe6oa0+Vfp+bHy19Ed
iJPbwauy/Ks4A2Dg/z6ou4u8vZuWMNuidI5aWnHNXk+QnKzyTcYkCvOFNhKm
Gv9dm09/Z13CCTqcZ1OgEWoWSlK1ns1DofoXdrzJ33Tj2w/939LsHsRseALa
c/kOgRBbMhW5YNKHuUStaZ0B78bACIyCyEdvU9Dha20gn2+DrbeAo5XA4Rnv
/6xJRbW/M3wyNb8b2QtYkhPkf7mqgHKlk03tKNVRLRLKif0QaevezHOhSmHB
0IbXbuX/FG35LSAjhPugSZbW4+Od5j8ajHNFNJi/L+Ls/+sZ2SzQVB6Wl6aO
yDu4CDcvyWgPnihjPAaFgEaRcmgsNtrAY0tQAunGEjklwdGT2ROrI9c8KVKO
NQHVrxqoggiSRTbsD3w1RK/Az347Y4Ia90j2r9HRK015JosnHYQDO8TWDHqd
PyER7DTvC3d9tbma1bDIpNhhAE9m+h52Oca1cH87Dk/7zsxnmrVQtCxqsaFn
puccZaR7RnpJmeI2AlG4+1h/Raywz+vOBoQZOP9gep8c0Ok3hwmykmT4lj1I
EhWToK9du2MnZAn18xN7AyVNmcG6w3OzsNqWXsGYd/jkP9eTiyFwYriEYtIG
5Wd1VPWiEce5GPgSjAfrHHy8dxkqusUHebQl993if0txHUeZoNTIhZpIUUxl
uBLdL1erDyufZH+lXNJhX1bOJokjhTg4PYVbRsxC+Hcaq97UY0dke5wkl72L
Akzh1EOFrA9Szi/LBBtdDc/RAg7b2fLNq1nAawpI6EOZ2XlOoqv3XpARtnia
RmTeg86aqXWuCLVOsr/g/d8ejdc6TJ0tBBgtgWF3XxVSjxgyFWxI6CyYF5RV
2oI6YiQzMLrLS+dpOxutZ76vxzIAIhUagpw1e0yBrSYDHHNiMlQh5WNFVhBh
ZzKuOBpOf5dYSdB44HBOM1CAJMd9xteiLRSUUwXP2x6Rj+lEjOB2YFOQ7OxL
VtJisp1QZt2zHqpcvmY+mudVGkoJkO/rLwEkvTa5cjE6b6SUy2QHo92eI62Y
ren4UbmfCpTPYM6CuJI62t7YuONa8mXWINvB8W03NKg+zqt7XaR88+sjoAwC
Njnoe1YdbYDR8SkcUSEyVasAzg9oYRuHHlwQdjnwS+LrRm+qQ682za5SzyMp
48z2dri0vvwZtikqx5a68qiMgWkLfWkQmtXdjezy+ZIiX0n+0JkHzHrMFKSy
XFqirFHAnMWAIE/+VkekEY8raFzMfxbtG/rc+HFX5LItwRFHWLKV2leM/fuL
RTcNIoGDcj+GpTpMU0910Hj8HIov480ZN7LYMlPXwUF6GgLdVvILBloDm5/A
fkux0ZP3lw1XXftJAwxjnpZYj63RKiu84kjToSiua8HXCxZyOiTeCUU1EVTI
0zZ7Ep/79n5Gp5OXsJOiFcZTs8GavJ9Ei5G8X0bj8IbdaZJPPmTstS7W5Ykl
eXZyhUBnvk0SG2/Ld6Y4uEFS83gYRQQvmbUEc+5sWBmImh+o+meRo6XyO09K
TvmPMzxdAbf/tAmORrrzFdac950Yrd+Sbwnx3AgOStXJeYfJycNaR9uIG1sq
VvA4aNJSwPPo06LEoGvnP+Bm2l+hwJBfy4l1FsTC56Fezaut2mG8UkdqG/3C
wq9ZEIi4/+lBXgM6gyasX8r8zhB1q8YZf98JDMSOyYo9jI+sk7FqfHria9/b
uBcwdpcpKne/5e8W/yfyT+gcpn6uRNMOdFoGSW2PRGqpUKAG7mOxkWsiXwJ6
d76mIsf7UFE0PCl9nLzATcxN+tHkVm3FM3Z+Cviz4vfTGLuDqbVbD+iE/wHA
1dWuuF9y5BEgbOLZM3ezdcGsOGY2ZVLw6cmPbPmSLwTCkBWME0wJE2Lu+xh0
Va/I5tRQuenXS2oin+y1xNpi6/6O1Fd4aEuqV1Vzbm+g/iFcf3+jxYNsAHFx
8iMHir1t7UVKq4FNHwj8p6pvbLusuO6RcwoAcncfSNEyvjdeV51evoAZ2VK5
zKbLT4eTS5Gc71M4LBbPgWRqxcMeEZJddXyGPhdKSRAc7CbhJDkGGGfnbAog
I1JxDaAzLqzk+CGj4D0ktF8pDcKxixB+LKSklrg+3r1KdqkQ2zvKrWQ88//E
zA1WNHHQw7g0DTC2vYS/xj8LaPANdS+j9AJT5sppY5IY1pKGX1VqbnJuHF3o
XW2+lrJMxmo8+FtzmZwc0JmZJc9HwumjERUjvypBFx4O7tsOqfZdb+3BFatX
ikiDH8/w4aIkBkr82w9cWaIdvcN0e307s54imf0GmspUfeWZZVymhHu5SK6a
K7fb+DPj5tRUjNjflxajRemaqRsdNWrB7u2o3P1CzWe20rFJCqTngbbF0llO
IWDRb/TdOmAURe1mWEXAf3L8kwc3S/CcluoHcuDaf0uBHoDiKlVxClyzHW8L
GZOvB55+sGZdUb7j+3/ySXxNTx9+Zf1HzfZhGnb3OKD/XSWPCkQ2kdK/5k+4
s2B75R13vX27l8emj9o12BIfr6ob/4yksY0o+xQdQcmxORRP6yYGJzOb80s2
zwaQswXpt9mYpVH2rFihnOD5kUf2zruti6PIbbzQHwgYVPCgBe2s/kANFkEy
aOXVLvWTpK+hQwO6NHDTmyEgRLrOGPu6AHd0OIlxt1Tlb38HNCuNcXLmldks
X92AuDEK7qxHci1hJkXaBU7CQTn236GgE6Y2f8N1JKvhQEF1/cEx+E47qlA5
kudiDMHN9QZ0D06U87yCLWIPPbI1dL3u/PBH0Ri3VuVFjmyClajtuOycz/zm
cmrN+UvzG+/fMK8pdgXhGsHnoJHz+oABD/mZ0XPk7HEUpJlt6zhvnFJUQk0R
8cYlPB/JawdnCLuvcP4A4wxK3fDV/YqIUblu/RZO0bVCMX9e/KGrC7dRRl/+
m5sVV7BcCBX7SJ4D+duGw58fq9kQTAVG7kYVjd8FMOKd/nStulDDEmmAJzjZ
+d/YvlqsRvkreSI5DMzJmIPHY8lyOO0/jDF5bQnbJGa2b+e8UtEy/rmhOS/L
1dBdGCx+vjBVQZK0RwPXCMz1qhix+5Wxa+ADQXKbTuY03evwhk2+WYZgDs0h
C/OSCrcPcNcZf0TgHcZJO5/LQNcDQKQ/wbrud8hlf4k+I7yB8cFwudz3MHq2
8XGjLjFljvDFj3NsO8jx+yvBIjfUpY9sa4mIKGGRz/Jmt9NnfgICADaJX9oe
0c2/u/dzUW9whqqZPc980BtmbIbzWt+JWOV+/BWD8XmjwnsZ4KxAmJVpsP1v
ktE1iXmQ2iD4If4bJNCzGUnaUSIE648mSH/22DT6r8nYd3xVqyvW9gbPcLGA
LIYYHAtYeLkT8bncyaLLl0Hg4/cAC4XHftMLRXO1s5iz71TusFwn3eN1aa2i
TMWSqhrd7swCP58nbSmGCI0VT89il4aKHL0zmubcQNr6itHMXn6t7PJ5mu4g
nsD74BK5WEjIV1idTM0/VgAgqrLP4+2AoOvFhCP9o6aOr8Ovd68nhBZaxB78
/5QBFZjOxMAbYgH9rdaUsaR/r0Jm0oDlizhi3EdWbW4MTJXn5UULUY8bwKXN
ueEmFlgtaitOvnlgx18Uhr3llQa3Ov1ej3zWF7lL7zYNtLCNRLsmMgJ2b/hl
we6+dAa+lBQ9sGAm+pr25Uwyt661688MrNEcH1H/EojXMP5CbCb5nwHM5f6L
U90xrKpAtyPDhtpth4IQ51eU84xnddQtlCzsw1NeoY9EPFAZT1sChD1auN5u
LoLuBPEdHTwbAQY+y6lsdBL9A854/yL1EgWEmc1B787kSqVVPOKQugfHQS5f
LZ5PotkZB2tVtH2AyCECUk2smBei7BnV9IAuVNF7+gFbwoh+fdxNdGXCWN9H
9D8IOdrnCzL9tgtkhF/SIZV/9PWe/zR1ziPZ4E1vlAJgOb4zMgeEWkGLcA1Q
NWomDnx0bm7mVO+zs7lEzDONA8+lbgr1ym5A9PU/SAOlOgjSEV4+o0noYGTe
EXOVKdzHzqSCmpJYhWJHFhV6SOb8NMuOLT9kIpsuvt7OFiN+7c+2y4ItokOe
Zx7zs4wB0J8/HnbWugvpiiiHVopmMSarfMxxho7o/AVye3ibR+waJ011MloT
UkGwJ82oafy7wlX6LSOiZZROl+dm7w94bFNLpMHEk3RSxZtDjcVQNBG+O18p
Hc9KqXk5HDW+VZDnE4pVuiFZDG8JLnm9O+lUM5y/Qx38lceamRRPhzQa9yiT
it7cxBjsD6Kd6nFmGdDLevq2icRxhJgFsGq2mkFujzBiV0qivx4vq47y+GSD
NRwpxklg4/jBjvrazEjaPRLyrWT+XCC8RtpmUwX4jNGYu5+4IkPJfWOqAUdc
mA7T/oaq8GjaNPLuyN6aAY7G2eAPRrac94+01PDBJ+A4Y23Msg9BksprCERM
64L+iO5qYHQLx6/Xe7wemMmHRjojOc+D+KBSLc4xP+4h+zS+0+NJ5tC64mvZ
PkCdmFaTbVUkOx6tn1wVI4f53oZBbqh6kjTsN2QR2x389X/z5+TucZffrbU4
HjGYCxE7LnC0EyNvqifUVPL2cqshudBOU3CfxUdjPjDgMAvyKbC8py/aoOog
TT7bEWhyXwl34d4IQOFW9D6hZnnynKGX24I6qF8qKNVA9n4qympCSwK23JRU
QmILgEOjpdHiOOFBZiF24SC60uZOVV3ZZkbK3qu4pbs/UoykcvFBhCgq9GDi
tJNtyH4bLplrtjtln7I8shg/SBYwZ4IsoHvkW8yrK3SfwIv0EfKsXyYz4ffW
NyWvILlWMny1GvufF+FMnT4kEXUUsaQWznuYg35ir1qdG97GniwAl0CSFmA0
IbJP0+9fuieKaqn4Ksc46czwF5AJ+uupfLOw0ynijE+18f2YrrsOoelqWBW5
hkiM3jbouzrMEQTEqNNdUmXcp6M3j7G5i0ZMoQddlxF+Q2dZZ7EwDPBMer84
BuSsvxiR/LLypsjO3lmkMPfloDwcqMiOmBmPdVLzHxPO3c3V+1CPV4OyeHV0
YMvoP1oFJtdr0twGL8P8Ds/qieVj0iEXFsKKUKdRYmYyMiFNtEgKfjv3svrG
4m2QzJnhLUuk7dVuYS2Ydj/8EFG6SdOqTS+mYvXM11dL9RojN8JHCeePhIqg
dIHUUkEXuibxFKjNPOxMK48On7wx8fCfGGWqUibb7F9Xz5dKX+8YlRw7Ptly
NHiygODZU+PLlrdo9BRAZO/YiRdjGR+v1soUyWc75CTuxcCEeamuJHQtnxo7
4tBJWEVx3N+ytOckluQbHQoDLZRO0D9q07aaCGWx1JNmDQn6Oxj6LUNcsY/D
Isw6YzYK/FEo/jLaBHgvsZavkjJY3C9zucX1JHf7SZX19iOUeNKqyLm/Pjmt
z5aLJYym0yoAqt/7bI+KPjD7/LFddjo0h0Ai1egMyj5QBFHi0Ip7JYmy1A6t
UNeCWTBLiZppHwYoB/P7+sAidnuj5clj2+3xND28cTObid3c4r5J4T1pPDNm
18ZlJwllW5YcYC7UflzBwJPCmgMxFM4eXoATJtHQpATJc2DR6c1j2X0lsJod
OBS9fgpJUEh7+zNxxn+tv7vgpi9ebxeJ84uvwvTTpmPC9BCcYOyiewBoWAm5
4cVjSHJQIesX0MWujDZlxXeNaG/6NBExxdd4tqm90pJ67zEe4wJQ3zVjNhLB
3knn+sft/EBs8JkS7RnRTTBanL34zXD8ji4iJURHJgx8TtrKzFsDAA6MIYeT
YZwyC9EL7rGF9QUtk6T31IvQZfUG88wQ4l/fHbIRF/WK33Yvrq5KZeiDglkf
YslkGrfpzEHf74ncnW69myko9q84qmKPbZZLHVf0GrZ0bcY1Um9zSQZO5fht
8ZDNAX/dFKANVYBBrzvXLBx9K8xFvedL5Y6dpdV/7hD6Tvd0YbLcvdEXXZuP
u6xlNaJ2fKdAC59Cwv6KOPMOvLDIVXXUBvcKhk4knPTQs4G4B7NK3VtKSaQJ
yB1gqwLvf0H/BYk1DvqCoORTZ1XIYMy0SiNVDrT6gE47jSqOLtN1Go68yLGe
B0W0yIdZNsR4kfkc1UpHPxyjIpuNXY/Hq6G8sujcDMzqvw52dhyzzLlK0ZyE
oiAsouh92VvRsHCCqHDN00tgLumypCsZYmkgCDigZrINEVrw8R2Y9TN5BBaY
zlDY8JAENzuEbiA21AiPOXHYQMKxMlMZf+otxnobfa1pzZg6kZANzN4q3THJ
cmn6zLlMKjdTBk+rimyJ57RJwaDq/wrlfZnpeAJI89suDJKwQBOBoQn3fsGM
WDJKmwb3W2/1/t3sihbm9xLqCR/5hEadwX65Suxf+HI6WlLUaYF/nRlDW78X
MdXs8HuzuVFOaNN1kRQrOUaBx3RNWo4DL0MpZ5pxgbPTfgRWgrBPO+1gFy6e
XQtUHUlF7RXW/76OKfvtG8EmodYZGbQmrt06/w4rgj6KY/4riYooVNxGjz6/
CmEAiSTldKGR33Ym7FhoO6Z72WymminPeNH9XDZ1ReSqAghSg76PDtM4FzCL
twelxgOwAdaAN5JJi4KWQcPxuiVuZmYYWM22gcAhOWZR3ZskW+6fU/taNO30
yQSU7Mar9PM9BvzdRB8JzjRZRMJZWuQl5mjqDjYpJ6nQRlseHjUWKY817lJL
99fWWLPWzWFKBK3Lmmbmty0wRscXko9upwu2DUslcPQR4uJ7JLp3X/0zRl0u
q/ngrOr+n/bngo8a0FCECgaZu6zNZyG8Aqn42BeewTuVtFHLZedAN4rnJTlC
BOr8h1jLdB7yogLb2HMLCljQlfZpToCWJ87vdBKV0j3G+66i0uMuwSBpR2LA
wCJc4YWRKkEqutrYMrOMDqAC3AiY3fAWH0MQ1u1RhyFPfYKQXMj1FwQYeCzy
X8CzLT0qYVSM9TM3nh4jjDNzELtI6PDXG7cJUcZ5qYO2pg+wW74BrWQBPjJ8
8iAN9vvfMUSyCx2xAVuZmSKbHQUcLK9GlKfGnkpqtxN8hh/9Omf1Eai/17Sf
dCCr/bsqAvYEmcAL7vUhCIsCgoUu/UQGE48RiuGdp7UMHy7qe0JBLLLSHQTr
pFwz2k8z9jXVxyy+JEWMDDdwodwAlnJSERSW50Jq2oYrAQN5FFV9Fl+qpNKi
6aanJiMEO2zsHSF3AlfURUgUv/tzBoY7OpeWcJ/ArqKv/nB+nuOuro21KWs2
q4yxoQEy800AWkyKg20SVGTcqvFBnQlnUbXFTVIMPnLeGMWWgqIQSaFTkGjV
O2UdP49/3j6YUVl/C/3pPZhie4robA/XG1Nj0KIGweeiZHjSDb7DmiJRSIuZ
v1BCye3GVdd4Tkt4Jlt7/cxYufPNel5Xv+dztnAUvCBCI/3hH3Wdgvj38EtD
RN3X3aqwzrbpO0hLGCYHVoV38Rry4uIQtG9YsxHHrqBJRfHLItrJU2BUn0GY
jiyDy1RnO4y0BSfIof7XNn+LIqz2umMBn9JQMOonuxMR7nEkJfbYMNTJc5OI
/+7UYHFhFfqeM/FB2nkm+Hf4gF/sJO0NKDmILgUAxbMpjZtAmF3tFE3LO9W7
KwaK995y7zLbX0XQN5IHOsisluk7MjCPA9d+yEkMGe6+mprJhF9t5kkbuNRw
MBFYgtsx9PlewNdXTfVdKAJVGREL/s22C6u9e4dHU/9UfVzNApuaiPps6Ss3
HpsvioqvVotVzDE8+DWRNxnIsyFKYtI8SjJTXOCxzSKfeYRuTW2rMqAndY5c
HIjnuFQZeJ2hdCwRdaZb0nZBcDa9ZmGdSdqatpdiS8YdDc7fVj98CZu9rlnm
WkXQYWbClr9joavw97ZRhgGsQrK9l5Sw/dgZ154LW+6P2KZVYUOMPbgua7KA
4QqjbTjMr1BzTWq/l2K+0HuOrNVjIe1YEEdB0XMvzHBg+QvgbQ7jTdCDUnie
2q1HOKvZxAAaIjTt2hiVZsKfxdATHZ8wVc+UPWZmKuht7xLXjSv1UFkA0SBH
MqX+Gyvf+qhuz2/oIyVxxbCh6izE5Q38/DBVgx3gUXkBKZy/jT+vNXGEv9+p
Ej0/aSNC9q2ZqjQOrQCBiUEQhnMKD6Q7IPWKuZhrFkg/IdW922NvQVEnucMV
Lie+abmfp3EnUWA44AJMIbzfh30skTG5fUvOc6ek9DQ9qDZJ4thdOkXpma0y
lb4Lvp6BsdobuW0vRj9/FPPsuSQvg7K9z+HJEGed5rK2hC/ywLiHB5fhNQEA
/0tigcYywUhVIkhat0bfq3carWSbzP32Cvn3kEA0F+fumJOc93AnhI1iN9Er
PqauufBQI/wWfwnnmEoU5tdq1EXMXJrMmqY6tifWhbyFN3IQQWu71TCZl+K/
rlf0iBNEufL8Ktzm1Xbzij/ctz1pRE2Ou+9c2gUbqglL2M2q5+HHv4P0yX9Q
+sOsMr2BmtiKWUCqh9A7SlAKRv4awtC5wq3VU4v24GaF67LcMvCz/7HTKw4D
X190bA443ggdwV3+gqAEdItEnhllStfybMnxpyC3AuAwXtU9B5J5N5iDGMdy
bJakwBzuOmb0WMjrL3rq06clPTrtIoYmtLwRqL2p4HAoZ0mx5crSkfVQDHUK
4LlyHrL3y/ADJ6NGiJYjMo+BG0eQM0hYmE7HST0lpXy66mGj68PI8Pyz9F09
76bhM5SixUH6Bfq7h84RGLvYdIZ2l+ChS1s3D3nUJNcKkTcHZKi1/UafIJJM
fbLlxfEnHFcm9TaoMt6q+v69XasYBAn7i5xK/R4i3uV8fnSH1f8xpAUT7Pxd
ekT4OZbarOdPCfDgUYM6QcBdJk2KvaC1uKyNAQB4w8UiNDm+7CdfexFwX0gz
gq0AU6f/dLtFeP8Az+AAjpgtkYMLbSdBVtoWTgaN+CcGGRmgRf96iYkNXpCk
HuBoNcRGNRcAJRY8Nv+pP8GPA1QcsJX4SvRcmS1j28yGUbQoW9JHjknd0dkC
dWIm1kHo9/hZ+4s2Rgwv0u2SYbIw4y2ttNwK/F2ZPgKdMG8M8Il9d8HCP8VX
Bs12dAgCazBOc7gOe1KlqEQgfWkkjk3/g5Fyz6OrcA35oGmSQDLBByzJ0IL+
0348e6u5uH57JwPWFwNEZ0KklwfpkOG9m7UCzuWs3IQID4J8WvHFW17aufMN
fRpmsRwNs/TPeTXeGEEbVV+tppo9faCyVhk8d8oKGdwg3U42HBJQH+XawueR
ffFpUG8aDlNLkGlryYnHwyOa9XbbIJRW0S2fsOTeGQIFHEnSIi0MYukQosSq
g6rHtZ55i2QtgpqNw+MQoaBCQS2hk0Zm6vaZ5rjBfzF64rYtK5OJOpR2dinN
YsJMg8rKBuKFfacId5Gi4Q72zQAd+X/GR9fFCAKPq6ffP8+HrtJ4r5jrSg0r
5bcH8ZiBuj42YDvaJZqq1UBW0LzL5C6yOXeHnToznxF0L0FGeKV539fbt1K8
bnik+ei4ac9hcU+dlEqyJmZ06DaqDofYJiHjkgBXjTd9p7xzB6EQ8bGhNocx
xCt6K4H0dJouxrdwVhm6LxZelYBpGiMad9F6EyuXgDv8Tno2rjYEyc3yxVI9
wZBzU2qnkAOgQhxSY0WpZ7kdPMzrkrLBHYFroWZFr+0MRoaMm0YRqVoZmZ8t
mUU/qCpCkMSc4bm6REZ3T8I0iW8O/vbOB7JC18o5XlgXGr1t/WOo0EZTQkD7
YAE6MKG2+GqyqAsKsm8Zzoo7PRmgdQZE90eq1cqUrgDAmG1DyRXCvIUc4gnC
WcN6twFI7Va/Oy8gjaEljEClgJyXEf2t0KWUnHrr1Bv4/Brzt7hdQSTNQTCf
4OypXQBMPj0YgTZiD9rCUaxEYKW+z/MK1kxmSUM46riSfODaUBgdleMrP37y
fn6MuLIJZKAkYk4Z25g2kTQTgv2tHDdyNF3tGPFUIhE5qNHqCxUuD+5iYsum
QZciwGOW3adhmY3SIB5Dc9t81Ul9BhyEDQpNzWWClJLVuKSxUO/OeWB1P8Wz
T1w1hkRBfD9OF+mzBjXPDQQvknyGdvY2p6aIc8djGQajxDQg5tmde6cds/fd
JW+h9gmP8WRUeCfq0qYpkOzV3GEhssuDiPEq/S7lGEBD/I+45uTsozdXRUzD
9vGvNsmE+K+eabGSXKXN48vJ8henRpQnX97lYQ38W8VePgu5fBiPgNk8WZDs
HJlSo34MwvBopw/GNuZIuLUo4sfRRR80geUv4UxszWR6WEJ/OuWZ7mdEudvy
y/tQD4MwJalfYB8kBJNOSoc1uMATYrmpb12HP0ONornQDqaCCPHc9Rjor/nc
Yb5s+34Vk2+ITAQiFERla6ODG6lFH9DmU1eAOXlge/8OAmnb73l0KL5nFocZ
NzL/pXijRaqO6vqwTlvRsE0ijhYgj9K8A6FxrcnQ+j6JMq95hLPbCQ4KzXAa
50Qzt56+bhhS9CoeTKcEg+ml4OhtnzC7Kx/NpraNbx6MMyKSSXY/gaBPTbp6
6DawpebpKFloJUrzmk9rXXF8NTHU3va22e2ZUeQPtPx3pDwoL4snYUW6nKYi
uRgr2HP4zTyk1eVf0uOqZQGR0joV9nFRPfC4l64vasKxP4swOfY/bBbysvrz
AGx1yUzySWbIZvg1Gky+p8sSCeV4G2Wqli1s6fLazd1WW9Cx97V+WK5jTPxJ
CBLOnyS2y93TWudZ4/OovvDFah1KDyg+C6/YJZQAeLoLJQqTgw4tAVPppaZl
L17jIrUyNEugieEok0IyUMK2k7SNY2bfKp97KY3ust0O92VE999USnHTfJt4
jra67tmIjw05rpxqejodbQb68zb8A7bqdA4/mj7rPzQMWMPHZdwcADZB4286
IXOMKJ4Nr5TGTf4aGmaAsvyybF+j81kY5PaK93yNf1kk37+VIWHsvAMaGRQP
+9aTf4G0VESKNml0XulBeBlcj16Ok4GK7+NgXxFEkkDGrLyF563KNNpMbemv
uXCrQNNp7swUX/I9C7ORyEq2hQVtBG9x8gwSW0An6p2a2hADsff40KS3vf2b
n56tqw2lSae0Ac6XTQxTuBhgIO/sJoNfV039+rfYc1alSDQGX0Jg+d1f1Tt/
DYiGLjfJBofNLDyYlyYfc/KSmy7UgrxkfEEFzN6GxIx8fE2OAJM/5WufeDcS
iu/XeeSnFT2NLi0VsCuMEqRvyai7XoQHm17wdmY8KZxzdRW6hjlghaY5iah/
EDFabvJitATbpbTyHDpVI226N3EipDtRrTTfSrCOmSAtM09iE5qb9uPPi5gK
mmywCwaQ9A6jbocQ+fAzRSy4TkiWsjRR0e9way260DkgQexIbGdLj3+jOn/t
O28zOn/hznjFC+lWkZ7SS79SZszcVRD/K64SmBNssT5er35ZZTvL0uBn7/vJ
r/bBh2RtCojhHCLSROoqshxlst33gcco5ppsSVzPuKWgTdGBjAFoLbLbJh3j
sEOuU2AnJAKcmmHWfB6mSC8PyE84swpKPO3YeUq0B+WtdUjsgVhm7vNHBnPP
vXw+LbmZf56bLzf8sEf8o4mwv/OstALql2TKeztWx3zBVgnfG/QUlX8g/WMI
okhsm7b9dWG2Y76VqbPvSSiGFB7CRoeRakUk0UNrekSTS7p/U/gg6IXu2km4
OYdyd+DJyylx0vul+AGMM8Hu6GuN/bQmDIMQKQs7hlplHrvfehb/whRwXr4g
dsiUc6wMrwL/Zua6d45ZcA99FpExTaNQeqsiPJwtl96AOfulhebAu+/5BVsh
6x1eCNT77Cm8mw5kl2ksrknBNdMT3wdPY38BsyF7ghKnzREJwcPpD1uBN4K4
RjBHFz7vPFp4m5sMD+BBjP3Mr5y2IWQm2V1x1PaFAwGRvb/zPEFZlxpCZ4GE
+6Oqz/aPCUHX0QrxS6pdsVVERSYHYMCVIuRG4dTrT0y0Mx00pBs1/zeNHPj8
DnBghHtzTERaxZaAA8DjpjXXWYBV6CGWWu774uOIinGLA1UvkmRBDLhPQSmX
m81Q0IaunVkuaRr45ZFYkRLOj8bx6eqzJ5KrhTuTox5dIjIJ99gi5YyxHn+C
5Jk2cUvBv185903GYPh0OkRwcYf7UWWwOM5DTagZx/WCbi+TEktxOTaBLd5F
9MYyQOTk6k1+Pn7Uesx1gsfwTPFat09t7uMYxBx0bRl/mk3otPkFub4kTarI
YKzZcZ5kczYfcP60zu9HBxyRp4FnibEQafJXxKUd6ro8T2qDPIVxLf/aDzXd
19UWxpKETbWqqh9GZbn5IEKCFOWDHnZePIVg/mFHVRc3gDjug2AOm3RPxp0/
fOApr6vmFsEj8GPSpadK0DexlnJBCw1eb2WQXdh5GVa55fEu88Aj2jMp5cdz
p+ofjDOmREE3oU+kPSGiMMaKHIOJxmozeD+vcSODWVomVN0YDa20QCceb+zU
XifZuVcDW8ounohbaFAmuvdzEv/nzCYtiP4cGcUYUrhgxGElUMnvTY+5ToA6
vE048qAa+ThUgKcgFkHcg9lZx53gJ8ImUOpe44KzuTnSQz/frcRYL+YtxmPi
gcmxMYLkpoPY0shibLpKnooO4R1gbCpDccfpoQtngtgtQlXxxfbFB1yp3bxF
Cjc1QPBE1vceNQ/tdS31FBeyDJNGRvbT9QFw/30IN+n7oO8MjaXxzoMWsq/o
Xu0/zu+y2tgFQnK4pEReVIcPl/mh2LClUfwlasBPnus14xy2ZD9Pe6gr7w+i
SveG++hAmT44dAOaqNfVvxpDIaRKE+wcfjqL+R6GbIyRdE5cwQ+JATaCHF29
gngiZXkRl1veI3IzhP+sbhePIlFy/hmWljFb9zzGIU3IBJ2DHbg3ZbOwGTa+
8mJtKQk9lzCIfa5fKtkAZFVVa3XaS007debBDPUD1Z3Oun1MV4C1iieNJ+JQ
okdzB336V7/3R5LIvObDPjObSryT6XmPL/+rXZPnRgXiTZKFBZc4CzdZ+QjD
IMS0fBQuo8zHyNE3KSOstrHEELV7F5+oApesIVeSHEARK7HFkNED1Qlh+ifo
CPkaYACSssSSMB+lm5QdPS1kBIpdWtZsux83QxDpJ3vWhFyiPgGouf5Ua+hh
6VrE4Gv/5/CrsNYAjmgxg8Za2togbgjl0oSHeONN0CKTeRdTIt3icnhoPHB9
sDIEEdUe9FUZQ8Pmvo/7YOYb5/9xKqrlqxN7h/gISQDTz6upQXho68FjABvh
Hwyic70ETL1ShtlHtjb0SJ4EMF0fV4B0Lw7JsuMi+nhDhY3HRBCLmb9iDQ08
VIGY8OP4C/YijSJnItO4hB36c1CltPUI06yHRAZVVyK3PWwt9OLbAlNUACjj
tLbkL/Qj9W1+JqXdiUz4mkOuZTCUz2FZokvFivQIoHc3JvT+OJ6aKYk8Zk1W
qPQfRc5oqomZt/fN19rldar+xyPB8XY20Mt3jUAELXbMQ9JOsLnHeGGbK7Iy
1m/yQaK+zenzzyMcfwP0rPMXGr8UZAmggmI+0g5Dxb9ev6LIRrcdyTEIH9L2
vOj4c6Z3bZ0vW00784J7BITFKHXf57ok5XtEK0wcUDrfnh/KBqW2nx71la+p
JqtKQ9+jzHgjpxRnTivelktpwf3BoPHFvm999xVvur71OHHY/fKdA3W6TzrY
rh/5uZnhAk1qIF1TvOv+MO1mROwZENPstghqvurYfBNZlYENnk0/ZouoD+I2
wegd0Za7mW6eL686ypsNUdSlBeBI7ez17F7M7OmIbLGR3sieo6Mg8e59XVWn
tj0o9K0CYDtQjCHyPf2OdgEXm9tbJmaHRrzbXXFv0keSSXA4XdcQLyOZ0Lf+
YpEfhoZUNVUeDUzn2VkzeGmWr9G6+SF50A+KMfpTBg8N7QkAF0v9v0q3zKSX
uEOwNLKUrvnUK9WwxNAJdM5ehMFvRfT8slkI/Wcb+iLMUY/oE2YNAM6vzOMB
x1pujWZhdnSbM3i7IItedkPcokZXlgBdpN2dv0sVqqEWEnmu+AFyqQttjJJK
fz/7RKXCC19ILKBR53L+RVCVUjhsIwU9JCwOYAXsOPezBvbmLmQQvHOaHfLk
aFm49r0v+4ffnlEY9I90pcrVnRMZXx1KUseZ3VoP4Rgfl81+uFlUZCJyU0H7
KV0jfnH/G84AElfcyG318eUuHBEs9sVlKHlJjR4sHHFysGyONHKTUdL2/Qs9
5xvVdIWxacN5AZ5PJ55z9zFWDgh9TRj2ZLVMAKlmZrqtCRT0NUBk8ilo/26F
zpweieBfiwsDHodRmm2FugrUZ7DlSSqSWNA1H+nibslCQ5NKld8mel3CMacq
ybV6amhIr8pr7wcpmlAQZcz6rdR5UHKBiobtL01Uv0cOCCOEN5p6lXQ7fGaG
wiUv52LFQl0MEr4LjI0IaALDDxi/tbaDo2+yfHyP169Synm+GcRRTBZJWb9s
S+EaEOAD/WEqbSA57eWFHgVKOroB8eeKSidN6AJAWWTnh0n+evwGyQK8kDF3
B0OUiHXW8JbJkrIQpbSRVlTRfxQVvBD6R6Bp2wBR8gF3Gtp2w7DD4ADPTQ3N
B8fzjESSLCcbPyqSarQ1uPtgP+fYA3GsTH5UZ/yXoRWDYXZAVhj/xiiWzb7V
rSI3WYz/40QP5HkVkkCrqOKg6XZkYzNn8uls6l4UawvL9LDqs4pJsJEQaygB
5J5fuFMITyOQVC4ZrGphJfxCSaRpgYRzfyf0P0KshpAJW+NoQeYCMp3gwRtw
Gkqdd+W+crterlBVCb60YPfZ0PaERtlDduJhqGlQ8fEC1tw8G0CM1JTW8TSq
nCAdFG6/ZR5j0G4d0DM5x49c+g1ORhsQ1wVljidPTnkmZJdt94DkVpjL5HHk
HaAmecvVtmgYCGvcosXBXnv4LLfbfXJ2QaEjRLhMs5LTtADPndMo4xqFHEBr
YCpu24tWDTkOOMBcqtI+qa7sWUANhg6dSSsrU8xfZIrzE3IyXnSmXT4/A0oC
RU8cqzRHxTNXYUW9t07x9+RWrvOqySTnPvJXQNziUjX3BvQkBx8lbWzxja4B
eQc09KkOBKLhS2gY9Fmyd8wE7ox27VHZokixJ4y3CU3jm+hbYA+9EPUXl9Hv
Suc+27jcvhxp7OHjBhgkspFOLEYgMl0XK661TzAjFJqm/dIjJsPRIjQ3WuT6
X7F+ES4lHmrcaGQ0o5/LW2l813iIRQaZ+dJeksTBwSPKoeeM++SRqUuSClc9
E5T8GklpIbZ3rJ5uphPh5E+Zlab8iHZ43wQyBcy5UOYssLMB3g8z//DVw0FM
yI6s/EEgGbpMIHcd6WWceXB4f5EvjWf4y6Ar0ajmmY4kHY4CUO4Dx7kv+4mR
xlVzHQkQ01QM+LX5Muzgh5tiFlLypthR32JiUWCB+mJ3ZQ3YaZTPcVC0asBu
lspycHgkak+ndbO0LFIuM9qodmhBpPv1MUClVqyAgTEt6zd7GBhr9sLbfIzv
goF01W5nf1LzQy73avjYkOBylcPB4IihZ096VOQcfwJR8uu+GQtNJ//NDQ1u
l85gTH9pZ5UA1O/ngFR9f7vxE1al9z+eFfbB7zRZrhc6+uIql4XqJ1kjSnKt
NPEUOzzXvLBfrF9ucRwaTKkrwLM76mzBKvJcotFD9/Q8mk7GO78/PEUzPMuu
fiaT+3E9yAgZikUnNb6U9KwblKqZ0F3XhSYTM7PqznIDQrD1/okcGVaaykst
skKVZZ8aUa8k9rvf0QwXZmGe6axQchD7UX0LdkCC/cOb3DW5XjsnHV/D9W06
fOTeptEriw/dIdPV23H8NxwcMevhYmN1iitud42J116FGwWVqiR9uYlXF3Np
KD1wAcM/CseQ2VFs7aeN3f5ucO1HRhmYvLzgZx5x0GWcLN05iYUVRoX4dYJm
jpoX5JJXZG9OSnTAIaOrn8uRyJG2MVb+TKC2PJ7llHvwsU/ESGbycJC48GeX
Be35HOIIQOGg+y+Fd/n8/5Vw58UOaiU/O7yZSp9KjPv1znaEOZidgZ3qfuXa
1eaAveKqt33oB05WrCVBzIl9rBoLUKj48Wr+8IZWzar48wZBFG3vdXxaYgh4
QESs+jkjrLPblxnWzSHtBIRHr/NZWwA+8QgfyGEDt7g/C6sBxgx/97ct45tP
nuJTymNIxHiY2dD3RQMz0GhL+fn3i2Z7/Jf9rpd+bvqgjtNr5thdOzp7Pq33
L8e4OCNy9XINAZtcOalDitYuo5zoEzL2MmxP/A8lbEh/E1+xAvF0x63zUaLd
rxeakrOrhbUXu9tDWQsAlNxLBgTwOTs/iVxUDmItjgsgWeC9R4zuEDmXnnzE
J5uNcVu5gCVAFnVs7IfJ6Jpon0LDm7eBl02xzJIBHdYWQdx2kmSGBlVwGXDN
1b0kYQ4kCklTZSg1r6nuQh++PL7f94VeBzipgTps3a87Pm7xVA9/CwZjRBJ1
6Aqqf2PBqXxf+TCehLxqAzB4luaLsjenPf3CQk639g9zciVDVhlw1nBbUGQn
98c9b88HnXunm5rr3a2zEnvuCGwTiGY2wcuqax1yYn3esehZOnDVsJry5b3H
Poxy+YscKVg2kNtHd/FZLMRn9XNmVuwG8xzT7fhBF9TLdM3JtInmYCxOOuKK
H/BK8eBno4yDXPPnWtX9Eahi+YAEPI2jhsQL9y2zGwq8P6n8wZY8eEZ3Q4Xq
A9dswmz9eBIHk9CtrwaidbOpzHLJqOa+ex9ND3LSNvNr+17tIiVYihuOhwqJ
i+u4OrNNunNWSplSTBSh09lq/WCbWvi76IId3FXmpWWcllhTOT0eEXOf0b5T
lL8/JXZDJwwpyL/hab7vw9tiVZONJz/wYb8r2BMAI7WtAC7SFdfeKcwbNFjc
hrgkCQ9A5yuVq678DlCNdSU28xPrugYuoeLB07wLtI30FdcwQvHmCaBl/6lr
hvQ9KgDXWQ7cJ0b7ARqcbHaAUV5zkRISOgtKFv7T5C5UCMNl4ghxc56/buOt
i+XVZrVlBj6lObPwAzUk/VDKB6gdSZ6v0n2qaeHenLSuT/wYD1cXydBqJ54L
JnigdR2mdLlVI2VzYQIVxm9mNK7pIGfiDY/SCvT7Ye/CkmmI75c8KloxFmgD
MSORO8RsTCAw2HWJjUGf8oPCeRU7LoFIzo7WCCXsk3p3DUTNwp3EkNQWmLvf
vwR9F9bE9NCiXgsPOyYKbroUIaNxAKosKoLbNkS5o8FpRk8VY2EHAKZJIlFo
SZx6aUv5bjnGlZfmbeiHj2GUAh7/1JebDUeQwfFTZIFhe4SwpqIJQOKcYXJx
XO5nMfsGVmOL4JQTp/ybMVZniyGatTVggU+ANrzYsX7vWxTt2z/VNSSAcl8S
hfDWThmZVsUy3XEGM0gxmA9AdjYC3PFmgolMux+Cwb8gS4GsJGYcjGpjqHA0
f2Fu1CQBXvw1YSfWOra08C2Zg5d7a19KuV2+veA2XsG6I5CD2ce1YuPwvzZ2
VPvAsBmRqTlEoQI/H0gddN/nkgOy89QhniaGt3/f6FWRVyBxRJeW/a8jlwi9
/AnWzrg5bd3aWJLToagO83Wo6xCcaafic3uCTLO123PVLwRGXGBpW5gR5Ke9
9mY+EF4w+zcfcwLTgwKMN+Sc6a2h7saojyW+aMMlgw+0nHNMrZlK8mvLmkaV
+hCqr+kdEmvR9/elXDoxehNCd5gzOxurGpHRKQUt8s57K7jZZQylvMDzgaP6
ym0v/UFKPqxIBewrvvipT4QRDe2gad6eOSLBVyGsjDD+SesFeGV92vwgJreQ
tIUiqDE0MreVQuFWyvnMVQvtWMp1Ie0KiVL2fUGYtB9uODYFFq1Qq+AvVDYi
s/dTWztjAyU/RpwKgq2srSf3rgEY23e4Qi4sVhdT4Cx0CZqx58nVhKrQDfWQ
qomjD2e5TUiPU740+3ixXDdQoorzR/vbcvUF1IjhEF18++EhF7m6SCd0k+fq
mI176Oz/uDYjbpm24GDx/l5YiR6eR68XsUoXFPLZKXtB+Rr4EEg+0Lv5khF7
8FRpcnDdxWbbdIvTYARFpkewelRR705NM5WPT4gNhk5YlT6/Je2+cRNFYcHy
fvjOeucIUDsJ9rdnA5J34vlZbfiLM70OdqUBiQeAY2T92vFWMUcBR9ALT5W2
PjCpsdY1lPT7ty041X1BcThrjd5kbpiMhN9WHJwX4+WG8QT3xJnFer5bBYST
lVEu0V+CFTWtW6rt8r5Icl6iE5fqSKe4r3he7CzV/VOzMukmrqydOrlk+YCL
gt1dJ6QYYZXlsWPhMdPH0tCIcQW2Gr2ig9HB2KT4MYOy/t13ckCzNnNKx/xg
NWl7jRm9PPqSgkDb1oSZnCquOo8vXfw9fm6RnVziCiOkx1Wi8rxeqPgWU3lX
ur5wsVHJOY6Wp6u0ielXyK0fHbhqWWNcfNPPyvPLBEUuVXLpWZ4cwpV7bkI3
Q5wxT22Y/QgMpYgqv1EqFS/5eVHHfLLnqLVvnNIMocEPVgAVvn6X+23pWaA5
oAI4SjZ7D5OutAd9kWCEGq+SVH8UqrPicpmqkrOB/9NF+62Nz6L//T2/NuYq
mfVZoiDH4h+tFExKZG/F/gEETwjYQM3kCiMTZUbmGlpaCr3fw1g1kQlW2Jqi
asTqH+Vq8ctDvkB6+oTVbAENMimRkpETvXDliKM3fHT1XtHKg6WbBnx90Ipp
HtkgwfvSggskVv+LFLiEL4/j/hqIw4DMK9tmcr4b/qa1EBongm5FCbuCi4aG
YLjOjk3qzpLR7rsFXYBklBSA8VZO0pkqURi4wkPsHPNQZ6ZfeFEyUhDQw2xM
eqLHaQbyc+rN3cYhoUHAHPvLFVvtyS9jbiSX6sES7PGIy+v6EbEw0vyNmhgj
R78fqW/u6wwHCq2/Rn31H4j07Id5J5lsW6FapA16QSLciZZ0C+ghfxqcmTJe
W5ny4lYdlY7Ny3O7dvq1fy8/0q65setyxiUvvQNVtKt080cL3zt8CHpyqpBb
t6uZfnRj9lWZC/0JHwvYjpfbNFj+ETZIEJiJ02CZz7kAQV/2uW9JX8E6z6Nf
elvcX0WnLDlKc7UzL7M7XHLAR5dT53Jtn/7wDTZqo0q/PbcYxfftZ4UgIl5B
SlADRTR7NR1zHGGWykezbvGiRwU9ygSAFaTOzggvQdgATp3kbeEb7RpuE96i
S5BEQ0/qGPSU5qGG9UZHqPTHNnX2ssjf6X9obnYL9mIgaWs1X/rnpnTA6y71
b/XLhnYEjP7pEQBfu2jcSlUBRCTDgURGs9v+5LBuMgknFR71C4yHwfUnpsPE
Jkw5KPA47ozu2M7FlpZPFxYnHhinrTm8daoUqE0rEcYECSSzXRlrkKeCEGsn
c6nnxDc831vXkPYc7t8ijpNuC26s6THYgU0HSOQDld20FSrMxJoiHx8yiw9b
OpbDcLW67W7m4Vxm/pG+F+/R8MxuGiQAg4O4neZetLbkgdokE7f0Ztt/Nlqg
DAmv3q63cJ1OawCtoLTbSJaEWF9CLeZwdhH/1fgE5Xgt2Vd5uHDYC4X6zMi5
lrrkbhHDpp6pn7zdw+Bd2Bd568v718MsHUblH21sS8c88cKgb7CRDl9hunL6
je9EjOrUCh4A7MFTiCRnGr4BKqf2vHpO7x5qFdQglGfT2hiZrbKGvcqRfnAy
zlqUrxVTgXbmdddUkMBDRIIfJusik9L+tkO7hEkEdJcVF7sFgfHraRBLoJRF
iVcOHtXdpawdWyCUapUMXRFmabrQmIjaZ9PWobbCvuTRFEqGZN0m9bakWMqY
U2J633LbuSK1R6/xF42WaJds/xeMDTokgnoVhAX9lBYVHGhb6EoPTG44JfD9
wk/CJEoioMqKU8eTjT+sM2D4uSjVG1O7k0yXf+GHYw9LfUHQrpopd56kIAR0
KrUkn+wcwhTAxiMt9949M1lID9PYhxuoOH9tCCxEbmfNtRfVC8mocHF7TIga
8HrmSPrEficEndWwy2oZM48VK3oryi466/qpcwt08Z3Y+RFRkaBpmHQHLN94
NvMW2Vgpc5EpmTVvlbUrXPac/jlrMsRcnqX9zxI9Hv3LnIEEodYqDHlu/MjI
K4yzUwvz8F2G2Pv3DCgW654FNVy4YRjU5U0QS2L8u7OKVIpbRpAOvJaYA/oL
y9+3Jk/WbtN0eoPAlDSLHAmiNmwmL33JDVmKtsN/64fI7LM2tbTVNfMjv57n
97E7MAc4yYzdA2ew/TBswPIf9en3xmXsWWAlCJfPyGCQK7sbyMOdynEqUorK
6jRuLPifv8ZnB9s81T8MFbFwXtDxjFFf8BupvIfr0LmWfDOF8IEBOP/AvUu7
PLxd4ywvAk8vZGFIZCw5WlhoyOszRgScGRgnf9adcxUilCRoWsMvVw+huWeg
YOIkG/aHwBC6ouBQOW4GLhUGosAHpzRXj2+CCOcAi/MNmWolZBdyEnZnd1Q0
hdq8+FfRsffXunQNVQmAcYRUmeAVEfqaDYDfBa1aCQN2Yr+EN5P3LtG0aJK+
eLbbapGv0XLSYRCIe5MQEwUQk0cwqk4W042JzAc/8sXzlNZf09Nnp7Uimgwu
DYqdehGpKByvxNP+uMs6nzhrVs5u1oc1t0ZhvX0+Fo3Ti2rf+pOsMIxYmNJ4
gnzHX5lj4GtR6SNQj/4ixM9SAvu+Q7oLBsWu2ZtPenC8DyV/xUhDXlgndkNu
uhvoThaS1e0hhxyK0cnlzQCeyYJHK2QfA209/cOzcZEVWDavo7Jj4B6uGTIZ
n/SUy2IE4B9kicOpiEwPrRuE1zPGikEf248nnCfM6jueOnU8/RzCUeH1xkXT
cPDojXqxjaotZRVfx/3gKg2qQm6QKDoPF+EF+bt9WhtlUtnMoKciSZc3J4s6
V/HwWD4tN0vOXSZvU7oQvTVh7+rX2drrBmFlRPd8nVcn+1+iWzLq0Yc6mHFI
9dw/ABeMAqhCYpp9PG2ga4iR+QkHP+fwgtcE31VjMcYXXV2tFXhITr71aif+
fptBym61Mddwp1lQfE93ReQZUFqh/RLLGm+vz9BwS9KdpdSPyKYm5kSzO3s7
mtCL4TEXykK1HSIwhbuwkZDmMbgLw9YUzdfXZd53OrRDOw+zEJMzU8DQJIn/
h/5brFHHtcUvKAxn2NoD9H90L7ky+JGEr8n7YDRFcpgROEb966d/AAfWxle8
uTLDmbWhFBPb1bdzhnWI6RYejVI3DgtE5dbIyMz5LYI8O1DGbQ8o/LOA196p
VpTA/b3YOjsh9ZpDTbGTzhzFfWGdHNI3fY14ksq4nhZdmB8tZZ50ZpLcwC+m
08YUxsezx1VaA/iaJLYtxhAamLvVH1Dd3CDLpDmTQV9CZsPFWq27H1/C89Dp
GJZAdKwvEO0lp0m/hAU4JuulDDdPVBKrkwamH7xvtjkjcXrVyzVYL3E7SaNQ
lGVEkPOSQasfV8oqeAyiPyvsB0/lbUJx1MuvjAakJEEkaTAzBDghFNGF/n7T
smWNT+glD9mqxw8Sd2Y0EKNdPmfXvNK4SjuvZ8oQs2NlzmMwe6frmLbn/2yp
Qrq0jj0S2Aa+yzks1efHqo9WIEcUg/g+QC2r0BMsyGErtuB6XohwD1zl2PDu
iJ+vzJXX7EVRQu6pBwE7yCDOJmNakG1Ip7Eo8zr2JJEHG1T2k8aS6LG6fuSo
oVrEz+Lm6go1azXhDpLSAZ8Mb64k1kFU47aJAYCMubxZZnaHCUUrrH9XjGn/
Vvn5ikb6DUcaNs77RBCOIdiGYyOQ1hDG8nIwRzz6NUNfhmDX8btFwMOlQZkm
wtKFdawKt90u7kIcsA6tIlD103BrvQf1vJbsVFRZqshl2yXz4UJSL3cqA4vS
WUkvhlfZKGN9JoN9Sby/YU8DKvd30VIeQ0/cTjHWze6izdkLYKm8rxozsIZn
29svUQPwz0LYMRFyLVWJ6gynN7w9dGb2T+AWbY0H3X7E8GFnMpWzkC+NcQUD
TfLR1d4RG57y61gXFalZrMWw9ybfwasFxQzXWGXbfpwkMpo35MrcH7ggDMkG
lLaDbb4iwlg0i/aoT4jdYTpz7URuKCFhhBzSQR74QeE7ZnYFQhMB2qvQgeCK
YnWvgtaakAIpdGriWejvhVzQHpBbwHVNcaKLDut9rIF4gqUPskafQsCAQOAE
EtdtsJ1wuf0+OMsgY+3qos/oUMfQn654Cp+g9wTmItrdsdcuBG0nqchnfpek
Jxz28cZOZlszvXT0gW2HCVNmspCZfQ5XbURbNk84bHxur/FIymUBCF9VPrhE
s7KHUxzqUoUgbijPVbVKrl6mVomyls+ocAqLblu0h/JfQJVscMh2/kYEMu1r
uzeWBub2bufGfFZwp5S8tr1LeP99Cj8rb6tuIjYxxUS4mCLc7fqci8xstvLi
fjXuk8N4bksNyRLViIt75mQRMFBzao3GB7Tx4d2RCwNyH6fzAUmnKrmLXkDf
02rMh/if6CMXPzScdsISb/Y0/VsgpqzIND9ndfeZAtqeLViZWNy/2SAjltU8
QkZBYEYYSey9AbDgh9+E7S2Bp8pPvON4K7FQ1LkoE0Z4iLUAPdmzAT9gsBek
Erm3NgQbu7tszHgR8r4E0L8zqoplOhnOJvESqH8hf+I8MD/u6oTdQK6/dXat
/ffaKl9nxYcqVJsbH4znz5/xAORBpUKfUs6WYtx+7f8p+Tp/z+0EeD8sDEqp
4i5kACw2IgpzNgwm9gKxRT/N61LUJNRVddUQScamL+MQe9gDXrHL+bFthZds
TnR1yPj7IQHebex/62c1rPkqizot89YTumUBHKC43YexJggQ3a5rnoVTqOue
A1YEKC37VG46Vvlazb/gcFZjKyvsDr5FRpHOT56UVnIPpa/XGXqxZ+3EsPHd
t3Yk3JfJaiOMklAPYF0tfLqDy1Xt06/GM6ZZ0gYxYIVAtBqGlCpq0d14wF1X
1/oORpirNDSiT0gHIxA/hV9GEslH9PDMKIoiorSuWcCJ9opf1NU7brhLwifl
Pz9qJ6qk+OqybGrGhUFJcmKjLmWW8iTBkEoyQxwYP9XE/LmpUTPxXlXbfMQX
gk+dfvPXi8xloFUkMctAmh02kBW0H0EefEU/idiljpH6Xp2ui7N3rcp5kNOE
DDKUkZEPTJqlrJ5/NR5V/PYMe9DhBSIMb3K1IVqm74UrF7J7X4xr0bxRZvgE
rxJFQqiXRbEsM9e+OTAjH92eEXlPygtmxfBBm325ot5lgfXK6eFbyw6PS2/4
Wf8svl6TB/Sj/UQPeuw36bWJH9Z0qFPc/DiEKZOECBVj2YM1n+FyWC2xdGH9
bazzZSyMvj5OlzZDlFmmc/878Vr1ORnrz2tFM1wxkLA3qKkTBQ2cdaQy+vCy
Pw+8PVmbPJr/HaONtT3fbB735QcXauWRYzGeGxT5p9jQP35Yqadkk7/yM1yw
mtT+L+VrzQQ8iGPFM9g1rr1hLt0FH1oX7V4zCpFUFbpugeslvDAZpxwEHgh4
6BOjgIyK8Z5W9OVk5Q6LDIAg5tye+HPBsU2PQIbg3eyQag6TrMtnFKi692+M
WZaHcX3aqjYaFgC25ICe9T+U5W959qK18CuovqqNegU3dwLlnIbxHc/YS2vY
Vee3Z3jddyEPNE2C1xb0QMG5D4wBtsf+e2PStr/GjLVj2P6xgY95/DePahGd
fZjHKI1XK+lW6nVglxS4ZiLN0v96yCFLfwRclh2YAjJW/EUK6Erq6nHA/3qn
6nSEXk6sWJUPJhjfXyidQe3BbcfVTm58wTY/hvzoP0rb1VeQ/jfgogyDCJml
UoLvYPHF2Xxai2Bd0wCxOWIFd3o2+2+tq1yaNhNDC5RmO8QWEdtSVLyK0jWW
oEKsuZhSwjdgdt6IWTh+QxJIO28CQCgNNO3TgnuAHDPYSNwScUNsU/vflZ2e
vqBtGRgtln3Q3u7OoRT97qVGe/rBOyXjzKCXF33KmIvgmq+zURHwPUaq0O0W
l6LUQgHzGpKlbKvzMrD+lSbnRhmZJ7m6NjS3KmJz3aueJyKJHq5Eet027qj6
niH14OvYQz8lHBR2Ir2Ue0CYiJ6ytFIBv7A4/Szq4zi0XT48dMypAVDS2k57
kSkuCEuCb8ruX3ZMgvJ//oo8czl/qQVacH3+a+X3vvc9bm1aBrf3bCf/d1G2
eZF2QmbbzO/+GOWa7xPICDT1X8gKue+MAgRRuTwdaHb6tab5qDsqEXrWqcCR
kTqr84JZohpCdm0f9tk6g0QA0YSYw9VJrajiQgNzCtAvH4zYHuvQdIW4u70+
AYokDmzV5UjCtbIv3h9mk7BsqfLJrgDssc3h1dmpcmeOa537EGX6kSk0Jyvg
OJ+a3mrgqfAIDi9mXPcI/2bCrYZnF5jhhq9FWrZ2nr+px6I0XGG+6zt01U4m
Lawrct2+kFwkBpXCgSZBlKDdATT1tKR2b6yrDdqo9sQhSRXCVUXuRmeRCBpc
MN7JO7+XgTQ1lL3Vtals4SlKHMOYtpBdWqR1JvHfmZ/JytC2QqxusidscuH3
6rrqeOlHkIlv4lUwUMmHDJhIoDGdTF1JlLs9tqv7UOpS4PMhRaQnpqbATddV
Oybg04UTutp3aWVYiFpr+OlkcztcW9Uri4XZ4fPt8PmoFVvEiPOYErCMgnAO
IdYmg9zaCo0qecMKQh1GztdeWq8HcXG61YFJAYoZKMvNdTOhpcJDPsM/Aoa9
khD/sCB9FlMpM3sUicdnmYo7wYaOZVS2+2r1w5DlnUPc9iABhT4kiZar+QQp
Qxnirv9A+zh/JCFC5E5rsQGRE2ZR4FhRE1amKKcrTHnouPtXraEIfVjC5+7b
hlk/yQvUaaOFD+NKWRPpaMqD8i4fzUCi6cBeagSOJSbDpWo8IBhXeq2Pv5Uw
mjPMydc0u1/48mM/KJHeXdMEnEkpCFCNrJOEq7nxXg2eeBPOwrOdEX9jTAoT
PkrmrRW8XE/3Qi5AwdE5XKtJiLfchckOzIARtVnUr5sjVabDiMeLHN6j3HoR
krpp1D/IiPKgtasSzIwpExQ42AZaX4xlxavlb/RFfQzXp8GAlveslAVTm8Dy
VQbLfF2vwxXgTi8vjM2YZnWjZynx/a31Ym4QiZG8+ONTaMyv/Ko30vKNLGnq
itUBzzusKWYIU1wjUUMTFuhjrfDMz25SMepcbhG9D6btI08YPFfPgA486KR0
7g44072YMASkhgbADCvMAnzLOJ/Hk/woE/j2ZDxYAN3qdjdWFF1QABTkDCn4
9DCJYut/VYi8N5rBjq+CURC+9s26NQH5M+ek59WfS4PV+NrMEQ+ewwJAzseP
gqI8bQEBL71VBu6GklicwBaK5VGyDvm5ei0RYFxCc0wD4fK8dlM5WGUdN+gp
lHN/uZFzHAnHtpByJSIaGg5OeBa4kxlF9sX7Fjkkee2iNGMF+EjJ+KP47iHs
a4/Ljj5OfXNDhvZeGsECAsmbXeInjjVrr8/WQAy65NX/376ZeGDVoAX/qXwb
3DA9P1plsiZnQ7XFf/q/AHzw9mU0HIKH51fB5dbm02TbJwVRnGGeG/lWWwkE
XGqOHne8cMYEm5HO7VBtitiPAiQ3lqtGbwRncRcDRSJzAUaFr7MCwjL7oyRP
X9cZp1PezYGlVeSsfHl58SY9QBHlEKQVQ54djzIyju0xnLILg+7HAoUKLfUo
KDlqUEv4RHNxwMiVV33fPKawbWhKBOub6MselR320suX/tDnwec/oGjQ43ww
yf3/e7t8Ndk7uwPbRCTdoPhuUYzSklcqd4HAIMR0oVkWEDy1ZZy9DGRer4jy
FtpbcXqZM/ZEU6+m/g9Z8NMJcSjUOODHgdy7LqjvUI52bkj48qnVdMEeYOfm
VZLLxSw44CnmBtXbch1ia+iqgJRNLSgE+UFBRfVGAc4yC1kf/063EbW5ykvC
/qr/puCV7uXKo4R2o5JKGY+5ntN1lMDau+3IHL0yD5TWfiZPDGDoCZhKNnHr
z32OTafTvtErHehJsvlt4/kKihng6jpV5L30IdhcSs1JVesNpMrlSlNmYbQ7
AYqgY/u+J+gO1Xci2keXCcsDhdOri/dobRVh5xh3ThaKEFy9EXy6RvsD5yZ7
fkuaAOj1XOFDXNH18RU9GEOyCTtJbVPtdNULs+cK4GqjUpl90vHm3RGy694U
ncftOVDAnx5YTVZBoJ/yj779V92GW2mi1IaXETfNbrkQd1IQdzW9cL6QeGjf
fx9uSfhB3KSo+Rix3akTay/PxiDZq7fbuGqs2XxshiZZafL9EANPfg5sWjl/
gQ3nL6OzwEwrayUhwDZhnclHL+hWgx2PZVF4Ed9gnhrL4pQWfNt7+9Sg9+ec
YfYuv1L1/gYKCDjbdcMtHriugRFSUo5pGOtc3sMizIJKYNr2r8KZOE6IDW70
FnDZzqxELFoeAsfdxtSlhyLk348wTeJRvD9OWR4Z8JSu0kogugCAPYBhttMP
TvpR6iBBxAyZ1hmReGvV+5QFKca5wfEnZSL1mkkIovKoXcWoIAIlBUfGsXZO
FqFiVcja/74pDFo8m+2kyxPmI1biHrju/RX1wrg0QM194ROyNn/Z17kGoq9O
Qqm1OPlifwX4MzS7zA0RgRwwRwwZzRaa6z9BbPqIjvGOgrYGlnGZNa39Sasw
Cp/kIjFCoeRmcBcMtFpgLsM9phgP0QWKKKUSJG559dlpy/7oVsG5b1oB56j7
IKJlLUQZXPsBHCoeJvlKEHoBGtK2Y5+FdusqefKfvvuDrXCARIudxMyTY0Df
U8UsESe94RiHJuyxdUnYdvhedUBhEo25jT9fwoNigVrADwiQzZXS2WUUTyy/
hWi/IPn6GT0BfwBO6Oik5+Pr3AvAQqAsMAN1kyOopl+/mURt1svwv0bfmn5O
J7+GrwfMYdT4m691ZkQ8FQHLxoi3D80CzcENgLWF+SwPSioqtlH23DigsBcm
MtJZCFk57wtVYrJ7hH2Jzmp+388fKnUBTwcU5+F+Te1shLTrJEQ87Py4Ancg
OnoMVilulG60zawy7RQc0R+BcuC8njhP4DjDFGzVw4H/WZ0MHW/Bek3XF4B9
aFNtc8miLBb+eaZ9l6GgNaqs3Uh2dKAQcyCwx3ll0UMovpg5y9JomAGJ/Jua
l8zft45VoFrtVcNmNjkdc9Pzgnggx6UDTY9yLmpRiHJGOUCXqGvLsdsZhBm1
TrAeCGV9vPmKtH5ikAdW/hI5suyEvdWU8XpxiNS/I4ayVzzop6KDjdlStSRH
sUO1QleIKCr903hlo5Rp7KlJy7r8STXWZKdsZ1KI4TkOlE2vmyk+VHH91CSu
mpd7DJEhfMBVhal4vGhO+XYJi8lOQYDnC9EqDqNqLy7QCeEeJyfiTJji4KQa
P9k8shMkHiFnSp7PZO7YI3oyR5+Lm3sFv1pTE7pd8e4voPnvieDUaRdKvyw3
Mhnud/xkqedUQC4Y0SHB+uuDTNbluXiCKAnUjzRV4wzXZfliXCJ4CasMabWp
izsYhlhU2mTkE9aXSNsub6zIjjJxi1oZJFXbSsSXQ6vcfij4z+7jGFokAARm
V6kUiYOHzgOumktoOpYhHjfDDD4vWul5NOX039/tpYM0IP0UjR1F7sxXxC9c
2Snw54f4swsxsvrFfjZg6Mh+39OmJpp6Uk7Ix74NyuIMCRfiDg+RssSQc+36
jsrLnwZHB9zgUWL1PMzcYiaQp1qOU9TyEF3QNAYRKl8W82vboFS1MAvhc1Ih
hefBFB1Uynd3OSBC2+6NlFeSX5AUDJGKW6VxIdJyLMUgI3oUQViCN9DYJTt9
tvnbWXjx+Hm5qFaUo/sUsccjQBWmND5lDxao2YDC+w1YadW/ykscFzYOie1w
vZ9JBUrjvqZl4QhYQImodXHoui4Suiiq/AW8MezngEY3yQvs4pecrKRLdHbt
mO118SAeWAhkPc1yOwRejW4Eo/mnbsyCnilHwr2AYNoZIn45o+4hNf/aZLPO
JvyB8juhv4oYQEFaUSzRHnOA6p9Razp/91QYeRrioCsoJb/6TSC2+Jw2q1K0
ZAZGiMt0qFKLACDYMkb6sAWivNBoJWl031fUq5fUlAYW0wM6M0yCJXnJPAt8
qsCXyo27DaFpr0vUsgPLPT/0WfFFx2wLDEa0/Mea9w8gIDJmiRdjbRbKxiF8
UdCgZVbQGMQhYMrUWeOYQe9KfCNwROdT+fe0sAo0HXf1TdFhn+N/s2eEY+lY
JGkzhzzx4+i2KXBI72lNcUP2GhhSdvu/+1121/goRX+wTrCGeh0z6hd0dJZ+
dM5CJ8C6lqtO9BfzeQc9HWKNLgy70W5N3kbhbj9k2LQ+/nR0OI6NyP1CAwO3
ebDUx4jA/Zxf6JIbhef5N9XHtcHkyT0Qz46XQUZQ7t7xaFmEYJit435zgx5S
/YIQgnvYNJ4DPqKGB8kHqc79/gdVhkX08GHER9ZT5oR5leJ1icjUiIaFXD3/
LJfoCfxIGWlg1Hdw5RVn0p/cPPlvO7Icx3mRK9vqXR0cGBcLUphgkRmhOAss
Q7fcY688KrLN5W3mgGGmt/ScX0LUjSFL/I1SEht1+BXmQOnBY3It7TpYo70u
QL8jRuQIGag5l61OhiWfsD1+8Y/86c7HcIx89MlOmXIFawqmCX1JyKYf+CL9
+O5HPKQDu62iWhD63SS8w+DGx8ZzA8zSUGnb6sD7Qi3X2ORavtB7wDjFWnJl
eyBA7ybhwHdLde212rgJ4MIuEf5AyeEqTdDUiy6LHn7ABF107OcZBHGCIHF9
IgpAU5ak1/jqxnjMVb+me+4/DLW7O2E0jyzjlZsbdXgBDBnQJnlyc48p4WO/
63cwHwA83ZewkD2LFi75/Bqbb09BZw1rZXteElKk1Yp2EFI95bYm/Id33Tw3
69d8AhI4OUl7QXT7IckaEfx9lyrlaoPGky/xnxHrVGQiZWWtxIyrymUS0aFt
GSVPJgSXqYOZaiVggHTirdHsKuCZ9t4Uc6nJCU3AIeaqNlItx4N8SmLL/kRn
KjXNLjyso2bBiKZhxlCX9PA7NNhaNP/yTFXNCr4H39K28xOQAVQqPY7Ssyhe
a7jEmDs0Ft1vpot/N0czvj6rWOY8FxXNRextiN5CYaoVjM6is94d9An/q3GT
sNfwfzLcZahhZ9qtHx84YWnaVx0PAm97sMba+sDIXiUoMz1tUS+lv0BhK56j
Hwl0HxH2xFo3Mg7WrtmOO7T2QVjfJQqSKXspt7JPrp5negloP78wrRZbK2re
WxralxDe2vqe4CSSiVGshorlxM6w2Zs3iQUugpNmwARe4NCqMA72wvR8PrH4
nABtz9qbCPMAE2Fyoc785DvBgQn0W/AQVu+2PWCDitVCQV0G9IfQibTgD6dI
d3iD/fNXvvJGjKGOh5TCZjesAzhdAGIflhEPp8/taB9iefZTBiOXL3AvJaB5
A8R21Wv9WYvhHkJ1ABzl6TILCMIttdFpnoANvv3Lp13pnfFkkNQ5MOlv6GQ2
i4WuiIdpUHWH6v76rqAwYvtIIBCsnA7+yPLpbwcKtXQllBB/gOA2fGzTB74r
aMosAR8gHK0j5l9u5J+B0k1b+/hS2lk8VOtu+9elPG8P83blFNAYD8N8hiqv
y5cX6bCJPGfjFTo4uGvxJD9FowqXTU9SjqAKXDeWGw35b5UoiGztyczyTxVR
KNBeEY74hmh5+uj12R9Pp4R8Z8y8nXgEAELNvMOPQY6KNDrBsikNw52dd2ja
BE8CwETeDdwGYWjbWspjA9pzA8l0AanVRsSNgcx08TGItd/8CHYATWDW0xcx
iDVuOpuOETOWyI0ygKFo8w88LwzroanlKP66s/GPB0QTXsEIw5ixV8CdLIe6
vX4HtBmmzbtKLIG13zpOSqgU8oCnq3dZxulKzw4oyW3zDlKdZaBJr2yloR6w
TM4MZQqSi5bVIUclSbT3gGV4J+/SGoW/rDqh1dSfhvWzznaKo4zbaZvcyNPA
//JK5M6uCDuy+MpRr2zIH8TqcZoWF+bPrmJ/wBvhQVNoi8MInHr4HITPAt58
Vpbb3PmdI1uFZlPGYmVFzlIi5uryDUE6sH3f3yozJgUtqBM5uzAUcb7nXOS5
ivvdnUwVS0TaTMkkRPUYWZA+5zLzhhYmzwzhU0QnET00oGCh9CiAq64Qa12L
x0DBIv5nDdt7TjXKhoIHTF5jhoz4gkPM5L32ADcLDyRvN5w3nZ/gXjwPtQys
X7NTWe/WXE96lWgvB9wrrysWFel/VznD9CjQiBdAsHDmxWvHdapMVKRE9Rof
7c/qG0aFYiBaLnAh9mXIcLWO9VVuRA+kQEBGrXn05GcWO4EDMIR3QX9gMf40
sVU/p76TRvpTlZCiGoH/X7HnaBCNDwn7y7/wqkbC8LR/CvwpP4GJXQQeqHvt
3JSLAd/hq1I87rgQt6WPYyl1Oaj36DV73KrMp4mde2Ev/3i9Y9YDADH4JKij
2hNoiZ9p0jeTdRaxofLkPZanmKBS6iw8qLDzEZ7xLyqz+tml+Iy8l0XO0Sbw
B19JpElIn//CBz04jCOFptqEFYxEhWS+kLQbZj7uTpD5dmomDGVoy4iXQVGp
Bokr0rES9YU6QAKl0p4irHvgQ/I2hGwkeIa9ybTre/ZVy58vfD7CytVrY22F
rXqjTrCxeaWXcwHcqxPjN1J9ilB5Zydn+RqHxVTiBjebL0Z5x07Bi4NHvvFb
4nfJ1VfYCbnvFaE5Gph/Pp9bG+LaltLpYNj8CfG6ZnZ3qjyf3VBAWiEz3Jw3
G8XXq1gaQ7nKHZZRJFiYYFZGZDmWFO78gIG0RF+/CPL8JX708KV+dImbeVW1
DEdq+DxqYQvudoKQ7J8ztrdgyT26p520Fv+rTSclMNOVLFzWeiT7wNVXQh1M
t+vBQVuNvzKnzBXvNc1spwxoiKgSx1tYPn0pESwzRrILyxrDaJj8RTzDk33k
72sVrvUoXCmUuQJljcjJsWJZZCZPOkC0IJ2G0RdBWe9fGG/jm4vuvmnuGZgb
XJBdO8M8wLSuY/l5sHZIZg22qxOaLk3DKNVOyvPmwJv1BuL4scpa5uOCvoK4
TAkCvluI+zLTfo81w8AZ84k8ZFsfYxVp7krkJs1IUyvJymM4xPL68uBeJIO4
2ix9aLp3nHMhm7aMbA/6+o+sJ7mMKpxj7sT6y7AYYF5wu6aSTlBpV2JwwRqn
UxrXUbiTtuslsq/+cc9C4i+kKqTwBIJrUXt9LUocttLAXxGF5wouYgXTeGsz
CiBstZrOXFol1M5XF9V/0GNw31RfzWsp1ODAxxQEV9CR2g7YN3oywcag9/nh
gExk1vGq5/YH8kDlLIzRGGnDxPqJC4FtNjShcabw6Tu+xxJuUsEWMOVhZBf4
TgRGJQx8BlXJa4nd6b9gtfwqA5dOD0xv+v4IVsqq8ntHN7DAMCzoxi/5YAt6
oWgtV15lX+x+fETkKp8CbgM4bt6RHmrCdPqB/3oocRJSH30YLpxJ5yOt99yi
7N1Oi10a3HJ3yMuw237VmduXhgphQsDJlkRCaLKzh9LOCmQ2+tHVPkbNtTVK
jAhp557oZN6qCANfyd94kWGXDAErdoDSJKAtOWUpKuIP/Xy3tT3dXpm/FQwe
jIdJJSFqSEahjL1KE4eng8ZSkmuceIrvo7YNhuz7H1eEYFv2Ik/bRAGBuTau
OwoXAwIHgpmTG55i6kdkBDLjglx9HgqobNkIxA9AKQQZeqUqG7dMeEj68NSJ
Sb/nvtKITXR0Irrzg24G+VMRnc03eHdlKFt1R9Y4MUmdQohdoNoQeOM0u7q0
ESyfvWySQ3WmNsRVOIT72BMEvzViMkRq3Bs3SGY0s53b6CvkB5emY52fbu/F
b1PFby65jjwjmlkdtgyGeWFak3vap9mYug0+bqGDYFT2bt6vwo4QXERzX1AC
HAbssJoxvUfWt6LDm10bB/F2HvBRbLOhnIMYAZdunkuC5Udtz4+bDnrO6IFE
f4ZRngJUvVFFbS0SHK/ONZ7AHL2kTfPdKAfPYD7w+RZOYlYAKfDfDCRh6sCf
0N07m29kQPNpb0Cq2AzdgH4/vTPmcJbyPivIDKSW6GW4E6SKsCaqSgVqawZm
hTJ3d7Ivl0SeShumAkbjvlLACk+Q2tklgH3PTLloUEXiz7fQ9NA1ljKivwcg
j+C12haflmUwyzQf4+u7MyW7NkGeMvMqGwbSi9pvP33rQ+Faue8HNgf4gEYy
Utcw+uqOgE6YCtZmLm9z76L8e+3aCsWiJhyQxckLRpaRpJpafzLQAP2b2jf0
qQG/JGn9frLTa6hObUOAQRpujDdbplDnok2XifC/UssS4SuNI9XXLELABxTz
6aJb0zQ7JvJgtqnSEJrI6Ajvl01D9Cv7g+rjFKB0MBy6Uv4akpdhQXsx1Vld
az4fWRM8GdN34ThSj+DSfcfVwFpWdSsoaGEfI/enQOM6y/wNGVrymhAU52mc
WzIrQXzzWW2W61HvUBSHSOActgQiFj+XLjBnA3KMdNl1UaTkOAioILZ+G5Oe
dLTooeMhryspngM8xpJ5QdrO3Cgsgo2Pl/LDitHivFsq5yWau8AANlOCHrzR
SHR7ueo2bELRcNJfsDHOe7LcVDhS7DQinoqhWmsw3uSZsgBsHjeuPk1Qf7MN
lz0If942C+FoSiLPEcUdsDm9+Umb3dVa3XK4NuQGv43AvFC/76J4hqUsK70o
bnb5u8JsEF5cvo7CdDXspArL0H+Hb45D1BIS1MJtL9sRN2M8hOws3HUgtu87
CjqwzY/VWqNwzDdINCtC16in0scRLbZ40a3mZpX/2qkOzvo0Td2BQtDxmTbq
0wg4VRqJXOpeZiE49WwG25/05XC54+KAwsqPH1BlLLt4PfgPMGDu+85OQjWI
ddiNEYh7qoAZfYmUkFCYaX2b3r/s2LY3VUkhX9zJs0230HY57Sf7HOvK8bIN
T5ct78jI83jFbmQSxsE+oTYZ6ItLsmkCNFp2OYfuS9cdt4u9X4VlGlA3rgyM
88NghCmp1K8QiJiLAr+FumsVu/FltQdjL3cbLzSfhAar8DePoAzhR7pQeQfg
FAcbWC+BvJshlwEDOcsZs/ga1p7rZSu/OP+KXgf/8RbF8ASDfX3sa8h78ecU
jKDeEgKaNhNc3cg/MFIHfRwuDGyikLI+Xk1Z2Z8FyO8K2/tAwmvGvoeo98yL
cazngneFRCvu3epf0hoyt6RTJhg5COCmWI7kWDrdO1MK2EdF0RLbvXHIYkwa
U1RP4lfdaU4JefKe1WjyAH1FWfIj1Uh+5eaqmqQzqYfoLJzWUs4IScv9Nf3F
IzMC1JUjxZQrkqCePty0afEi9Xmmsc2MchMuUvuykMNHOzM+pzoiGk4uZGDP
9TNhFt7jBBIGBAKd//1kUX/iw2FPX9bClFWlfj7G0nR19qt485Rqwd2ABIFe
CaZ4zkLtZuBEyKsH42K7J/SoiemxfPyM/nY95TUxuj32c/Vm9xMLEcZpX5qk
J51qrRLKoiSnfr0hVTDNMdD3D/x3zJDODYh6sUkNxfMPvoDHCbqzFAj2lFni
BnLeUKHb6hedJsjbyofuUkK2nn0/2185xsIpuLAQFAFLMyQzb+w68asXEzNy
OL9do5TTMKik3U13Ms1odz5vLLCwSbnvGVV+djTkDfhZ69ns8TsTars1MmjX
xTZE5Sfra4aubRmJdKGD2C5gct/bF0glQQlCL0YBwSY3PHEIAuIB65Xe3kbf
PtHIi6Weklh3biSSqlrM4ShKCfKBIjh8FxCPzeHPKJttIvZg7O+nGt2qSgwz
8t8D+3gS8GH75X+Pl+7IpXzxLQioSTtqaNjmNc7eimKRXIAWs0d7lut2Ie6E
mHQ+hRN+RBS/HrHeha8GNT7UmK6wn4m+LQ0v2JoAkNa92ctJqUDeJxOEuSWm
4uLsGxVd0tRnG5ZmNQ8Xy3te00tbgAs/L6PR6+N/RMwKygzDpBmwWydPVbV4
H0EX0zG3y15+TzqIkkkYhPsVaV3ZY+EOFpFCvFov8buoC/peWPzIrJ4oBn3/
A36IxVLODLRaGHWx6nJXk56e/hbAVcMZ7oWePMwxQWYvXkAW9J7fc9UVPNUY
L56afOIW4jg5Ee9UhY46MtAMShAKyBwjijP/NdkLIlRBMBSNO3aaNm/icXxx
PTg5avpyGMlnGvPpgPwbZTauXQcivxC6sjXRk/S7GacWIn0N6pXpTlFdniZn
FZdS7O6uX0yNfzK5MchG1Ne1FMQG2Mt6WhxuFrvx98v7BixYz+7hYV7i1q0R
E+rMbi1VTqfH9SXyU3qwtTN4mn5Ia4sPWzdfk5qiLtUuf2t6xLKvs7SXhXUc
AnySAp8SM/FUM58yH0zjnCNjzRla12p84TqLHWlmAORFWmugfTBOuf6MXaNB
pyvswVzIyAxxsV82lgYqpOo4E5BHaKArgYl3Rfbcvb3KdbUnP0xotsYVDyQ4
XR6e1VJqx8Wl85nsi2vXQF3TaABhYIPePu0LKZS81Id9Vljg0KtBsg/7eSVY
C7t5t48EH960SemRlrPuwHPHiqtJILBHM06C7kX5s/1qiJOTzppqgpQjai1x
3eKeYZSBP4RVhe9PKyd0D/F1JcN9NXLaVs3O6wPUK5zlxlKWci173p5HRjgc
Hb4OTcXfm62XOOlS9f2D9q1Op5aKeiiznypUNL+y3AsVBnCn4A52Dfzi6zEl
tYWCOrStVHVAYTRcU0gbJhbcoKFfgCN3FBbw9jRguNmGomILksT7JKtwIE4g
336tg23AqDXwMVSpE8Kaed1+D/GIni7h7w8MZSii73/r/7cjUbBObtnF7bZ+
H5oTp7kntZu4hzEhuxrXG8xUe92QrhF3I6urFATmVnihhC4jq2M10YCkBhpm
5yLNTtjS+SoC7wPLdNI1UNGWlKOMGNqq4ParyFOhBBZj8yIPKoFn57ZDl13j
00/II2gBK7lqgct6B5/DNKkTjIlMtS1rFA/7Bh1Wn0GLnFct8y7oERnCan2f
+T1qCpshgwtt0clnhi2dLfCCCXNSZ20ugkFOwQPyUjtL7eVbLQ/5pEKx1701
MsZlVPcmS189oUoaVHocC7w27HgxW9/g513bRYxnDQWEpz1U7EPDmO/538eG
HPzoHpCIzxXYKfmnyqU3UL90/EkwvDVxWVSbhWQzvC6bsp26BxBepl71GVa3
u+nFaUKBBmkmBdtHM0m9peWMDOR6WhR5oUaeCuz/PF8ARvwNaREgETvQpg8W
O50VqPGuHqUpSsPLAKU2f0Xaq9FYmw48iHsSnDdIqPwUpT4ezo8gu3kQNHN8
ZWpTRZatfgca0N/DfCaklOaPq9Zu43LXff0cQym4PUqV8wBhTyKCh3stWndr
7MRaBSPhcRZ6zuo7YsOl7H3u+LJAtw9y8fxij/j/iIUyt0ZHul9Vspb3DW+4
G7bFQHlFnRL/zQKmvDzxIXS2tY1AEGcdUWKkaDvKAtIwRKHtydpC9sysjqjS
IK6KeJhGeBabIyOeuOk5vJtxFayl7vA4zUa4lOwjKQW48MSLrJ08nFRaa6g2
wZlTfS8VnypyJOgBMNFjNX33yXpCSc7/+ZHecR6HNOu/5wxkG0UE4n8vc/6h
CsJWgj+nNBouAFAmZsXtf2tct7CRTjAIexjI08b5LF0EhQNp7tLiFFUA/SR/
heS+5AdwtJAJr1X8QGJUWIvlhCB6+MhqT8eiRhO4JJW1TsTuxBGePluy3o+U
r/sSUQpDmPOq4fW/USNryJPxlnsdlzjt+MjtnZUr+yKlQxu22/aE4AQ3ccmq
28iQb9ri4JHU9H5UZchP2sTCljXwgbiidqkYTrFl+j6VtoaL6F375UYa/YRv
U1AuW25m93YHYWx54gFRTyAx7i3pgoelVDtZC7502AS63q1icCIIWTXP66o/
319ndk5rwNQ5Qvijy3APOVIJ0XXm3HJzLb/cTsvHstgmznhDGS1CaXgUyDHG
YJnDw2UX+XRSB7jv8jiINUG1DlggjQ1e/6munKiQQnVPXiiApebv1I8zlSOk
SpIPbyMJ+hD8Rf9d4dMk7MBUwgHqet3DWhbMmKyvVPDa1GBTXFn4yxN9OAjs
VDYDWSnUXYotizpsZ4bGCNQxFOsqzJ81oiM9iRrgil5BwclmCIp1u3+ekOis
BZL00tc9ZcEjwlvjf136KTPOP6GFYEwA6iFwANpq4L2KOYd+0m2r1rwZ2PDs
Br2yeuv68q7DtCoi/Wf0HTpJzqKU/bMh+YKcVG8AX86g+32Sh3W+TKtcIA+f
2FA5bLZ5uyCAEjICtB9gjVsTXKiHejo8n306HBukgRwZJsED2KSG9VzkTe6K
bga7hZwuPMHi/p4aJrKhWkpwxluSUumX/a0rxZnlvMPgdUAYhtvl7P2RvS5f
ePdO9awxPKJSEg8WfrsU2T2d0jGDrux5LUCuIiA0hetqeZQ7Y8xWHlJJ9HuR
qEXfjupq5H8GHOV0P0VLubU6X0fWkC35Wy+F/X7buiMZ2yTh7+d4Rg/CDwp5
VGWTP+/b4rX70GmO8y6RYC3353yK0UOP+TxLOGUguiV6PvYPDvsupSKwyHN8
2OMrzvltM9CfiXM9cvtk3qxJrAdG9FyMIKtGa4iQWk1BIGQ534Q98Yiivyah
aGh4/EgSiaRLA8P1IniZvWGeXJ/epKmN8T94e5H6afCi2DSyHbjxECH/kPNm
cPvXMGPjW0ZRvzGKB39XrQoNaJAMCp6Y7V7yqdz0QMNJSYOuX96uXf8Hjql4
aLxx6hsYvMtxc/IoS0x2rcP6JrhompWBf7Qmw4H+/c2ACUSPp9LtqLEOspgZ
tGQ4zY7Se1oKsxDgXOKsNKBqX8cmXpw/ZqNC4IEwjGl7SqQuDW+lvJTHMYym
+gdLypGHs2ij/bidElTJ9Q+4ynDNXHbft7eHqA/9Rn76sC3NlvFKUEJf8mRg
Deh94MQOhxAJh/6mCRDxe84ayUtmKRhOvBh17GYw1iTJeDAmMUHRjnLeoOvX
BrTUpOaRmx/IzGb7vBs9aDst0ZaJBPaWI38aJ/oEFQ7AbYq/m6QO+lcxGabJ
stMrXZ3zWwEzGtdoGqzfZG66LIvwKgnROdgHS7EOwV6PR/lWBTGCgw73/OXk
TFu1e/21MuYq/WZGey3OJxiC/xz9BqBo+D47BnQliWIs4FkfsvtP+s8Ae1zn
GD1KDz1PML8uYo+wGgkjQnRS6PWC6unXrRISUkYW0w34quWo+A/aCEGf0Vv1
ICtz1pyu8riX0PTWEAWyRGnoQYGbBceY/fzEvjL7SE/f2TcEhHIepgFY1Yp6
aqYJZ4lM3wIvLtaJV6BRJ8EjOwhmw0gJE7dJhkOXa7p2EArHIxuWVKieiQAb
Abi4KMt/wKYLCQ2JCDzuElxPXiKADpGz2kp6FDqMWVlI0yE/c58LhixvLHSg
D0QA2L6P6S9bpFSKUUdA3H3PRWqf29iWfMD/PdoCMOgo5aj09TZqzxGbZoYK
u0dFOj/yv6ey37DSBXgZemg9LngCtzS60w9Il0A0VcaK7vNPD8mkHaYmw+Il
AGbMcFp12NoC2Q0JiwcurO+nTYx86l82fpb31lAxjFIXlU58FK7XL41YZr/C
7LWdmcthp3RImzis25mMiNqFWPuV2JSfXGK9eDwCB8O0T1fjtK3/qaTftSlZ
WOLDBJ24uF1RMtTzq3lIuX3BHjC9Hj5LIaMiqck+LoZuMn8BNwfCWP07BIYk
U5t+5KCLd4QJOj74E23dFAqUTThm9kasWwwr5EE7uulLKTjVAhQI2pII2W2/
ix3beZ/ORWpxTyg8EFXnZZWRws3V6aewMtS7+5FgYDkXq+W3brnbfd2VCPBQ
BFguXIfoV79AdP4rjMyUvNxJmqNmE432oG1zJAu6b6NPcpj4EXwcTCkHJB3G
UbvD5Mt5Xbp41zmrDLKw9Av9+cVpqm18ABgmAaUV5aSuSVhJ1rfI584SUmSV
/STq4ucdXBJA0aY4trS1wtcb1/UbWkrQYsCMqiS3OUXB5jKrHMrjU1vcMpgs
fpqmnKvO40h2XhSJ3RLGy93fFxKaZsEIUEnuJFVDLqqWhXFlI6psWbjLgR1B
8kaDwHg9YQRVoU0nrM/BPKX0FQE7x5zDaVHDzCEe9Dur3sXAMGRHADJfkfxu
HpLiMRSbnmg6Jq8QFDFNCPm9kWjMHTfdcKUbNXS2awUbuhWWhpd2vv3asqlq
9mZXrmGVsH9eD+DOFxFsJ9nyPsstJh7aQsauscyM2UJO1GGlp1VNqnVlJ9jS
EETOi8+p9SAVOKOZ0sIFxW6457Wf0xlWFtrWHGkpO6MwdiKoOJFCnefMBOqs
mGMRv6SlMJ5DQiXmkcO6uvog9TmlI9MemQZUe7fCi9raEnxxiGr8tJbDzsYT
V8axH48RFLQSBux/HnNpACG8T8RYbbDQDN7k8hJ5ntoCBcHbega4D0g5CHxo
dQ43yU967lLRWA8djcmZgkQtlydLgfua6RgEzom2ROFXg+yVY7G3EoiKz/34
G5JZMftmkKOw9WtSM+Hy1zUNx96A8DUKqrd3KnWJig7+Qg8KzZ1bFMqKGH+w
4ZTR7RulHKZUOe59uX9FXU/YvXLZcfq922SeiV5iEaCuh9aLDjISRdIaw9m1
JVLXCHGqYAYWRpsrEZjrT1CbQCzA7XKF8lZL9PrkWZm5craKVr4UEBoLKSnW
flAtEUm89hSAMaPBqqf+nCA2BXr5GAO8y60gClvDMqA7QAyLBmDf9Ti//HQ7
ZHIlfuO4cSuuC+BOFzDWWtowFF0bfsvKiWjao/glntRdTkC6G80LuZHt0WKc
ynAQDAbw15h7am2HMw+U4XlmspDiXFPogF5/bZ+lGGVyoX7lFOTXcLaN5guA
b8tAh42RdTBK1w9DV4EcdjIe3cADqlH139Th9GYDs06EXEgUhL8ezHSBVUI3
cnlWcGE3pkuneNnLP4nMko/UuGbawHZO1jyANct77QimNYlEUVx3dpmF9+QR
Zs549z65wUCquy2Woy6TeE21pi9qY4s295oKNWxt/K4mINeQo/0U/dJcIj90
lcBRyAvj8nd+M/jcw+sXeiF03kTDqKoz1Gu8puhcMiOnubvXhewXrtzSZJNL
cxGHnekSKibo2reFsRl+8jVdNZCWO8ron9wsoQmitGCDPY1yLCFSRs23W5sX
eekKumQrRYs/RKWFBsgw1lFvHdPKcmI2BDzL61EQq//oJZC+Fstlcn3OXJ5b
CsqKhMzX5BpXm+8g3hywIryJn4g7NrZ6VaZhYIzjE4IOCcZqDwG2lSy89ydw
BZKKWNUv78VcktNdQO+ZkNMVatI3KGhiBVSpXHbi546CfmftEoZOE3pgoGLy
b3diqL2JL8FKtcWXlfxfiuIVmfmFBorcCQ1xJ9xSJZc+9ScpWX5gNohlmPdj
6Tt5MCAXVZ7DtMmyolGZfs1dqy3iMbomuFoy0OOxoyLpaw6POc91GsLbE8Rx
zpkdhbajDNhpXVBjGaF8EqbQpjNn1TNZMy0UpE0mNgRz5avG6BAU5lZ9Wz4w
8x4GWm2OEIPwVl6KQXa87iAM0L+wQKZvojNSiHcerV4pOALBeWfuZe5DvNER
AXJ4TktQfBCKiCbGHrgCKCGdjzukCM4Vz2EDktSIf2slfW927khAPiSmWSVx
6GxsWNpCcFIyEfAqwY++ykRe2UP94Tpp5/D5YgYVtdb/ayHcW5bGksUQE6rO
nNwAbDw0XuLNeqITDmhHpdAPr8RvC8cIZdGv69ns+1M+EObV/z0YBxPJ/h82
5RnwZMJbcLnlsUPNSYpritVfYdLC76KiiOSf5OTKBJkxgzATcU93aGy6xaSq
pINCYkjl1QDqKCLu1A0VP4OsPuQ25MMzyt9fJvPhet9q7S42WNYTvdz/YcKs
WBn4XSug/5q4wBUsoO6Hsm1SlrKqylWa4MSBxLlzBtf4Q2ChTmafFEjz6qSk
cuXP5gqy5K/yGM0VQEyean9SpVro+JUQSsD7kzPkqQfrSwwVIJplMPPLOEm8
80VS3rQi05IQgcVPNdHVwt8ktlqdoCpj5aQ0tNb438Rz7gKrxgN34vN0EY3F
QjejWTYuQx6FOpSaxCLepYPbizlEbYEEsJR9Qj9vzSJcpiAKQt3jy4CZ4M2e
9poak+b9A3IEHWFWm34cy4Wz7CYpMYLOxE4ssl9tc12n2rVOXZFs9MDvsi/x
OOPRJADGwJbPwjaM++eV7tcHMl904Uh6THuYh07XFz/q4aQciIlUkM2F+o+K
LqzFcA9UnNI+uSp/Wud9QxMXdDV+A7laHdnEPoe60iIK21W/AbRC/MvXu8dJ
hjlZ7s8xmv+jzZ+sqH6KPwvs6G8hU8Utn5KFcqZJ/VjTeyoIgksdMwq8JBFq
a2Cpd8DAEjq5lFDaAQ1UsYDteRKlrR2sLJ8bxWb97xoDZp7kn+WPUZVfkyi2
cyhBLgaCplE5cRkWXj9Fo8SGnYzeh8kxLJO7SBB/G9/VipKlv2wdVbGAimzx
79gOH74IhS6T2LPdBHK543XFDu7rUOHAX9UuAug1vDxQe4oPxhEOJHjsFsFi
e6JcRdX16wAm1ltL1EDgxYEuYR2dT61qYG9YIUPDyN6uYffy6x7WNuLaubW+
ChYb9sb1qbBJZUgz3X3SUzTWJ3PYionneN/Du8UGEjyocpTDLyVxY87o9DvY
EnEMxEWcdFPX8dQM+Ak7dlK6TLD5VFv+1rppd1v8eJJNYesADoS/xwCYwRlJ
hLaZrsh75YRWf+n4UGD3/aZqP94Vgc8+rJYyVmywlxcFIGyV0Fk/RJ12PD68
iLez1WyrcCNPpb1ZaXo1lAQDvbK7cmumZdx24lXLXLeaBrlThQj+ToY5Ii5Y
BmG64gVZl0j3CEY5Ysmiz8gk5oACtrLi5FBV3KwtCPGuueXJgeWqUl8Prt+8
w4KixyTlmc2IyaYdrDJHHoGBFiOXCTg0kNX7LrxJhMORA1x9jt2e8FTJTfQn
NoFrNSfW21SalXWdY3OLd5lmGCEcYr6tLFi7T4isQq4qq4ZNpvOrjA2ETHoW
/pAR6qFQF/rlUYAR5TD8fuyIyhzJaY9NYAybB+t4/R2wyIH1BeK/F6hcafvv
jOQP8wd7QbMDKEZNsNVV1k77tX0g4PsJwOeQmf+xor0mE8kCATxU4FW2imsl
0iISDp4BE52wCWCsQMJUhyCt0imiLKxM6O3thzBYxucRZhCUiutHvzfb5dQ9
+uZuyYYP7kZJKVBM5kRRS6J9iOccF2BqCfCA2qMlPCB1PZigWspjxKER9sf6
DUQBUpqdXr+eu/anAcNrELGdN/PE3stciRNTBuy4k3HW4jsJY6QlQEGcIARc
+YbMinjf4+ItAJ1eo0wfGxVSySlqc7f9N5L6BCMSvRSm4U+Q1wZq/oDXbJAD
2t4w2lIx1GZfkphuk92ddZrrf1HY8joNFw7xzDIgVqzzk4+bKfI5bOskEzmW
WeILmh0cS3o1eMRxQS5JR1Hc+EK/UgaZM9ds0jMSjIsvi5DAHYCZ1rWk34zf
Q6f6wsSVuWEJos75SS1zmXE2QpnarBF+pm5Sh8g+a6XBHRXKzuehivb4SZh6
c45njoDJ2aGLxSlJkOloyZPRauQtteJTYqaQp9nUjfUIVfXoSQEj0OTZvVpZ
qU0Sj6Ag8qww30VOkpRTOseTbzBeUPqRDgVKUmJWbcsLz0h4RB5v7i+Nhzi8
xf2RpCR18OSGLd72Z3zu0fxMOLsMKZsvnyzW5D9FOlPLx1KuAHuxDDh2sN5j
ser+gcrw2RZOSE9zjX5OAYEte9qqYx7wbIGYOyONKlREWMwr4iFMrQtV780a
eyg4ZFmuexF5vH5vmeJ4yztDNl0LpG16WK9kEjY+7tyKO9cnFYpKrWwInJwp
+X+GSG7w/0Y5Qng8H+oo34JrNoo6JAr8wIszeO8GthjzyUC2rWH1DH6i53a9
RVgTpNGXQ6yBB9leqAZIo05WZjuuyxLGmU/G2IJXchpiOngP+gmmK3BMt0iF
DihNXr6wPWKBXy7n4SsEfpcwgK5dOD5fGPZpUjyXeFOPSSXM1O7TwLPxGOrC
mrEJGsaOQ5jjHIUYBaH7RZdOqP4/UF1BiwcbWHYIQfw9R2SDnjNdHmFPLSgU
RPEw0tAzuculj6sHONzY/IXuJe6W14D15g+BqCEpr2LhfgsE6GLSV2SkHOBV
UXMbKwjD5befP9C1Dxq2kKnhb2UQF7Vwpy3/BR3UG2N15OSsXOz4TwmTFTtD
0JxT4vknCwNvsFvux1SbvjuquixWJEbpEfjk/PSoLYTYnVBiZ72Q6qRsKTfb
j08M85vhMc4lSLQi6fCq6rg1qgOt2Dgr+SkL+YMdKFJL2e+liSjRkFBptOmm
5n2F8zNI0bN/lKwPgNS9Yj9tOla1F08qTVoqlAHZTFLi+qgqhAGJH7DaE21Z
EuUlgHffQ8qdw5cj5BII4mgXOoFyAwsznBm1fOB0TY9bvuBcOnWSLak64nqo
02pdKJ3zElv9Ic9ufeuHiW9Unv6Yk0znxwe08LFlT7sBi7SOdFg6HmVYniLK
/UH3NBWHbDZfofNu5E3c9Vb/h0W+5103RUyp4v44h0CfKnsF1UnxqFcAX85Y
MBDilanod6l1XFxQrMnMLsXh+5GQk2bs954ygD3OZhsi/h7p7AxHNN9ZSldX
6SHMHp3gieN/rLWfcQBve6iVk99WAN1m53HXw1ItUvr/FppPwtYlHUt+rusd
ecOug5wplA/2U/kE8fkw/I0a/Ky+lC5uafrzbgKLd2fvSuegLiHFcbc5It3B
TSCSp3kHW2BANPfv1pcLsoGZyj1oQioBjlx/KrZLK5FyTkaJv2Kurv2LCx3X
OoRriDQg0R6K8AyN+7LzuqZRAkIfiNMPZA37Y2Y5JT6l2R8LOSMO1AeuI7nO
gcl6L95e4SkTwVQm8kXz5dKqspKVhSL2M+zr0/mxMFmGagPVadAe30eDU1XQ
m1Iq5hMmyVO+21A5wmzkVIp9y3Hsz0321tk4WiFfYyjc4FD8wBr846ZKQe10
K6RKr2wfl4m/KA7D0okgsdez2DDSpp/BSk0cUD+CCSvSBUM2yNLWjK3wlD7z
/Qu6BFqEpHX1pJnHwunOdVNLagwS2SqUzqEQtncLp6s3vBfjMzRqWZ7KUP05
e/YdJ83dSRzml/68slWV8vnTlsiAVhHvSpIYUmeQPRQyj3hOzqQAbzYwr/E8
10U0KaUeI94LsiN8UVvmCOJzIPV2prErCBdFno+B2VjVr9nMwD5EFLaZTcPZ
NzO2sEZqtEzYEBtcxgL3gFAxIuvQ/MzRRL8GAZq4CFm4SeMkNRydpeboMLJk
2QDbGqEOpQA3q8DJkY803kgQSWqT2Li7wAXSkxqciTr4EX0aNKu5cAURdb12
2ato5Vh8sMa4SsFi+Rqv5TW71G7us4cf8OeN8gb6VDBq23wWh5M2u2tOeZ01
KX+/l9YZm+QqUTieogVOIhlr6z29orLTaQhAV4WN6Q2spf9F/n+p0wwhpbg4
bNUAhHQWPEiuKuUV5AmkfoXk54szUuQxkSygkX+9oWOQskk6fthC6SVlZ528
hMuFIJ8nIHEsRegaPaY2qZeyzCb9moBhhMDBTe1klWaHjbbg+xGpcr6Rp6ys
ZA8/aK4WlTqufZLolj+QxSkxwTOfNa4F7AZk7R9RyyrIVu+4Qnc8xpwKOJfw
wJDbyQBvS3rtaW1h8cBjDTxpBstjrTmAd1rs0TVNw9YQuBB5bWZpEBF2GoEn
S8DisGBOvgR/ZP4xjC/k6gFkTKsWe51fwnSWGosXybeC+vWEuzLsIagkDqek
NDk6PGqC+zurK9uzhuo5XhkfQcGVOlaEIt2+RXK/kDPr73ukEh8uyj6QEpgb
IytrX6uzX9WgmOg2IRKnvZKo+r1jxJKOZr9681SSLgm2KQqSgc9e49m0/CIz
zry2UtXBkGX+dXbJ8j5XPF+DL84FlN//QBDQBJuiCVycqGSD9ixa+3oaQ0hZ
8dfOpn7uHysvwGY9TxwSQvlnGBA32iV7ZIcTYnUDCOk4l/M6quHuLBDPgF2P
4l25RVnUhYrOH5ImSO+SQoM+QTwyA8Q6U+mmpMb2X00D44AIPvHQrvOrjjbS
44UoMs9p605KKTsfr637K8mmMxpmFj9Q7ej9B/owD5eZLLjAxwezv4Z+WrNA
+vUutUDnG9wW+Gn0auayX5LqaFh0fzW80lRxOM74BHRX1P35k2xuFcO7x3i1
R7hLWs/LMtJk6PQqaSspkRn59+AZvcZQiQ1x29xdPHmq6cUNIC283pTJsLJV
6p2YTlX1q9ankjuY+qzVvPqwvS09c725Wbp/TCf4qYA6z/DSYXNENxqvGbgA
PidJwDmTnkK+zXuRtzzy80sWDsmq7DRvN//J29XMopRCw/IKJrbBOgn6xVI3
XvvG+B0T9khmb6XsTNK78xrfxhVdptWfK5H0BlGK7UPeKIBu9zWdQFKhSFZW
z2MjvCSFN3me1PtR/W0mv54Dq4Z1mzTBIxmLgGpL+CFEJyMEKtl/JZfKlw3H
jLLZMnFQ+Kn+43ALsltcXBFiCVxGC1YLHt0jgM3MAiJ+nGptP4ifJqlk7Oi/
S+S83dJsJ+zBHdrGwVL+W5L45w/4BDiqztUFezAwMIuz2gqCMR9kYbtZrOqv
cTtABvPlor4B9prUZvVEglKTDrEXOp0TM9UnO6Ywvw6JbSwfXpjVIK/kW5lz
TkD7u8BveD4KILtEJbWUOVqD03KF4+B2osl4RIPOJyKlYtp/MsuVO3B6DSeg
yygZYH9wEcPa5REc45nGo3QgJ8WG/RyZAU8BuDCSX7GtGaUaNW5VCqeuIwu/
iY704Vdt6rWRmvpQ/nt1sbMIuPbneSuNU+kjqZp/keIj146F3Hi2f+OqoN2z
3WZTHJYl+2W8TaljsWDELpQsWUT/5+aI0PCdbi+J7hjovIQlpAtvbu/UQ4jN
ftRarwDbe4ULLn4Trbz/RGFPGIH4dHmbnWje4GTRybwPiGCjK9BBg296Gb6T
JVhpQugEpGKeMyv6xovPxhFN7o/1/B4AQEoAAMzXdG8yc3DtK79HfOl2ULnn
Jn4l2MPNEqGLoHu9xp2fATHZdAfFUAPQvmqHZvcMkh9SuYtxAcMOBtyLk2vj
oznM66C1Nox1TmcrO3qqpKv0IVsx3uMLxcrWc3DffvglQJsc7eTLRyunbHr9
K3JSU10HZLUroSMNAG3qlZvuqWkK1fULIMzl/du5NY0XaTQ8t1cOehGqgjWV
mUbwF9N5+OZQUaXY8Xu46RsNMO/Kz6sITxcJWGs9lZw8T3bms2u6xvi9egip
23XXwHCDg9cRq+Ausep3hZOsiWEbE74uwOsTtChNu3MTBjOdcysRrwXY6bEZ
H6k9s/V6aOrvyy5QUg8jlIuGkSEiUifsvOpDalWDIfLFL7hkXKJA/qvZMemW
n8/oZZDR5IWeU0rwWZpb2+kc0wDQnRZXeCnlooqjVETPG9utNhqjjwGMBJ9O
ARo+7o4KiU+5I/2ZAfR/QNsRyuG8eGOxiE9l3QykgAYQocGr4ffQJIkHq1FH
zl9CW4CBzdHAPW4ohxeREE2QJOgKjcVbpYL7jAqMLsSPwRskDb95X66mXJan
z+ASmqQLXkyMnNAA2B7oqwwfQhRtT/EXgxZji6ewPYi7IgFn

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q499h2YW8ZOJqGMcR69kpVw/iN/tQvWCewOMIoSse466TjTiYjwzvqQomECEpz+9PbMVw6J4uijLl/njx7p+iWXn1BfQrXo3vI4BtnXdcxGgmjwJnPycuaeTsI4bQM9jxffxfD6wcogo2roLpbxFtr8uRnL4YspchgNBRliuKR1rxWWkQK+nu/v+5iUKQFt4anPMOx9KUZokDt5J3CaWspAwiH0yJV1oSzHLFeCkSObj0Q/gBAcSuLUIBcJtBVjAnCqXS/kNNdvz82VdJiiVzjUGxi5Ko+mYmyHjkAsAxTvXyWC1f9jRh5gJcKhU6XRhrLnpt/NJ5ZQ8Cfe3jhxcU9zUcFLif7FCmz+dlZW23GNhhD6hxY/30N1sAo3a9o2ID1Ox45As/vq5/jQhy415E/ER2F/Wsvy2S0dawXdHnN6Of/KwQUQbjURA8VAU0V52IAkSZMA5MtemD5hltdUInAuHED9zE8VoOzHYlApcw505Lr/HEmlZe1iLQKOW9L7kdojqqA63bQ3gUTqOiiToxCTEZL9iHJguZm8SLHaClkSSYeeT7N7PGjzDVo5+pD/l3LtZNm6tFJWYGPHS5+hnqwo24I1umTfbBBrfNL8plJJq5n7bXbOyzNY6eD32fcTfzui90az48Zu+fam28qIX2ThAU57Vh/m3KQHsUTnflBVVW2/I8aOaxfdv3cGzrxSOMHTsZN95eVTESdi3ldZa0A91UZrKQhIuJAubqaa7KYrWun9HzyMjtqpoORJENNsWw99YvAgei+BLbzjGFuvhg6n"
`endif