//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iOecM+EDYuDV3DVUfX/Ol+qAedui7BdIlsp5j0WbpXNkiabFWcT0Dd6UXNfF
IKhTNpYqzJg7LWOcnXEy0oMqDQZnbDwffKjAYNkYmgnOq+uNVKJSvfy33Znp
JJiOck+TM3WOPEeLb71HpnIYKTyz9cEMEt+eqk2G0chPGzRHesel47fjmZZZ
Qaa+JRfsj7ddt0hT1DxnG7vYrKOBpoMqe8rzoX20+WEC99CeCDtBjXUwjEKI
v4nmwZsBqoDrIj4J3/BkiiS76MbLMk/FF34b4QK2yxCfzezGVF/aOnZr1MDq
fakYjhSFB8Wz9wj5bua1JmURiHqY6JmIzdASS/HoMA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
h/y9qdJSvlQXHkaqS0KqslPwxh9U9H83WZW0VeYpVUdhkYhe/s1orbm01n7o
hZakrwn+eZ3Vu5kcs2AWlLkgKZuAdE+Botp1nRk0PDr3f3u8gXDXLPWwKzDX
z64AqbYQSyQ0IhhPclPSmpptU0nCLNKxyRTfjZZSXYIir7n29fc4GuvsPpjm
F/Xie88EGBsu18zJNKO45LfrjNkwSJgzzs7Eg0oKvCGJVlFKKg7TCsvsO9lk
kw9P+1GV4CRCglJPkfIzn9XHPYslrh1T0mbim41fy/JhgaUQlSbB/5A0q5Q9
vdq+/RozPlKocbFvUs5+nqoZc7jTJdlJi8Q+08ALTQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E3mBKpYeI9r+Llu+H7pXYkGmogqfJk2zCQ8Bu1Hh2H6oC2ZeK6dnkhIu5H1i
lmO7a+cfts9iKJmpYZ8LivGZt+cPY97p4jm68azPmzK5hIrNs+ml7b3ZN27j
w+/n8TmSEbVkZB02ao/yr8TGLZ3TUqfcyPeS60ROozmbC9/pMD8C0QjD+aZ1
OzAXVse33hfpAyjYS9umc3urbuA8xguhv1Ng/W9Q8g0L8GSpEoofguggLMfF
2KyZEckxtaft6CcMLYZdw/lJM/ayanf5l1V1Frn7/jV7hcTP570vm1nkBxMw
R07pBpjnwe6pHHptbnwzSpAIs8sC3eqRSXHSfZdB+w==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fZe1NEIVNm9Ng3GX7mJic+/LxFkggRI3J3TqFc2SnkRUNv+QQzgDuboA/PVz
kkbYrSGk7HsNIP6TN1DJ41oQzalVomEHcDL36+ZU5zI1VwKulGe4M3nvn1q4
HBuIRM7ZYq1F/XLmMZBPdS60IcYNH2/or7rs9fpYbHWeekgSrlU=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ueKsNPandDG0g52DBT7t1cCB6QizktrS+/XOr6ZzPbikdMBHVLJniTG5cBby
76uLcf0SGlISN/JWFnLH6IVtt3fXx5f3RcyF3bulY4gWXKzm473DUZBs0UkD
82+88gePTe/V2VOv3Eh4k8UwVaWz4V1wxPIwwnVEnvJWyNnKp7JyTzSp8eZf
6yGECeC6tmyAyIkGBYzUx4KHTIQ9Td/ykw8qXGl6SPwbvBjO+d4+BZafR8oV
1KQuFZ23Xw8EcASaCwqi+XOKNgPJArKXvD+YGBxD2mD8KnKyhZrdP+0tji8s
Im0O9KzEI3nJghHBPJZG1ETIC95HiqCII9WIA7gNT90ef9j0Aeq/sOIYfBby
BXkMGpneurboN07z9BAvgb/X9zMQJzZmxdQuDAmb40da5lbZ4eQeqG6WIoSW
+5QxoYsOxuvXwm2axPvtPSJ0Ob46Ijc5Ps2XfeG97YejnlUGOp0UeIJ37HCm
C2qKzXpD6Y6lWGbhge+L6CiKxrSnnaT0


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZB1yRWVh5+WrAW0dn008QL+or8KGnnPm/DP4i8pe3ygEVLzOZ9HTazCdkI1g
jZe8j3BnKU3FJ9+MiNuCAaieDc/LcD+2IGl0CqBFi5Go8Jjg4oGUJH7l/vCw
VZmrEpUbJCD3qxyNguzkzdV3gzOOC4EoTGZzq3cyx98IB4bJDWg=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
KLCd6/LIN9JStdWA/mJURzFSYDnrLepC1Zzch6JwS+Iv8JuDaA4A1cB0r6/n
MbEPoZOgRhUWjwbLu2pkkib8WvHS2XJ0ZrYKqTJvTbf2GlpS48yMWpB7BF1L
vOpfV+SiUvYrGjyIu/e0Lq4FOqX81giQPkBD4hPytJNs+6tTEC0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 1376)
`pragma protect data_block
+eH+uo4qlwh3YxR/Rg6HzBBNCLKvnujrvDIKSHeEuI0kC9LF30JUuSWbrl8z
RloS3Tzdh0cK1vinlObtRKS/0MzSpdRzjCWkUsTJSe93IWs4uFDHV7BPDeXv
zpQAYk+k84xNuLYdK3wj3wyQ3qYk6N72JNz+5RSYvI+6Go2BwYWmat1GiFLp
bGSdkGh41dWSFcDzUgzGyChxpzQfjUG4UBdT9k8gMY7pSTHhr4kJu1MjZguA
uxTqBauU8ApalLAIVkMm1cjnK205B3MGiKWn3r8cjo3ZdOoodXRD5SLoV00k
nl7IFNyWnwycP5bC8g76xKqVRPK5gAWuN0uiuO+eGbYCINKIH2RGd5sLWMtU
Fw9brrOm/VKQrq2gNZ/ZEKZDZcfzxMe5R6egP6tpTpHi0cJLUfdqLpnun5eA
4T+0G5fxbWyz/d8oUHH4EsMyx1g3kgTboDteJo+VtXxiP2uWeHcRj69Abw/L
C4cj9bb+IyzLjfFM8MrmsQ4J/v1I1soBTQka8raZ3dA+SyW5B3XBdwQM4dZT
he7ic0DBPv9rZ5y5nVgDzyuxPR22zqMnzgEOyruIt+dDxNatHTwsWTD3MMxC
vWYnwvqijLauFax48dJiqPDtequ8+3gRMnZo+NMi/7CgZTGxR1v3tu3LFcRw
wO8ldyMqNgO23fBPMH4z/ThKZPmXHr+QhtXg+nKbbdL4ajMHzPY4Fw0SH9Tu
mY1vxLukPiqBam2Y6q8Wo4Kj8QLQmy2lYN8vPqqYIjmCt8Fic5/DjtoX+q1T
Fx4E8DPMgqOYsYENI0a7L1bQ/0UMPPnfNmaOKyZBz1hxvC5A9o34at/ym0lq
FWYnYD1cOfxxGLg4u5yGTFzL55+Yp/ZoO3wW8qnVLSd7uxcXnryKwtyvBiXn
/CLIi2mnPhZVJGBsEZQFM+1+eFCHDupBcCq4Hz/HtvTkJGeexuNGM5H7lIgA
yEyYqOQUuS/JRSotgpRGh3QjMuwaWVHyuXvHTog3F9bcGRIGqJT3aqOxX5sJ
ym1dwrFhwN+She9wRgmUbd9s9ZzJPg5xjjsY7vkKHCxrVjHLHeT2dqqFXfCk
FrahcZSiKMI1zcYJhH3L6yAt9hTEE2NE9uzu/qm30QopdQqzoj+hnFCVFBw8
Uxsj9ozAHQg0jaeZanZCtKoZHpsmSYbMWLc8quIKnDftiJ5mVqP7qlWYUK+q
s6cIgl+3HDyB4G9r8p93IRY3+xpko2LEhJjP+UWR2EMI3rS8E9ko1wH3+EfH
AMBdXauBQfugTXR8oG2hwdLEHZljlZ78AY2jZ2b/8MHXqfzCQquchImAAtSn
t2MCfAOeVg7Vey4SpAj9XsVOEWGYHXcIXuvrwYXodfWiFN0chYEIOLJWPUXj
j7O25imQtSxyCnUfToeTdqvp0GEKy8/ZDdXyzeowI8tR48zz82OAZcdhLu8B
m9n1YUq5R+DM6Bz5Blt046KrUBSafCsAzVLwNz/iVewzrzdWIipkExs9uwZU
t+teld5vAvLB/IYVl7rcR39cQi0Qi5tu3ubLo2xnAIdM7MFXjSyOWAbx0yp3
d7ycUiwhKQUujHWF6K7WnrSotQnx+swwD7+wik+NBxBTEjsSdvDL74I1G7L4
dDCLy0WnyLjBupcezA0wKG/haLhC1O4ooHPEY8L8fYcg/kKrIhZEksxN/PxC
62IjWGotVcdFnzMWB94CIEJuOIwLgmrLBZDL3vp8SbmvzgDqbCx92ApnzP8F
VsDo6g2jC823Jb5REmRIqtD1NoI9PZfHybUwijpSW2TQ0tNJWNHynpgNdfNz
WUZ2i5EGsf/EzLDGpNQVVd6n8hihkNydva0=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG0+3Yn/K6IgX5tb5JiGvhSAL0lBnig3qTth0shL5UGiNqXtQu4lFTJDD7D7vh9nDO/3MCOhn4d/8mYq12xNXDM4iC0pzKhuZH8bXicIk4xlLILLM4VX5NcfyK/xo6/+U3+hQmdzuz6szKblWNBU1eiGrdwuI86tsQzrdTVEnBCyD62YglOWCtj32XJWbSSVpJGS89TyuWf07LZI8XnPO9sSUoPgmDL1s5PeU5/TdOniMYYOGzLS1qd0Z5bTHWghbmApTpeeylry2eegTUoFJ81/h326A99RxkIaAAKzPzB3Q2VQAwbHPkpYyhGwfhh2eBr/jLFtWMNk9VxpF+rnrmkUsnk6ee488bFazDNzfHnIKOyvtPVHyBN6G+dpdsd4LFnCR/8Q6JTgBMJSFPY4cEY016y8jeM+x7ov85N/0ru4ImbHTPvqriGjKJGDS0hi0WvFU+CNaUlzP+VNEG9V31SsMjhHSplFB0BUIyhb6x++XkiCWXBDvr7H3JYqGmVBh0MVwr8pMM+4mFm1MZkLZe4Xm14SsNGlxvyhSSqygqINquYGbmUi9xl2KrRn3680lhksf1IRfV07bvXI/aux88oQUEz0n/84Z/tuuDxaLxLY36TGD1OdhO3X5Iq01IIGL88DTvcyXUpUPR53ElQHjerO6re6sN5L3aIVSqDVDJFd0YJdOgVJS1XCAC6reHT95kiydhWZnMO985wscy+4B6GuUCgLdIAiVBj8hoV7eouYtVpLAetqhCoNKydZkSYmGkZp43ktV7sXC2jZZR8MMBsI"
`endif