//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
1CUBNZ2rjQPFJ0qyJT54ShtJTB2tgLRk4+XaDofPBl6tzhq4au5dR50R9A8R
Pfeb3wPmYOC9F7BkThlTztEeGEv8J59j7KLqsmoOeDN4fCsly3pe6qE/8Q9T
WSbfHtc5Nl3qxiMcSku5oQzHcikVMxrr8/pbaBDhlobujqpoqxdYvUdRKiv6
0ANbg7aUbkG0si+10z8sjQHMfb/fCPYL0BmjvlnvmDC3tSTgk7kKOGEiE9OJ
gZKQG0xbWYoM9TFkFL+aQJu2yAdYP2dpqTqYix1iA0bR1p0cJDd6k1wQIyWv
QsjgDIISkOWzlxhZA66pLYwLpF/jiK3kOD+amWGYpw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
bfgjtA624Udbq2/aBL+iMXjGdAsG/xBGEE83nQn+xA4Kt45HvgcJhTGBrOxH
2zzXHxAduOnylc6JDobhuZqUgQg44NnDdzdZ/RtZvroPzqvHiHkgePMtdmVo
89NAlGHUK+aDi1n5NCCk2opTwcza0LlVEgQ5JEwgaaYC+Z9OIvpNtnfR7y+4
+zMxBUS5h4kTaGe5NLWS7R+dJ7NJQSaBdQkRrFVl0yF06I4X+v2q9ieuPQGE
VGpO4Z8wSusmwMCxwXZA9/LN8Z5+yERK2IqFN5xrSwT/hAb1DGLwZaVwkQLH
1jToQK6q5DC9CliFUtuXOqZE3+8s0lRuB2SZwTwJhg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
c0EIsMLMloq4KbWIcQpY68acLc8q7MxBiyzVe6SJLaLFqPLPpTbWyDckgD0I
nmtr5iWWA1VpQCxaWYMrJ0Kz+A8YDO+GhzoerrD3DC3ASYeQS+LD6mhwKZsG
pfHShRfNA7gUzTY1r600SXPnlsw10Z0PRqeHO7lm0QksrNkFMmYmCIXkGMg2
mCZi8MrNeXFzdz4Ba+F7SIuPtQYi9OekUixR/nW1WsAhQUl5kEKRBNhO45F4
end/pT6v/DptXs5fzj2U9oHMYC3MKCfExFgI2W4yYjhdVBcf9BEEqbcYPYaS
jpLhYqbTBKuulAGHWHieE5MdFtb0mFskWzdun0HpOA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
ZjHXF0Z8Tv7ZrTVQHGQplfSZcerJSOXZdEoSUheG6/yeQwJb9thB11VnV4fC
HWnpWR31Id+zjh2LVJt6Rbaf+zRgjtUBcN5/AsKRJZd4CdUdgEq/+/P3AlIj
crb1qh0EG837TGTFdPm9Sm5t1c6LLxx1UZm3m0sldY60jIFD12s=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
qk0dh+bAf9GKjBkx4O2HhP9diz8H58+qJX0t5qGOzTb2UpF1GtInYjjofAw9
mLbul4tkptI61tngO1nHRgozKl8jUEsQWWcC9gjbdSiafi4XBNLvNu6dygOt
oXSFBTP62+wrWQ7jV1zMQltEFKhr7n6GStNJEIS2+W6t8o32GG9DIJ+vhkCF
bl3tsMRRiHGjWcoEvdcDQVJkN9cLwpn3BCGuK7doxROxWuUMCxOckOsbsyDh
wfYmM79Ea2zgEm6l7IX5tjJ3BMIxK6pJiPyWnJlvjOP/sR1SVB+evca7+MFb
uqX3cF/rQjQwvFVH4jwnDQR59aD+3F+Mnk5rNTLpJZDSt47BMThwTjB5AUb2
eeS5ugIW+HwQ4QiXzXIfcz0BBdz7eV3YPwXhdc53Hvslh/YRh9zM9BJyRQVz
FCQEhgL2LyYTdqqJiPCsqCiSLTSaO+q7eQUY2/CFWqB5mdhR5W3UxrrF05U4
wo4Zqt/JzHYvxTzod8bHokU1w/+JWrgr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
b2RS2MZ9Vv3Xl3gw2wDrP+J9ZZ6vM7voR2M7EZfPESx2on1jyxsVewRqxvRd
qAQTHEZZYJWOZvOv6Fe15sSoqIpCWyST6mUoWqwOGTm+C3UsoWXVSFSuAOb+
Oy0VyvZkuQ8VpHaQZuLyLBvUl99oQHPIjPF8JqF8EFTwFlTBc+4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Vsk7yD7TOqF/NXIgfpjan7d1l7aFsWLY3Jm3qm8Dqxn0fkRetvtEL5RqK2re
BmQjJ/13BqNfjJnuYWM8gxHPH6Shu9AIDEkuTaJHyYu3Kzvk2Mc+pUPSqb8g
So8fTqu9r6ojTeUjJSBbcZVNCjLsJdTq3vboKGlspM2JVUJ6FrA=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6624)
`pragma protect data_block
pfbTR6aJKpRvblrA5jLTR92PHF7StiuIwAC9G13JRHXdh7OsR99aODNSk5fC
y6PxI6aoA8gDDULCMCnlql2Sdm5R2Pwys1yLOSGUyUkhVDIouECUkZw9Qr09
WuNMr1IN4HTKfpWc3bpIBJwUmQGwbXeUQVPH48sAN4/uKBvaM+uz9gkrG5T5
b0znsc/s8m3DbfwjFzPTsuOwu4bsMzIHLLdNksE+LvI1oj167IoigdqtqgMc
QXlBZjjM0S83SUyN6JMCl9rYVoi1OEQHKGEZpwWXs7I8N/fgiDELfeeKPoqs
0wWPuSs126ihhkBxftyEu1rbL/ZPigTb4sQXoUJhxk9qxAJ+XVs6Dn0ip/OD
Q6/+Syycuk1Gg6n0CuH80YMza/kBb/uX1MOMBA/bkJ20rm8m45aNubJYNlrQ
QS29ukCw7VIcVEfDM0+s/nGD2zyGrp0lAgnEeno98Z2EwSFgsfKP5OO2qopi
wg7XKbEuukCajWCwFTQ0a2MgLxxapd85FtJXw+s7V1tx4nToSqHBMszIWGwI
Fn+AtSSsgfJi7ymvcMJrn2LyBjJvdSMRTfmCMruYxMDPt6We0AOC5xqp5D0C
YKY8ggEWHNFIh8mkVAQkXVoeWm+9EmUzlZDaPpLMOU7AFRMPPmDMSf/HxzuG
eVcT2vqf8CGV5QCX4C8JbCuJ3h+IYul/4fxrBeRrzA8kB9RXQ3QCpNgX4GLy
u78mPMIHVZ4aasu3mqW0rOUBqCWtAn6LUTiHsGeJaSkDLFPHmVzs77SS2dIx
1Isdwp3g1MdupxUYxzVrWbUKhQzydvFdTqpVRw7t5g/9X399HANxiQ0Igiu6
AE+yVgRPIsAbQdVU1LL6iHpMKQr6Mc4MSzTnOd5tdoET6IlvZMkDbgwlXjkF
sjX0/c+pEA8eRP7W/tf+uTvSMQoBRUnDe9ttn1Xw6el+e+7YkNO36q4IdHHh
y5UsRrVRFTVOViQzzInIj/dVLetg8F+BU4NPlxrDT2jBB61tz178JK8TZNep
eTfupY8e4hbXpqOipPIDMHJUzwO4HedWr6jKLmDJGOytGR30YuVRAWZeIeRH
dtyEZ8SZ3qyqKNA8cxBGeDGNHgAvRSNWqyY9AL2ZjCZxt2yqKfSoucYIGrZ6
bBoO8vOhq4Ei97LI3/1vBEw8eOwC1J7jbfzETdhmbh68xNGgxzNRmKShJ71n
yPBt44tU+dJlyBR658ARmhcSAIS1Xr7HP9BZ1MEbbhCCljrq5sawZ/2IanW/
N29Uu2ejx/rMWhSIFvk/vsdCe0+k8xL066kVpKswj418VJAMbdiA9cNbnS7s
79IcQ6oKYPWMDoAGjyXoA1p+sMuTbnVd4nFU4PAI4FhZDovcPOKpxkg5jT8w
aUiu+pNmW87oRN/5nAdZI3CR5q9SVAYNo980/DtEL7Z1sXuDLIOhZlrPxvKL
gEZYi1mk0Mq/Bc00AYIePbbmyTb/kb36uTCQE8Dqt5ZhiP6P/4ew+ljQCZ5I
ZtRuEWk3jfIXs5MEg9AA+wP4grsA/LYIKqBOzVgz3c/akWpdvx2gUvLXFQHn
VziKLOBd3nYrNSUG2XF431YaqEb8jcjT/DMhc+os6Zu8ukBZUPgnG2mMWKlW
S9MRbFztmm9/RKx4yZ5f3sJJHoAT7FNH/GuvAPLxt2O+ToKHUJcDSuf3jIUw
JrXgakcbng7I5pVkJHi6xEtyVWZ0n/KUbClKIdSUCg9JxML7zFlClsKiSLtq
SgufcZ/MMtAKNfVSO1F8n6cmRlODb8yUMXkI6Te9Ws/yrtSFOYlApE0C6i21
5IAACrTyref1+H6TkK/yYuzlSm9sUAHE1TXMF9I2Vg8n8LLVN+SemfZSb8Y/
iT5T/LjCFf/Zn2E9W2Vak8BjQyq+S5ZteKOMSKeELoPpMxTZgL23HJoeMV+o
wjhh/FY9oLbSzyifVKcdLA5Q800QgNPQevJIbFfS5dxkl9imKmBvwNg0JCDM
4plsd2WJg7Jlm/tvh0H5bAMa+O2omd1N/+MnejCwGMcXZxvwVZ/1Vc9/KAO7
2RjjGAEweuLMpz4hJ2mgd9LsgYzUQyrDGdudUi/zj4USK1jcbHVHZssCnfAX
Vf/HJkUx7Vg8tXxGVV87Z9KHF9co9GKUr8nrogLsSztbTwALE7H7Ark1WYWt
9J172+4oWU+71LfD5U6PdboxPQXKZ2pId/yhsivs0HSiDyjL5CqCl9P2M+ju
cBwoMvM7YhRDk0BuHY9crsF6faRXY+42iKEKjmj+fGZG8qKrDwkwmJB7RAce
fksLd9EENwJ7/LXTPYf/7WxavymEqgGMI30B60tzehnueEDf8+lnofy8qWgy
rgvycx8BEU/TVYtgmQmavzd4RV4ycjIchrkhCCpGSInoPoj5bYgpCqr6C3DI
WKkhBmTRD5eE+PAI7aEaeiADnhntPwQXdX3wUHSdWgFrNfKj9LZBKssf1W9x
/Y6N+q4EFN2WZDfU57U4uRfMjjwNycSCYIZAqdLC746JEjaAq9JY0NFEwzKs
+4cxcKkvuSYpoWRIxwkM3rkvQSoSBJQt7CNuKmivdlZCGTQSYV0cMHk47nWa
LiUU+GMply5mKtnFzMCOgZfbOzyigYBQB0FhzkiZuTvQQM44UIOPBVSoDPyp
1muDFxvO/pJQZNjKG+SMhFLWBlIL9JTQA5VIq8tP0lbx3106g/o7RUCmk2K/
bEiwIJF4AdhasY3nnpmVf46nxduebeBGy1/KlHxqenrlBhaUzzORn+sNn9ru
yazdYy4e2fiCpyGnRvnQPMUChJVM6q4qgSN88qc6WYuvW+COJhB/b1PQWNWm
n5eSRGicIwfAkcKq8lgWXYYhaXuBFXqihg4kJ4j9Spp/KE1hx/hM6vydw0i+
dp+sE1cwAJ9AODiKnA11hS+GXL3Efag+WUXndFGDEseNypTd4kwn/3bHXvE8
bUdd5lCzZ7XXQZBm3oObHKSOPqAvYY9BQI747PKucPCwEmIqpGzQ09pINVh/
O0aiGuwotqy21b5i1tG+3gXyYsu1DLhe3ld6z/S6wkhoeuB46Bh6UwturBWi
hGWtDtep1Q0rou261gGlBBVU96zGXj/icmN4tQktlcPJY7RLSerYxbUoFupb
pQvUbTpRmkIE/kiOwaqL5pix91ln6X45cRXjYA027SBnZ/HhjVA4jSgnk5Rf
SNIf5HJ/gT6i1ALkcMNKLZwVb7bfHw1005IaDMzZZIoy/UMrpb6HlnPx9HaY
YNGmdthX4aR7HqsXjrAsznJWfxm8omwSbqce4iJhfl0d4yV0LjCK0bsBakMo
L0Xwe3xHO3OQmOmg1asGN0HZMN74subHKtYqDj5vlvKD1OgQMtbxmA/ipjB1
3ZWZn0O+gJ2vOTEAUedV86VajGhHQG9I0y0Vc+qinf4OktqCZVU8YdPyxi3D
dhgTW6O8uPoVO/U0sZp6h8IWX9PMvdU3yJEXraLWt2k8cSK++DLIigJt2YVN
ABo/w/6IJ7Qmmv7BFm/LWsywlE307v7JZjIxqYimux9aJLNgkawfbqo3/c0Y
jlzeirLmLA4hla8x4lqTlcacnyW4DYYD6x206FzzmnyVeLamrZZ6JiXpyUTD
5pBeRUvab87hXFgkzFVuLnLVWyl9SX21Fz6QGunRDTP/c1yp4QrBzBQHdYsh
g/TXrNrH2BKwZyolbCMd+FlpoBKMZ7z2weI4J+OUq08OqBBI9sj+xoJLgA47
6agT27VG1JggkUbqqzTEchei8uGqXXKEHXPTEeaB3BF58mG9v4T9mVSp41t6
6pCUCNRWzX1BsHs5sfIX+qR9jxiRiwdh4224iX0hjJ7ORAtWlDZ81R/oSttL
8TpYwY63kzcW/BwGzjh/qDsWBXk0J22LJGxCYD8jtgJJslS/jAFk4UwZHTGu
oscW+/XqvQTqX9rbIslGB7oEDS6j7UENvvKZ56cRkXE0JvDmDghjyv1/IMqL
vxDv9vd6taYCC51kZ6f+pyI2YNdXPp2CCk8RdbFkFBe3Ne0aZynNdCn/5EuP
B0llgaxp5A/hSE3CMo2OKzBmI76/kkan7/qYAQsrUgruS+zUncGwLnTZkz2K
j4D/eAVgZUvHNC0BUStCaDboR9Rwag/z6w5C4oWeUAA4RUzmAqtpMtF1Zny5
XnryLDRCm1CIIgACwYdYtPvK4AYrvbPWfxHZ6iHAkzuwmtCp0Py53a1smxe0
La4IECsblxRp/dXvtRfanyST518lOr2etWLf/xuZGJ3oEXUVFX7VQDk4rGNe
o6MbTMb41WKCtyBHVSzZjz0teyvk61tbPZlylKeOZrd1TcP0UvLPWULzN45P
hwx0Bl9FbSvNcois6LwJjxx/Mqfb1BJR5+zKVl57McLoXLDcvR1tE8wv1in8
q5wzotmK3Z2CS2hA0yqEpHNLJrLWWwPzovjsk/zMMP307FvReZEdQ6l+lXE5
Q/gdLUC0+5QcABoSvYIp5wH0j6BsVQ6D5mtJodSRwnn70UuUbobU7aMv3pQI
FxSfOQauQmdYh10prGjkrKEwz5oZG2Lp2bRI/e7sdi9MVbpeZEJ1VxKB3vjL
ch1M753aW/PUerA+SY7iVLA9awN8W6S0E0SOceAstxpZQc71Y3kNL8H+d6UD
Hk+o8yBrfkeuy02NTJ+uBpDYO0SEBqkJ7RkTR9yfVEcAPe64VVJgnIrC8Wj0
zgVUPjlRaB1JIHloLvgk+OrgTCJGkIi/4VKBwrQNhW1PKYpElhi6XjAeafdh
Lcx6b5d4qK4rfnzV0doCFd7fSvMMirrUy/v3aTiPtOLIvKE58qBX9pKd3ZI8
XU1OhCB3RasYlmlFf7efMElNHcn8Sn5kEunuiUAa5yr1SmFZCLYXnAnJXQ7N
GErvY6mOWRIOnvyu8tm6Gix7fs4635W2wLSF0NUA2PxGnA0IExr3h+TL11XJ
SpUXIJy0Bo1ob5WX3SUj80LwlF7cfIi3V9boBDsAEgMBmkD0p/HXPAu0Qiqh
f61118mbS6tQtD9M9gIevy798MUfd0p0Hg+EOIOCnBo1smKT73NRMWQn0yjQ
re7d8L+/9YxHkpiyArUj2z5zvCvRtS7588HX6azTzU1dxiaNWtUqJszq2vaE
i1cPrpAK5qP1vr5ahE7dbjE5V4KNlxP0X/e9lEKvyiyUQSI7dLRdjJT/WTEC
pL1WyK8TV6qbC9/lsnbWq+VvLFhzlwBBfqvqzEmi4yKvZ6uWQSwo06T4g5dm
bUj0jchWVQr7HDC6M9P9DxDggJ1rrZAK99KD2jFeBkBANK8tDDB7p91vjN4g
0yCn2DrnizJfUI3u/p+BuMGqgXhxBdyDdRdIUhKx42hJMAhmrPvM5LsvQqmt
LwOz46IBXwPhKoRH+TflNV8hB1ZYZXOBPEm1piqByF7Zd3k+7VbARMCz43ZV
Lfc9sRhTo6pEJOUWZdHXvEhJNz0Du5L1LA3dxbm+IaYLZj4E6rTVDGCtpsD7
1Ossl0cKYQPQI31rD6ifhldo0yIuZaPmKpKJkOMo7W/nzkATaKLG5uDJ7Dqv
60T7RKF1F53yO/waKYY0zvdlVGWWUtmZBZkss0Uyan91PMzWQlcJm1W6d8AG
4wDRKg6PXBQ8sEFyAhI2wKqXAbWZyw4iMRckjni5ROcx8Go7hUFVg5lyFJrW
GTEBmEgPC5/F3NWRI00VYwRw1qBqeBdYrbeAxGQrS/MbuT7n0CPBU57hTRHO
HvcXwCW9xgeoQEgwi6jWmpEruaTaO6IagVAOK8qEy8Ap+VV/uLT63G4Vzzyk
h0fxQ5JUa5YQbwcarSk1oDAYjED88JmHdfKx+XW6yKrT+DUxXUMWGMNsjJHG
Ur+BXUzkwj6XOvkQ0bVaRuHkm16J3cs2fRCrQX5gFAcBmo2uFHULjiWweNjj
Tu1TCNnRoxB6MljxTf9U7Rmkat3TpPTxCsaBOl6FVIn2bmNHrV4dXEOevS28
6W0B3L89IacSqPVaC5SPYZ9ZF/xLnZvxqFP4/omtAQe3lr6kNltgsgR9Huzt
O6/mzO16ireKHbXma/10qRa9uWzfuGZF9QOQ7XfM/df6JCtEn8/fZcwIycpN
+zPIairlz3BcUl47Nepdjg7E4SRZZq01z4XCtmuPftzqTaqQpsFDjVF2Bog8
7H4HC07wzp9QEArB7m5yNlVkkBBPc7ImWfTwyzg9E2NtP/7gG3AccK5NhE/s
+gxuxmT+sSTV6kas4FRaTtn1Lu1CxYsWOaalj36isOD8VsS8ARkDnxgouo9d
obBuUj4ma8R7TDfXm/wUXT9m7YwxSdFZGA2dihx78JcA1jPNJf3dRx7e4Ol5
ovkOSMTVn6T5/Geb5U3h5pu1TuaIHmJJjKwceK4y40R6PcmOEP1zwePOA1uo
GXLxqz0QPhGNfMXAbMdsu/li6y9qfVKZY9wc0YyYxzhk7M+wZLDogTsYj1ld
IkzHB9ZyNGFI3pOr9FXM/cx0JLDozaO2qF5vSWFNpztpzi0zoTM06P3T+UDh
fe8gzr7hybChvral68Cl1ElfQQ48oiPF3QmO8gGgUAimTduEy7rhndzvgWhp
OgbrssRT6iAovl0GeYiWN4j81O1dYCANe5E/BQ9UPLJpOSAuf5z+21cYbKBh
v+zIXRsu+RBlx1CnINPl4unnYZKEgvpn2Ncq+YoVh6ZnSlb6tFcvh5W0z/gG
QqFb0jgM862D1jK/KgV2XU/P+ZEjc5uvVtag2iA1OAsif435K0OCZ3Oefs1+
qOuGetJCOh37XYaBSSJd0DSeILgIfIqdpJr9yaZVnRFLmLQRj9/DOJ1M9s7L
IAw8Npvs9R8g9nFl/TkjZYCt9cmh+dx3atx8RqlZKHXeBtI36LGQVj7PIG8L
x/1ZKcRa7++t5sjzq94ZVg3YKSoihLuLBDEaGFQjgJ8RdfoLf5sUbtCkNZUF
TR5awvHFT5PAYEXAK99Ky9hgkAemX8iVTIa20bmFlLiQjSWKHtp3fnecSP1D
m2hmy6oGlQxH9ael/2vOBeNyXaUWaAkErvy/QU9cSWHCCIs/xPccW/1viu18
eXA9C2i3HeEQIdxr/YhYMVgWUu6D9Bi8PJpn6iAB53ajfV64MX98t5Nlqly0
Ol1t/6tyBbBWxgcwsQ+Ax+d7WfyistVO8HtheENj187dQa00tnZ4utFgEogZ
Q7pxhpGcZWE3K7eowoZthWvsaHhDWcPjMRmkx9r7Apq+slz01eNax3I/y6F9
cpDdvSABpSZ1l1nWOiAsjU8NwKT9/ruiDV9zKJy8H7QvGWSw8P7+642FmxO5
yNa3ai4LqTBovdbxvM9w4HI2d/5WDzOG3sdHW3ZEsXGchPygsC6N8QCD4SM4
dhbxVhvBfV+GoT4cpqga34YgCRhj0jYKsykrR2Qsc2T7bf87xdbfoW2sseA9
fhT1MnszlrWE/WrkJS26JuIYfrHg5WBu/xMxYiH1WBKTUh8Yu9i7Yi3Uglvy
+oVDMp/n61ostqa0m0AVpsjlg9q+fQ19Y8NV8GczXeGDxaILRIjyMOkW7mxB
tDidIcbF4okHX8BT+m/nT2yV83y/HVi8KHaKB8wEAIqOHvCQZ+955aJGFsE8
PyuJf34aLwW4eM/eoScIQ3EA79vOi2vOD2Z2G64MXFKVWbsctnPXk95m8+2h
k4eeHQiuolVanG1F/rEB6ApzfoSmojvG4yN2wXiwYOymu1pcWZpGFFKrfXeD
WJ9JZCca6tlaxLfD9hfDuoJiQgzF5RfxiHv39VWz6dQgAaVXdWARB5VPCz4s
x26aJU/V7koXtUvfvKH+xr1tuOL1ae+toXcKSZKuEmmy0z+rS3V+w72aywxG
QV4skhHCgcOK30BRrTg6IG4tyuO/6fCZAtV04A5177owowRUcyQ9M2euWrLZ
Rt4as4w+8CG7Y/zF5X3JVvDtkUoWrJ/uIzTeZ+kNsKyz4IbVl91njBndAheL
prytH0Mq510RAjfZmisfv2mMUcVk/IsyhHkq6IaEM60xzs8uSz+/QpjKmwmg
dNoWWYv0HXFsiR3+FxElrUxe1pgqTZ5GGDXEyVmWU3G9jAogcNaZotMI66io
zANZ23yAY5sVGtW5d8KbAItDijOzAOaukzmCNznTiZni/6rHorvOqQP5+t3+
aRMCrMtiyd1fJ7OeVGqrzBBTZbPEnSs1gbCq8owCrx4/bXju3JuuukmR2zYT
RJZ+e3gbhz/Vv4HW0O7u8+h0faMSynBUld7l4FqAjwkS1E/U/0Ox7o0YL8hG
LitekXAndrgthK/MzUeF375TgOqanUdoZj1VoUJZDvV2U3dDnQ8PT7lg7LDu
XHsLQfLOSiR4YCFiW54d2ynlG3SyBoZOuDKce321b3KybsBMxadvk5CJVhGd
+IXQeZqaL2yTX2nnh+cejvxJu910JsynREMKZGPemZ9NRRUgSJCpu92h8UT4
VIxTmR0gnsQIRnQDOHFv2HLhDG+iXq5Fm3Ncq1oLXz51iE7zTY/S3jg71Zda
fdEfEZqe4yWkGmZEM2cdqH0oUXWCRLk2jiWGlx2No/SD1cvQpefzWUipJ3pS
ZNk5yq0pSOu18oTcsTkP2NOQV4Dmc29GztbGiwWe+VoDiUo+QaNjz6xCUnyE
36jKJ54GcUVRD1YUNlCTH8pMEJIADUyznDxE/9JKW0L3i8hqCxNPvhHJ4gE5
sVnGP82axcuCKJhZFA8yrnIMotRrwBzEKTYZeV6JRZ+NfiW8FqJPWqBL/50V
gSd+EKwuLMNy4Jq2UU6rY0aO93CuSbsEmgWItmdZJdYs22d4MH8JIMhh6ab3
SexYRjqUIHLhiKWsGaKJ12GGMHkSv2vDXtGeUu6gXeiVVKTeS86JwPC+chg6
W5ha3vgu7Lma

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG0DCezUtZVBVMnFzM2Bm3Oi2jKAt1g3JkmVNMGG/5iLeJLqTkbCRDbaixKHCVQ82ZjLU2pJ4Bu1N9vKx2iogLn/hrmUMNEPXvp7One5OvF+QSAA9qF1FkV0S4AU8TFNv/zrqC185kFw0EQehTi13CLQ9CheQeSjZ6eEK+KWA1EA3oggscogC0d2y4wRehdbm9hoWviFqd8dFkjWwIVioemrOQYFNdNiwmyowJg3wrOVyWHdvyuzMTSimqUyJJQDWcWU937ktcUUWgY3feE+PqrCq3NAp0uB4OP/aB9Tmzf4nJgOdjlz4UCEg0LR6fADgNPl0myhgrTt2vbU7lm4yiaIEA/KEhB6swwCbMf0N+BzNHAFufAXGwfOC0v7kxoLVJuSWqeK3/DxtMcautI/xXJFoQxdURXO0qcaBBiTTkS341TfjjfsGQadtXoC6YBU4kOZq4E3kkVSoIBEIo/KNkbn8L/3AZbbUvI9kq41wzY0iigEda8nrqBvMUBIyNEKknDOsDkA0b0Vw8HNK70wqHy/0jERN65hWhb0hMgdEIXUatphSpytOdld4Uwi6tamxGoHvcM7LZKmYJfD8qor7js9VZDYD2riuhrwTrfq5vL6LGLLJlGDpF0uOnYAhkK3GO7f8IYKct8uUugByDUVL9j9QokjoYhvlnlt04eo6yGfy5yXsFGdpq9JzkSnrj0Ye5tWl7xDceTRxCb4jvSbwRWjg3LpsCIh5VHQadT1JCqh1eEpF6PKSB6wXvKQl/5LFJFv7jk/NaZJ7AV3s/PCXMXN"
`endif