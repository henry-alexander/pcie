module resetIP (
		output wire  ninit_done  // ninit_done.reset
	);
endmodule

