//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
uASC9H+1zD5suPAXZ49GOkKnPMe6vqoH3lOrv/8McmQCehIvM70SGhHhsIBH
Wf0hgzU26quWWsfn6W3qRH7tQKEaAjLNPuVK9QqAP7Tb4Y4F5Tr9awB+qYj4
58SqLy6mp64EHobCLcZ79aKtn1jSibzDjvSayFNN95amO2kMJb9nYaem3gFw
lT7favkX9BMjkPZAaKgTTiOKgznm/6QEf6yxHp/mHOP/K4msL4eYMx0uF910
BSOmuure+icavtUCWq/HxN17cFXlZTlOr//IxJI4iVK7AlyaA/BgGbK2f/Ms
1lLJfhPof7WS3lY5OMZ+6wF0AzIRM7AwlUll1h4tLw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
I3ZfJnLLml//rdAx8DKL+xmGXu0BFfhVeYMwzd1iXwmLrFoqIFKAWpmV94Y3
pJGAQ5m0JaYtTYr6CHTNUX8OHmPn7Zp5dCelZ3Htfjiz3YAkXinLQmXPRIjc
H3dgTbh2GSZUh6PZ6+kXFhQIRSRaVmvFJbUN/134MBTshRUqcuyjP7slaAuG
SLOnov7mPjqepPmd9wBi0RqAfKERUMhTXtS+Z1FckVEa8iPWJHNg4HzuZd0D
AfQcV/7Bwg0QRP96KxRpZKFnUSIfA406nHswkg4EM0hjaRnFo8JA5/aWkE8M
L032f1jCYEuadn2WXc8pxV9u3nHBs1Y8nkHOTSLahA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
LUk2nnWrmdk9/lSWH02CtzqWE37h8cuq9V7bud63KPXYMePyMxRnbygz2khc
uNEoZMyCK42F8GV9qNW8h6xV6eVrbR/iUhINVd0mLzKhB3/C2fGNRi8hyIw9
fchGb53j9zdJCJFggx09CGE4zWvSdxetqVdOpZsXCGZBJ31Bp1678inZ/wkw
ZWHku9gaXbGCxgqFp3s6DEFN0Tp6u0UtWR8IhKTQRNVj8dO1CudjRs6iGJnF
9iVclclWaDk6MgsnhVKekFJT60EHw0VuS4rxy9CRcQPmrdsakCU5/pHLbmp3
VepPV2DFFmNxAbZbMESRg9GP/02aBtXMfjKP8ooaXg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oyhoSGl1oEYx3FGy0O4wWP1qVgk4UiJa884yl5NKuBPQW7lIcNevEsp9SyzD
4HThW1HH3egTC2Stishf6xU+NFwwlXoGdWck3MM6D34WpnWFBFj0IgKzksEe
OdcZ18xV+ZP24TkTsn/T9PYEr9fzYf0nxSpfKd7OeCrHwdBk5zo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
ZZZ0gpjgxiyf6QNjJmBOGfbwdyMtdcZzUFJhb2HhdUcA3iTM5ezpE8CIug88
872Da/ahmgjYGLNAPXPsMmnfkP/23PI2V+oUZwDdK8dysDo/UVlAHPZpU0ES
wN/jfNHL9BFjbLuh5wMRwOMzUurg45BXN0M3A8WLPTfjqn6giwdK75NTtnx9
6se7+5L/sFybdcnGSESdT5UC6Lh9+fMhga8A86sO5/jW8nsUgfPBwVdmVbkJ
cv/iyrhaBFmmNszavqiAjMoIRGq8QYb9kKgkIVuhHjSIzED6kkfp4UNyfGdl
rMml/Xc25SXGCXOaj4mVnB1BaeH8VDzQF0Kphj10mdUBdUI9iooYcG1Jsu0v
6/T8XdOfMX/7rG5Dvj1ok+iWSZq8NHYmbReRxKBLnGDFFnlHU72kYCFOLWw1
q0Am30BFndrKjAEOm+TCd9frp9yrpKTlLTKes0uGhTASsyUdr4CoZLzBTtNu
ZxqHJ3NqvT9OM01LOB2nnq6vgIHvonFk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QHJAOlkRjedfK6vkS4jdtXvKIjPyXa0MpZCQp0ZMq5y6TtDiH+z2ghLLfWRu
2oSmtAW018eOIwBKskTs4H+R4HlbBhSyb6LhKpK5G3Ic5AKCdlWUSCpT0cYh
D0/uUytK0Dl2ed15eIOkBR5YK21rNKEN3ZL6JhcvtTd/RrZ90Qc=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
OAJfz5O9r1o/u6uFuEKdEf6P8Qr8hrt8QvWhljNmtIAZwgxFxfinFHPU0Pm0
fadW6mFO4xf4cNOTF6YPX3/ZdftqWn3jxuaJojiPetkq03AtMvnJ0Mdcdw0t
F9764KPVgWiwuu/adZJtYX3AGyxmDMCZCfXWZYI3vmTSTuEOmJU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4912)
`pragma protect data_block
sb0MdF2+XQRTKQc4z3C53kenLUlnC1VwGdnbST7kYsBL4OOoxQWqB+STo5fU
OGnTWidQ7IVgpbIQMTFjxxAO6WAan93P2kGB5RpVdc9DfOd6nOcAY9kaPzcF
YtyQTllhhzFYu7NEjwTmw2l+h9o+pEfwaYK2pe45LQok0f4BvPBF/94U1VZp
L8zhLZivi0DmV5/mqVBR96fq7pmy0GUTuoBNc/BOvnOIJZz68wYcokpHZfWM
+4rpvDGrVVSEqrZEtmv26+mtLiqeJhR3z31BYPK/+POkljycMI02Kuvg8Nmb
yvQEGsBV0K79KmKOkQsFhTzjI4JajvGADmAC/vP/KFnV6P7c/Ua9Q1eRlyur
VPIgSyVpFIz5b8NPvBwDS+PrQ/ewm/iUQaAwO8ktO723ffj2NLY9UQDYRN5p
zeszJ64U9ImgJxcUYNXmD5tOS/xOcucrDdh1xie6mZ2FGQEJwaE/HyNZIpHu
mHX1So4nAQdD5mXMO0SQyBEPsgSMfTqSbVX7FGLwOVR8RLmDMlM8eKff5T2r
nVnhDwTMlc3jkECrgUJpZWO0m1Wbt2MSuBIUpW8bTyyGCWcYxW2MiUZtbLTo
yCJr/ck3GcTrcU//xEa+I16tQ2wZ5KB8RHVbhusHGRcQ3mJu0ZSKyK5EJMkc
WCHEcf9APaROiqG1Ks93I02A7IJZOGbeXvTToz1cmws0kxTnKtaGv3Q0tHta
fpnWA2YqF9n7chxgDnmv4rDodKfGuI85s6Xm6KgscF1Q9Jc0wIwpW9gYa8cV
4tQ+vGUHWV3odPqLBHXSLzP/5PUV6pb177HbJSDlwALSfgBVHojlV4kSgQfI
OFdrIfQJ2uyR4JqSbyESDODo5j0j5WbClOi/BRXpJTGsrzi4VLQs+iiZtJk2
Rj/Jonz+9qCSgy2OB5t8wW6D4nkJxm/SGyxVGPf2/fohn+UKHlHcgmlilWPS
Q+lHdrtXtMjC4HBJbdK0uvhbXv/IKMMbdfF9+ziOaHMKjUYEd9hYIfJR45CF
5idNr33FI4fU3GvlF04fmdbfIiQkAWAI7upHfIMMJn4wXI78x/SRs6Oyu16e
7KYMbHot6x0AnhvAiyGpwzv5f/jKTZH+muB0EeOHJY4tXFuOlTDtqJCx83ct
G/T8NGcftjrxjG0kqrEcqbhNHtHZiWCU/JNhXcAAL0P7oHCoYCbaXwO8iEeh
j6ETUukgP8/wY4JB85NYX2TeHHEspODQOw16PbVs/yNTQzS2VyZ0Un8EgDz6
Pq/vIsPQz2K07Wu3NU6WEjXl9kmKbqDFJ/gE1BtDS1RtdgQRMVsDblHdW+0+
P5aPAkVcsGN6nITeDRVj9sdQato1uPeaWtQsGnIfYq+PTbt2g+cCH1o4s7Dh
Ns4tknWJN0Jmhn/efb+rcrYrQ+ukfi0SqGoAa2hEUlkuC34nj6YZm5LcThR7
Tlre2HoOo+j1QTMUJyOBWF3Vl4XsstEaY6hlMwCV7F5YlO7J8B5JLoPfvus2
n8c48rKKs0YvnnB9p9e8fu1dtKLf2QIfonLBTMefA1FZRw0U9xo1MsT3Yct6
6zoicew3L/FdEm6MllhAk7gOenyb9yUxGpOs54RCYrZokojJKph5s6Al1Cns
2AtmSBcIHd0bLcwisPef1/yUM1yNii2vM/C3iZ/I9lDWkQ+KgID96AM438OB
wGPTf9FdRdb9bIHbx6BKHPPiLN0qtvQ9BtVnEI4dTyhxr5bUuYwQbWr9NOjl
meDEfymR2h7w7HOpyisk/pvqs8c19XiVDGnZ2V5+tfj58sMxI+y1plMGdNjW
XJxBJxvXrKVHc8gpBt19GX99Qaun8rnbHvbJMcC+PEpERgDWBmo7M+803oRw
IfbXpWXvKxqCDpD4te3yap3HN8f4Ev5h5cbgga0othOtkcxteJ86N9dqWwwR
QhLTon2RuRUeYvxPkGK0Gi1TiQY4VfemiKMGzxWhNTYMSVTJ7Zw/Vp1hbieq
Ga3MSQhxorWN0L5wbT7YIzZsOtOspbquLKDgkOe6Zy8ty5doYbtOLeYvCCEl
/+z+q/2nSchVfRb/AsKqjRI1qmXRvv6lrnkT4jFHG55eiB98gqRZb4twyz/g
ax1itdbcvzjrDbjBLfAQDjq9Qh5A8RSfOqnibKcdJztQ/ZCpPvzTAdsXIVOB
Q0mWdFy0zkqLNwyVakK7oHtHDuLZeDMYcJDXSjLtDoFFhrpVHMmVwaA+AvXE
qzcKUq4FiU8kElMtEH8D1rTznp50zVdDC3ObPUz/b7l/dv8rouYYgnJz08o/
5mVZohW+9L8z94z+fYUkrldgu6B+x1znzj+KZcZ6oksXqhLudwMXJSUAYuun
aBEbMYdv27fh8dy7iFV7Oc+iotKL4TS073b8hPY4m3ktcTBcWUfVv1z3RmO3
izYIhcsS9XVrM6wWb4IyO4PjxgFCjIRCvESwUEhVirYRT0SzdJcENF6Awzm/
KkHoCIX6eXg8uwqBYctqgz/1yD/ZE4Uf2aCrdgQ8awZCf6n7I2QmHsRwFQsP
r/te0L5/ZtAPffRz3J+N4KKle8QRPZ6DzxvxrsK6g6n61B+5oQYsyeNG5XJH
KRY+JbFfsVzzKVNXe6J+IjrkB4nyhhMdQFTYCPO5EN0gYMI2W/oPm3ApcvbB
sRP3akqP1K4/4JJUxYsXu2li9mA50EomD7bXKQZqHiyvbbC+yGvCdnLmfVxX
XJRFz44nnV+lA+RwH3KrjeVxr9o6tm36w+pbIZEO9gEHeAtMtENC0M4MEXRm
/VFa4W12e7fxm3BcylQxCq7LCCgJBmaQGVkWgu5yOlZuXc0qqU7VEvF+pWlX
nzwINMAz/xcxmSV3nyQSahAYAlSGG9zII1bRQ0UxJoNR6YzvBVVsgMKLUhKr
gROO5ll3jXXDCdyc+OsfuLtqhc7fZTttoMa7C2yIwjWYb0xVdWuh9vU5RuKT
pFZ10IphvNhHZIeaLKfoMKuauj2wvsdOcGStVQ/lz3VGRNZqzGESRtDeLOn5
s70Somvuli/KtiLDKJUEIL32jQwuyAqErAiWubUxRZhlw6VHrUyKLc+xjSVh
GL5VRG/ois9Nlt3GSMD7vjfBl8sZ2xDsXmALWy68tpLCBegahfk68Dh+vXKz
iJORt6PsEmuEgiqdek99n9RgDQlww6A129ejC/ZyfwC4UQOgC/gVQfDLGP/M
3cn//aqccwroHKd6wCvI09tIrBntbYfT5pytVfhsE27kAlXqiF07xCCMiMzr
CYGBu6IAGQXOe/oNsiQle3fhrUZKnUzaWoknfW1SZrYSwIl252TKSVvlS6h2
6qye+nXFPmf67qv2j11rtWPvaTOWTm8O1f35uez5qEzVk9lx8lIyQle3QZJd
xCIlxb8fi99O/E/9684+9YrRAz+ltrd+W3YyfU79T3LtMC2FqetOP1pL+bRT
itEglffHfg82+wbDojYEyUJ31PML21WmKuiufg+OmJqA+XZWBehf1iTrswqJ
Pddn+wlQAuy2tTEIbp6mjjylO09drqDOR8pH2d93ae9J8eAqfoxFOeMFAdAO
g+vWMnur0aS3wJfvCvOJWcDXGUhu78vSqJcdm8oUle6zKIqZoRI/tKgMxl35
JrC5Yru3LrM7yzLbKJgd89X3vJ/PMxPz47tKkH0rB23O+2+bnvQNm+18UvP5
L5LQEnQumyyD8vP7c4DMtWEoNxwSUrjOOfAxTS8fvgxtON5lJq/txwsNAN20
GhTf71oVy4bzJv1Bu6lDUCtWEj8SUbK0cCnrnsLoW/0hCjCGiJ5q79mTw7cs
MUVNOswtDKTcvjzPmSUW6dVf5hMN2UMtvNLdKPzTCZFNjsXDQSES1Qr0AsvJ
eWKPjWzhllXLCVqn+UYBOLuNSIqkb+3h5TZPYpN5mZ7hDjs0pJV4rrvxx+Xo
mHDAtJWS0nBZZwhl+ZfuBrT8mw9jJ8ckFp4A5Yl6ZW7xwkPc4eA693E7AXqS
/XisrUN2ovEP0m6mlhiBMkBa43krYZ+CvJ3V46iwknVJOgNsFDU0jbU0CuDr
rYTSA4Grn95qk8wsgFn8mdJvD+X2H3k/DnbHFH3dULwtBJaW5eUPIjWrYf/M
bTkHNZIYKGZzcdl5nYuQbQGEtqFhCMcGUq3v/mMrHVjDKQyhqmlykYp6fuzs
7czhHOHIedfdSTdFSaqqAq8LSU+tK097aZ1gaJJchcK3ItUb230oKAbPWQy6
1EL7f46+C6jHHp5kVB5AvAsqvBiev84MsNb8vyH5uLRRvrzF/YCTPVGiD1WR
c4Yg8C4uwCrjTOpDug/N3JiW66+TpaXxcd0Z782hD8b/SF3Q0Uqn0fV4dkUe
ZrouN5Y762NtS+2nOF8tCyxJ+5rLaX37Yfvnm1YAq43tSRukeGDSTksG5Jcy
TRkV58+BRcn5trHjj/4l1YtSB42QMTbjwgC99lmkjHOctILkJsAP1CHzEl18
Iuy4m46qXOn4LCXPqw+7q7jTRtoNW5hTdZNNCd4P4v1YaYOUDnaPVWzQH+oe
rwyOHlDtI5enyZdLuxvch105+7v34HJdvZypHc3Po3WHPRDeSHqqFrCfgBDz
wM/cncurX/YqB/WLvjbZs543/1PsUpk0iTqOy5Mrpurnd2wvVTFeRvDCRllO
NHjb8yH84uKQdPKtTmkTm2ZV5eQn0+RequHxvpSyutN0iB9I+kNaTHLmhbQt
nHcGK0VIVMcbV5RqbTLe30KLrxotgYyb5IswzY7TN7DQFLg3ZzxSC+60qlL2
Z/2sPg04PNclm/+oM+REDNEst/TDQDRyrJVQFWJDOwbbkjeeSBn4GrXxIs7L
OByBjrOFP2yn5Wn2tkOJvAFDAqNe6J3pY+HT8K3q+rKeoL6QZunR0WSR+L66
GxAmL/75hf6XAynkpVzh1/eHPTf2L0N3Vacfg4ZD3EDoPM2+8MHZXXPmHO9m
I57lGBXDIgkqrh3HKvTTjQb5wIOxOmHrYCruuHLkDQpX9qNzYs07TWjKVYM+
xrKItLgue+aLRX68C3K0ru9qGyb8Oj2BbbKXWrmJYoosD5K7VdfBquUqxY4i
RV8FvgvEJ2p7lV26+pIr95yYYD2W4f2IQfbLrSElKquj0NtU9P7C6+vREmA1
3oyCtg5wLddoM+aiXj8nzK6+Rsb99KsSty3VzYrgwnmLQntfVFAoHwI2R92r
rlf255dtOdsMR7mirqj2QiaaVmtz5wp1aA7IXqXz7XsQo8GOXjCoGw07dBEq
Mc6zx/gN/vklEVX0qyQODjUZEavEr3SletagrY9FlDX3b100UP6vfTtJJhfd
aA90pzTpONRQ+rBB2rvx/BPZBvuYPszQzalXdTI95XqKz/bcZ7uJwjAVWVK4
xBO3u/N5nZvTZxjpAoKYrP+nIpuB8nxd9SIiSUTVGX1HxGSRVHAJATA1SzQG
UfdUo0O7TIO3y1jcOxTZEfGE4bE66ge1F2LAdNMNSaJWdJydUlK2nDi/npyk
Wq4mei6by9jNYQ/Zr32uqxbcGBSgVXjNXPDZiCJs9nNhpx6nNNOocz1iJKdf
E7EynsTBZgJnZYX9ACe1TZ+YWlmjo71NxxraWf1G+gSmapl/uC7aR6N4r4EH
WqRax7fBynXm+oSMOEqJ/WLquDXEZVGtNQTuTvNjt4TKDcOJ3CebOvGVXvcn
H4ouDVGfofhT/2dh/mQrCGIOkIdp0Il4zLokGnAJ1/nZZS6xXszcD1Zq6AUA
kia9Wvy/6CZE+i00+qW33/XjnFwy+1wRE37OBVwWaqov9Xl0VQC2zOa0IwK7
jfaqPtzyvZQS/SQVNoeYuR+SLIP1QPfkp/OzcLliwdseOLhVl9UKZ1mfA+Cy
QemulH/5vcgYPKR6010Dts2AQro7MpO6CxOIDi97JYaS9Ui6UERzrr0HvyJs
XtoB7hmv57emnrUnQN0Tr+r1/IaWKYgSTxRyzaw9jr4VV125MH4hqqIpbb54
iY3P7J7IyIPgmdUawOB2GyESZAHF0SfcFq8SWFmtLcNFqJzlXOVDv2gib4lq
KwJCdC6c/aWIwTPOUKHSlCJAJr/0hx/og02mtxm5gKtwTP6bqCnAB9sD8BaL
y8pPcRsnRqMx2fn/jKTIktqwMM6Lvf3Sa8QzDG220ihv6YbQSOTOQsrLWmfq
GwF65pdiZLnUcoV6mhZxj+iCx+tWzjAGxbCeYu35dKsdfiirVtWwmbIz9X2E
AmvThE9t7nwFWdT84PBhIqWsN4MzWEl5DrOvfLXjTpX4NDCpHy1GQAGZFnYm
3zR3NnxC7Vum3aJZc3+Y50krWDZsNwk2j0no1IYC9PS2pzcUguyO6Lx1HMwb
7Q7RgpBuKocmjkWxW4YRlgibu8pYraicLav9Bu2wXCKjEmV7K0T8uWnOss29
/jLHgrpA3zNSUxtT5jojnorfw82KjJ+uLrfACyjqLx/6fufswTQtmbNK7GvL
BPbLkqbfX95q2yZaSA0MW0ONq/8n2ykT+jfafdkJASOWftnxjNzx00I5SmWg
8SXVz00uSIgNBm+Ua4BkZcV2aXIfZ03Lf3lIMbtp7llF3N5eUogt6i+0A9q5
4UKjegZbIg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+noeinZwey8qi1kdaEoVa6tn26vnqg8t1gymUoAW9jQYBtgRk4S4vqgS0WwxnEM6NwhQwA6httClffHbewYDHbAJlXajJK9m/iTyHDf8Ptkc7FfQj82VZrxuWjxtSiuJKUPOmAvIQT2yjIqKZz844alvDBeaOM/FNEsdM5TgCJQUfKpmJfGF9cEJWzpNd7jzvkW0/w9pANiZ8cmvgzx21KHNjl0EdM61qEqM1If6Cp5IIMQwC+TJLQJ9m3Gmt1ZCboXnHo5PrNRnR+kGL3SiLznh1ehkSBOdemM3moIom+y26RMHMBn8jhv5GkjDERujoU11gu9dKTw0uMtbdQa0hywkx5iSEaL08fW3GWOQZE2xK7OjPh6IOSRvNjRxie13PdEcmnc+5Dru8YFeJxciZkWyrASaPjUffoKl2m+6mhJPt8iMpddd1pFEFURgnrg5HJqUoO7k4kZB6tnOV3HeU8GerPJt7w1QV/CA9U7J8bj5DsKOzQNY2XAXdgwH8rNNgxNHwxVgTRH24glQeOsm1BYkRYE6shil3tvESg15XH4zqjyRiBkOLkEfL0HcLxY04V+8qOLwHcnNBzHPFQ1vUty1Yb9zwW/KYWO5hkuW+yiTPpPd228aRx1Rt0qfqlpEN9tXwDJtXtlQCkqyRaFBN5b+RmdJegYOHMgOu2Z4QYCIgHL21sGnKS5XEk52NoGVFD6YD/ZhWpGUOyH1g2OpvkHtlFgqbV/pNsqvfMrg5NXHrwJ2gQkSYbpSOCQmL13tgTLBnfamlRVtSDYDXhMwecZ"
`endif