//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fMYSU5xBU2gr1jJ7IOdCCSq/vygy9McdCr2EVC1+EA6Ri6oZVv2JXBC6vPKl
s9A1q/JRx79b3bIwl5t8DJwFmKv+HT+TQXn8ppEnVnWq2J+DLgIBw/5tfAQ5
lVls5VkiqJOF5yI2Acj1cFdB2bOPLhNsCRzQN8TPb3dQk64wIKDpJ3dNqJMH
H9cSeFO/7Q9vAuhyQ9vySNT5Pb3Tl2sRcz7o8XH8Wq8ZhwuSFjr9QrZ1HFv+
F2jHYQ6F4CIpB0XtHgyUcAxcV2IEAazGgqHYGeXh7APH6SosyF2xOx3cqyvC
I20sJGt0ZkU7f0zl3rXIfGqdanZpfbDz9nO+RYoRKw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XqxapMo4CdPSrLvrFL7J62+KR3Vcz8gELZ91xfnaPH5v0yVRU+NcAe5/lBLD
b+CM3YldVipM7TKKcQ4Klf5g5RNfKEMPb7imlGnwNFwR2CRWSbK6mqgYT8QP
cTS5r5Dt2EhNuEZYzWhyge1sGC3lOhNVS8hiOQDlROmlRTJOnb3RGro7n7vh
TdlxsMSz/TabWvWLY9MMDXH79hXf05EGonpySPUuPrXq7h36ItWcW3T/Z8sp
aDJrB3sxcdDxBzBmD0eb3hGf3RuB3JnRz+Ufzoi/RKTwBKlRnIxREY6xl5dS
opgKh7hwOkL9RJHWJVeemp3fvwe65H+w13a2Xb6ZpQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
UMW5jxzpdYxLmEF0zACPMJbzJEzRwmLHJp8iq6VaCTSgABBWIyr2+YC+dZuY
uynSHH4ONNwkG/qXYZ557d1GlZ4RnH+nb7wLuhDx01IHysZ4gkgXe7DKh/J4
vzGX9JfEXd56dd83qG2v0ksVXRwIiQkQ2MwLwsRbDF3ZS+ms250WIIAYS/Um
kq1R0TT+t7Ukk3onpGJ92GX+KEHLoyq/sH+tCUgqgazoIcCgQs8AHS1cOazK
c8SIGBXhsBSAV8vY33bhV2pVpDT1YBBejTOx29iubcQ8Bas0MMI3b+8W3Qvu
73kPie+bZkI2/0qft0NQz6XdB4Of6qrOvJpZTnd7sQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
YBscRqwUfVZFeVGtAS9TTAoIh9XAGo5icdqROujJl6eWRdCgpEGaOZA+Bufd
2BgkGP12Ggz8+OJ1vAqECocBx1E2WexWPD2okh1COpPGqAOnHYHrocn9Mnsp
qNsBPKF2K/HNmZLDJe2BXbkycU8XQ8q3/lzOMvcvFOr5DBTaFdE=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
kg+OeuYHVsk/ZrWv6EGJ0zURzKZHZ50qqWMjYa/1xiHzUDF9xWaOOo8kHWc7
Lb3aaZmIPnU+iMnG0pyfOLVnPRZsfSYU1ALgZDzlvFb6QnN2KDzz4PPwhejK
30csC264HUu7emkRVNyVUINn2NpaeyI2G5Y2zNcI1J8/ajf7OGyjQcHjDjHR
bTbk5ndfOJ5v0KR8HTDwtqR/ILtcOHlXxJphLm3cTwwixEqijd0fVA9g3GS5
d1/lxcVNPPiZICpVqn3eFu8dKGP8sk5yDRaBJie01t43Ar4fEgeDrHHvdIfJ
Ddl4MVNinD8E7GOBfjOlUy0RwqiQVmI/5Iin/HcW75NatbgKBBUrA2KC/8xj
dPxtV3nWQ0iBbF2OjE/+tm6i5/DX8dCs4T1GPF3cnCqv9df+E/9GrsXBFIKz
gH4mXi91BziV3W7G7oy66I32CWuU7w6OkxirPonOYZQtZqFUbPOE61DedDKd
SY81AN/eS9cRLDgj34bNYEToRBxhwJTp


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nY0K+KG8uzA+0gTt48odofK7s9LoFM/xKoYwRv8GpyPQa2zYEU8Vyg3Uv9RT
lRxgrkbQSXaaPycj4A+VWqJOQAo0xmOQQMM2phzzuGdyzbQqsaKdird4EVet
3X9ll/4ccRhIFFUgV8mCCUlmfLgiCsk3b4eFU3tjuUpMwd9sBZY=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VIz3+SHuqwajRVr5q4y50inVDnikN5mZJrQlnEFJ54Dqoww2iUJAVZb6VBy8
ogzZeTIV4gD/33upOW4p3epuXwuaMYQpDG5kPdUeAcEgAeSQ5Jvp/5f4sJzI
R0FN8/ULfgVpYlDaFM67vcGEAtnl7NCbEi/0/fS5nyOSTmbCHvU=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 8896)
`pragma protect data_block
877tovNbZSQIv9EGTKdmzfOxitoKdvwtAVHF//iOyptznphA76o6AOOuYXkm
+aqoMhH0JGrEDMWbQyQRUOD1easychbh/B0BYneHaxniHHLd72ej438k119U
cMFnE5SobV494NJtXINuIKtLGqSANuEwDqLRmEPpNSNMRYWjYL1vUhddf8Jy
/5cAX7iOIiwqlFgRyYx7+4+kZJ5Wnpjj46g0NvGHwIDFaJ3ktefaOEr5wX6w
RtVoGOje71TSe9/Sx6c8Oy/Y0rHK9wrml2iFejyDLRQKP3LupzvLjQfPqISW
QHLizki0H8WZQ77tmKqyscZYNchfHIZ15JCe5rUMAhQfF1LEwl9Rz9hwl2b7
Y+V/GWdfI+wve+uqxgOCCB3i+45ScuRT5+KYxQcRvo18BH+jkbfehjrByb0x
EclGvYmeabbjwc7X/jBSjNlV+ivDvwaqsyDKEdSRMMvmXy04gN/7d+wL+9L4
FK5SR5x++lg16aSwbYVGg1JFaYA5UFFulWuI4ePojddDQlX19c5CVuThjDn1
PyJMFBq1rEkAcLTFsEQsVsb08f9HxGrcfgYgDEISk167s0/QyW8y+b01iFje
suOE+VPM1TpeJMQH8mQihMkqk5wvyX0oEMZ5lbXm1VnskIbKXRmYZjU1RfnL
mvcGyI8ZTVHEgxS4/E6bLuS3lhZtpip5XJwKj356oLM3QuZNjgvRgd7Qioiy
6w3yTwUNDzDu553Kv0XU6N8R3M/c4G8wgTtRUtzjaVwqLPQB2/79IUwzdYzZ
mjQHBSTxuKsAfa1puuQ4F5XXe97IazJjdpKhqMuKilq2pcN8RtWT2khXVrSU
1t2kWb4TpI4vmPsWB7xPZSPrzUwlSdlhTwg14SREUQqKPsETMMqx5EBz1adD
p889s+02RLaMB6Ii22BBTIluQA3/IjtAh/Mr96AEFAseHisrm6+t+Lc0xOAO
I2CxxJKAx5JjGANb4MDkmGdQcf89oG2hljKRIZ/uPaxc5ehGDnKlXzWp4Cul
JCbrkJIjmYDmHCcZ8OQn2CwjsPQoAu2dWqAaSHmvgaABs5M1gvax+8rCBuLZ
5g+Z6OxSOHTFQF+iI80VXrLEppeepSPj7rP7wZ1+l7eiWSzGaTrjKdz8b7Ou
jWE+gTfa+L8FOYz/RYjmnZQBmqEmOGXOQ4LY2lmJGeQDaaxPsDrllp0Y0C8V
WjAQ9ijsdbhZg4E78mfHfISpLdW/m9xNxKsMRTyySsgRP3szqSVsBkzCWEul
beESKo7EnM9o159d+IBeDLNMesN2/aH6j8AM9071Nh5GwPZRTgTdJQ+9YY5N
rJKnLfO3szpDU0pfyU6YpNuVRK734HnP97LmOkUlu3HxxlbNavFxVySoyY9s
P/gGqNpX45lx8xQnzr8uRmPpxn+sD8EzjrEqV3A+motmcdSEheXlg0xfNBMt
DLsY0Ut7EuJ4seKAk11s4jGiz8BKk0DSAS1f2aUyuJheg8pdy6+2a2ds778A
SGu3OU6vTWefYs1hVL+XpKH82zpWXghLWP3ey8lV16A1zdsWmI2oRnCFkSU0
bawdIAQjTt7wGPHHw2VPwvsqYHjgC8WwhoTpyFi4Q9KBfHLdNiYZA+LcPtI6
8E6Sqnt4TUj5xkvoCmD3ryb4xrN5mCq0QLgbX7NTpZw0hxHTj0kow2VorUNB
svlQnywr1yvNX8DJmdfrKiU3Lvdt6Oeq66mU0vNijD2NaoAvU/sOllXt/G1d
GtVtsMA47yBVokAWsGApjanBtiRr2FllWdC8dak1W1Q6LbdpsTF+Cg9uV2xi
RVECe1ThtESiuJcZriZ4BlQ+ED3GY4Aip8rj8PnpWug7Ddr9CYRFW3tEkBVA
5NFicfcD1RBvFFX1vfeAzYD1jZefUBZ7QvF4mfU101c7RK2XTIBp/ZXo3MHN
/wQX/0AlCZe04XWNrqzeg7hs59VIqNZxNXMj1iDeKFnkTe0Gp0HtQuura3MO
4C29vsQnuBK7rt+kI/Snzs4E1ngLcfmkA4lUBzyxhn9Do3dpmiMDE3emh13k
8/0uz44FAnAw110yEfTBeQjtsl0tp1RUexPuT8cAiDrcKcacI495n5NktVgb
DQhkkCjefZVkV1nnc6jJsbQa/oj+T3cLqqfgIy+3EmqTQ6ZZCsqy7hZgcbJR
ZfC289lY2+EU6ybrgn2WDej6Oy1swIEMXcs2sQKgGw39vGiA3qcEznru8CC8
ngcha48IhmI2ldqd4s8rJVrHlJwu2/pfNBWCXzKjsRPjBqEhxinJCa3Q0Cvw
iBSTj2lEMnBBwyst1MODB9UidmEwA1+oxMN+cJPT90+k7vR+7hABYzsV9OjV
6TtO1GVt6Tkbjhyc6eDE/2Vib0NPwpNcqTLJPmAA8lXMZzYfeQFGrm8xMuAY
JjJyo4ELGvpM//FJfJuUgIKsMU3KtPKsZOXU8ZLArNr3bB+GNXmG6U0vFj06
lneij4z6VMK6mMVbiNgbjHu6gqmjK0d2KX0kWL8vuOsoqZu+LvuL5y0lIzVo
2wZfZZocswbDI/rBvy1kJXyfWn5NacQSxj+6kI3BJrbMsWPeGidx3+W4k5XV
mlmUruzXIek9vxTZ4jn7rYE4ggmSdphQoK3Qsw8orh61B0mmCG1hFfHwFMvr
PzI21PXUALU2t/H8skHFtjjnrGU/Y2DwmyvYVT1n7Kl58keTlsacSpA1YuC8
lqUSWCA+BzXVe3yFGXWwE+waDQ75FvDyYoiIjkvpelCi0zL8TeXzC88p67gF
wilC9QGHIqy2moTEOQX9vZYUYYStQW7MtqGI1ZaDH7sMbeFWkr4Q49I5ITrU
FQQ6k42LkCMmxWt5hpS0P224LdxRLIJe+dyv4aTmtS9wedfy8W9GBBugbVIC
j/ykZlti2qvTAIRWw/N6b3mvWkT1ImQGjpCuXx2G7m1XICJwBgcR6KqO7w1M
vKMSjlOrF/eLdBPIfSxhFKP6l39enFgDE5akC9m1qCTSQZwxfShcOGq1RPi2
fkKWGC/fHrLdku/QDAd9CcenIesqEsoa2qP4zZPulXTsl+e7Lgx5c8E4IacJ
kv5MRFWxb30P7B4ochVAgMtsvHXdG2Io+3aQtzS3OtcJ41tZ7XzFRpI8e0V/
R7bIeMf3EHK/vnXGevX2/mUuQOcHEC0X4kVaVTBrln09g94813mw8LwVwx3l
CdFeR4JCPcEOfuVJvFmMC0kiov21jE9RRLV+DuQnOH/ROhjRG5wP14tJkrw7
qpzv/c1/NkIaUVXRq6Hs4nUbKkGuABu+Q14gH5SPqd/rqsDI4mtDgCZk191C
XxKQYB6y7fSlBNwqVHqcA0PJ25bzHj/AU7QC2Tz81/DK+QwA8PRJ00+Q8LMF
qkNt5zP0ir6US//0EE7drSI8UB5Y61rDPGhzrKPd5gHgqs2bA3KYYS/1uQ9l
WtWEUxz9chFDVVd9PzOGTG0Kbe8Yv/JNK1xtPWVxnLkRn2VcjwELv5njkRG9
2HrMDKN9a5Jh3A+x5HmOpD9cAPyougupRx9BCJrTqToOwcM3NMw8GSFdLVb4
pbFRhh9+2XQOG5z75IHaFcqYCI5aPP6wpNzsVkCakH05Seg6MmRats6jbfao
cURIJO+cUr6frIVemO+IhVjXS6o6m4G9vbw2DvJC9u5s+K1JP1KSCn/1Skvl
A8aDlG30jWPYeT9jAt3YZx613Co3dN4oVAs+pP1BMXqYyCjtpfLkm5LsC6aR
3vpg12nbg6Y3DexaqshG+QVwwRPLGObuSXKfnYSRTma3ZFUBNBGJ/t5WWqhp
g7TF+nr3d28anGR3ygtppOQYoaY6q+VI8WCFRgcrWom+la3WgB63o+MLoy/i
+2OTwaUT8qF2jBAbr1acyntSnaHO35F9apqr0/zQtVivHYfQ74zRLXZDX0Py
YV8UHyOQO9VnJZNMZbbKVeNcSpZ2+EBF6szhVyl/uV/W2QIiIbjXABJpfL36
vO3rIPaoQo0OAWiKklXYpR8v5YvpvlsP7D8o484HYZ5K+rLDJoQsM3D16Csw
T6j3hrdszircmAiUQD6ZtaNsJoWOg7FBodADMB4qod7gW+CNPjN6pO9Ui57u
bdWh6fvtGbtbmnoo/tL7ZUY2zkdKiR/I70Omi0D3BxD/oUOgah9H0oiycHRt
9DJZME/FrzrPqholobDsnWr0PYnQqii4fbZ1l46ftTqGQoKFOYoUVPn1c/9z
XnUA598p3peR/BAhLzHyA2S/wp7Nt85POBaN/kbnG6qqACLsCTBMBQJSEf8T
IiyS0oEbd5h6qzgTUjAreyfLEbkRyFxS/b4E44ql7EXfWqGdtFOjZF5gwSa0
PDUEln4NockvoS093nk8fZnSuzdciY8otyN+RSsqLfkDdiWDO1Tl9O83iP36
xAfFNViZ7BGR62W3GLIfQ2Hh3KL7BKacEbvktBjxaDsW61GjY9r0t+kxaUop
Sn7QD2NZHEYgnmomBSMHhefrxbU+05Bl3RiE12iPg3TEirpenzk3HcJ4XdCU
nd9RBzBcLwqqXmzWw6OUhC+hbb+tmVZdEamsdHYiWVm3/G3cLofv6Ka1tqSm
X9bfC4RTZjY14WD3ipvd0/DfzsF8zYR98MxflA5MzcGZd1qa7Osx/x91YQs5
HpaR36xpFMYzLN8OONl6fa4VXAUczHuaNHot4N4rtpMha74RNk33eIWD8WTR
eZn/erVj+h1051w/49QYNYGOXvIrPRjaW9q87cS2z20Feaqjtwngkg2642An
3FPG5jrMcFf0WNUw7XWXdT1qK+yoEG+Iufxaag6smkdDkoiKPdsuvyc7ymkm
jOstgPt2AG6yANE2sbqy6B4A2mPuA0HJK0DvIJJ9QABnX6y6+UTyOxMPIHtL
y+eLF2gInvgGkTQ4m2LXAARqh4r/Ukdc4Drfy+0Zar4NlIOc0BjDYFn6lXF9
8cJN1I/7eO/npB3RhIJJGc0Nb9x5LCx8AaPyDWKk7o0iKCBBJLCNOnbQKEJC
rV6gnCqLltNgCXTKIRL5xH6qgDIcGUCRtF73eh5ZH8RmSXT5wdgEM1I0vFWt
JWjo7mrZGuXyxLHWtwmMvtT/YR3RcmqfyM0COn0UwCcagnvCzlSppEfxFinS
KYDcg/ZMAFxFA3dJY5BdPzEVIYoDFe2BiNZdCyrWn5Ua9Y9NLIEcdPnztIJE
sxemtvv8RFw8NkFoBmoepnCMhbNqOgbgcuiJK5in9mM0VtWaZKZzqI8vqMOn
azDaIaqYwPMJK0eV2MRbYExLUIkvb2hbuEpcNOHNdyuwHrNm3lI4sLytBvAy
M3gpB0AYhY/wfm3moLMYPAgQbIruJFQhw+AW6gti9hOIKEaHxImF26hRxpVQ
C26sj0iIVCdHyCh/fYbsFreoeILHRACsjfv+vC1H2wBcYQIPXKQWp/0fH5yt
T6+PKyk+rJRGZaM4vWbTe//mdNirRVmhTIznDNptm5k4fVfbeYMsxEqWCCod
AczydIfatfr7zfTYNDWmppbhtz8wCBgFj6N2bhrNa5pc3vJsTgi6mI93ang5
v8Z1w6ET+2PoJAgjQ3x32hmaBxz3D5KKC6OoIqYQl0mXvYpcaqhOk6Cg3v0s
B9umYsh4y20fpH0o/pEcfP7xeYv7ZZeR9yLhjsqv3ssWs2qPvu/ALJ59zbHg
johmYHfHpovqd9YaUxkbMY3FC3/6OnJEdxueqwNh5BVofyBjGESfBbuR0NBk
YmzUhGNn3UwsIDSMeDfrurlxf0+rUcavQEHO2sH5riv5lhxsgwuP2SxuU9im
rOKX6ju5RChdXHu/XFbocSGycUKDSzxYuVJ3dvaM84aFW0Fv/707xf4bkCkm
o7Bc0R0Hf+peRG5BAZbwjj5Eyz6TaSSVs7R8V/97lYroHCv9jQuWIgmm7sCb
m0qcpOh8Yt9o3/VaU6U33M2T0wCl6DBfT9dc0Tvn+Q4qmUSLKYcKXTTNL0Y6
vIj1ZbZcJejVYkp3xzlOmQBUd3n0QtjsTdzH739mbeU5DucuMT9rcu/p95Rc
IDNznI3TnQMxODooqGlSQCaX1k5H9bkchUk/ZSg2m+XiAm7VzE/S7KXOFBEx
SAnXlHnixe4yPoc8eLxjhD6WR2knRKCBQY6CC8Qmb7SVADWVSSwFYqNqF68n
BaFQFu0apWHMCzn1zHcorVICKaS8D/QF21LwaWo2J4WEchI2dAy+tpKufWAp
zyADhn42gt9POKcs2J5n0cBABJC97queAwfUzPpeeX/gXxivj5UjWXAXJpCc
FGyadbdx+bQtWh51Vl4d8pOyDOCg8d53neEVdTWtdbWZ73eu1Pw19GdgSVyx
x4lZmJ1V/oL2xeUi3VnZ9Cfm4bb2j0dsWSGHkexip2/h+989dwaNE4EQXgRd
gmE5my1CsxIY5legJnwzs0R5q20w8IPRhrvh93ohyKS9A4/f0BtC5J2p6YeX
g/2rjJgOVbK2ovOU9eiX6iWEG9KMaDIBkjA+HrE0hHhwVnbu+mKCGvM1lEle
c/VeLb0kpp/mza2Ls3hbM+GzSNlq7zuHFeVrbdtAWCtgDKGI2pWISUPOSaMk
i2NLwrgbW8reXi8Vd70UycN8QYMWpqM67p3bJ/L9JH3w4nHTrXDN9fr+Rp/P
IgICJhATD04oGY9FmElSd3Za6NGK63oSOBVzsAiX2/yLfNPPdy7xr0GZPSd8
NR8C3VW/v7OeSPrW6/reKn5Sd1iKFezNq3Are5a16wOUoRbrRORjRlCZOVhl
TrbM497Qt9r8HXdgpCxiSetYm5dUJytc/M//n/O6tU+aLLxJ/N7V8cyf0V6N
wj9h3f2pk33beSWMgAI1YByIzBpOlzzlOVxp6wTTTjnc8VFPphLLeXWMGa2X
HQNEDod9pIZpcjJNgADGBI6FcgeaCAK7lL9ljbT/+ScIzIYL3ZQpyPUdgD33
C+8oT1R78SNdMOwrdnceemuh/Uze5CO6tB3I9AQSdHdBWVi6ieia3yatPZ3j
GGLaQeqEOW+AaZ6jrAGZMfCiLOM2LMmQNbX5dy1ZOva2v8H6De125PAx3EXV
qjxpt+fM+4RgsceVy7YezFWRs0++GmONpuz+bMNFsF53rFaiOqqJ6+OwgS/Q
yyNdOOnn899250K0ibDZ9jh7/9Px2yj5Ug9fu9lmU+plFpgdzxvnErZyrmYd
L/eIg1SzaSumkC9H3Sum7ErYhIB9GCtntXAgnwk9IIPbjnmjIQtE2G1cIQ1Y
lDqbZBeWBowmVk8ta8CMJ6K9oYASFoQuILMP8ECBQqLPNOfrB2TqkM53QUkq
Bkis4e0828mN4lXrSqFDQ/BSfMy5o8Q88rOAqr8eG3ncyIC/vNrd9FHD+8Rk
4ibkAsEmJYlOSYo7RqmfLj5mOfnVaUMum2oVjM6/iM5DFutDUP0daI00Zzbm
zh/05pHDoFLT6nW+/8vE41SiBQpmpZ0g+4TZjK2yEOKeFA+wv47y2yZ83nYw
hYR9sB0Qk44FYkVbeNNf3v8OB9h+Y+XjRzB5Yz60xRdgfffKZu7ADLPd5scA
/WlfsxuEQ+J0KZdQNgvmvL4MjCoP+oM97YQ7zQJZzUulAnvuJz13/rBRiZDC
gb8ojV9vUQolk19f1M+5fn2aIIDMgBfSGlfu+Tjvp9W7yNcXSrjykUuW2N9a
M5yZiXL5SnwYt0DAfhAusVRfvUgxsknHfxdfr3iNZUZRFAqC8AZYOeKzcA+7
Nz2+pxVd/6ZabmqpSys9DA367m558XfzuOBpvLhXXb72sk3gXvZmHjnTbcDt
MIyP5zu1UQCqwPqUFmSbCHiFKpH+6Jaf1pKyE1CXM4yV1sL/u+WXr8uoJHfV
TF0XvmqiPOL3ZO0GdDdOZraDaMvulUA4V55q6JOp0vHUDoKTxyFHefNOAP7M
iK9vTceE1TlTN2qnrGOxbYEEtzZLwUxZ3p4iJiZXKeM9DxVySJ9nzuWKl11U
t0O6hT+DduWxeWuo3pJfGTtmOCjGODL+Euf+7P3EvwJpL+qa4gFZKBS1aY8D
+PZz0Qb9sdQ0bAl4odp228CNUca5c6UhRimujEy4eXOArMgyEIyZuL5fVVWC
MkQkU36l61RvR9g23rvIr3jR5/IsJrhxxgFESt9VjLN+eSWUZShIUb+CXXR6
q2npqidmT0KqHOREX6J/87OHsZCUZAxypi6/x9sOvUdvYSvdd0Cm7YJNGln5
8XajQHowFBA4K/RvBWIjEQSb07bXPTvAS8GI57tJK2BhAjqOvmSzjRlld/gq
Go1pmXe1XwIqec9JHCaQtECi44SwYOYYQgT+6uKKcIv9RWZE5HIiljfssQJk
vpbpOPYk/yg0BolInGjAD979Jay3lbALSLWY2ngi7u759ny+Os2/siWjCOpH
wDhxJYfYvaWO9k+4v9FBFtaxVR/uQdqe+KTli4qFymv9ulWdo7MgjJcRoZgv
ykTEbpUY1WRv86OZrpRtEGg0z2zSYyrUBbm/kShPyaHBD59Tn80xF9WvIiHJ
VLTiAK2WT7OOgyz+ETyuy/Qjfbddc5+E6GeeBsfHOEOyUJ/mQwVJxZ1qXya0
c9gs6dHNkP6Dh7osb5BCdFKsWoVifd0SZte2vD3aT1J93gIG8+qthZecyczd
pv9VYYrn24wksW53FrIq1LFHDqCliu2eYqExCDpiSJCXyb6YhKaLc5JGHZxb
0exiGQICUg5BUsB2r4/QcuP97xEb2PG+Ge2GkijJQPuf4OfLrhbg2PkyLm78
HaiJE4JnDn7R7zp3xCXSEMsnyLYBqpbqOv4B5ci0G1d3ifZrjiQXz3yNAUfX
hJDC/YWdrn2vqKE1W3T92Oj8BDJyCEoS0owZBHWtrfZPqbwC4u0X9JWpVken
WP+nhy/hWW6DfE3hYUeXKV2HvHFhWmGo/Rf5IJQEfgCF5oJPbgAKRKhaeBQt
BGzkV4CCSmOIb/2rn6I2tMnrUkth5d4D7wW+gMWXx8TKp89WhndhH0Un6mDD
ePYD/9Idn9/9qtrOznoH/z7f0DHND4tUcq1YE/H0JK2hgKb+jtexfTIBIcZw
Mo45O9AfJcNxYlkB6K44Ko03VxynRTuf6QHCyst62/FxdYyKg+b2pLToQ7d0
KGycIkOKV4vRNk/u3bcioz/ilC70f2w51SX4eFTOe3pNsFgHvcVIQwFu5r4Z
F8YEbPF03dmDkFPwEkfntaTzf9mGAyGSywg8NRF7v82+zbKQeiT5MvcwgC10
dRiRD8CJaqhZYEssktkw6uLdeTlW/2aAbsAZo/eDC0IZ0+Gui4CHSUJ+oON6
KpiMEA6N9pomuD3fSyjs8WBphoJudm4b90xg5fnHB+RYek34lr0qJeUwG1xF
RkxONAyiFanQvBrBWU+2pcFM2TfruVs6tzXDjbjAEJ+NdxYBcFprYh8l6JhI
SaCV/dYhL9cXiL2FJ8Im5bHU/OAvjlmVP+i+vHye/ygtfYJdKGc6YFKIa++i
RSC8BNWPEyinMpGyfRLzCl0NPxzPK3gvyFagO11wLeogcy1kx3Ro6iBnwvzk
aZGgVxQq7UlfbrsIqVtA3KHlgE2wqK39YY1WQ+/cRN8EH8qKQmNPfzLpQHnm
iWtZUKbfNYTs2mEtgkGi9KurWtBtITeYrHWISH26ghuRNctQjGxWtfRvIMka
3ro5Mqw91bMgW+vz3u6i/51VgSGSBiVLoZ+CiQlHcLksIj6wd4M8f4qy7Ejl
3071j/puhw3AbVVfjxPhDmDLuNG0Xa6Hn3lftfjmKXzhveo27L6qBFObrmoN
m2Yjk25pjnyKr6N27KK2RggIoxa8qUC5inr3FVTeQ9kV0ul9MHVLOU151FOz
ezktTJnfHQPhS3VsW2drzc9gYThPY4BNdUfq9eC9ZcOfgTXiWkFiFDyvr/Lp
AZb6sJf7ZACeKI3lUnTeTqbccM2a6HEpsRi3auvOAWgoxBveVLYUkHQwRgVk
EJTfEhT5IONDuE/kg5fElw2Fq+uSHo8GOgkFIOfK7Y/8optrhZHfeeLtH6Ve
9gfMFiOFUYvAXE5aXEs+iY3E2dXL1zV51X1zwf0gsG0RS8/m8ZSTTwCa/Cap
MiwYaWpJvY53N/Y3p63TRRg88SoJYtb1PqeMkDo+HIc5t99UpFx4jCxNDrYM
kZdtkv771fWtM14oMr+wsnqPvNKY+q3HkHXgn33JHVq/T7Rzqs3pQ6ygyrOY
mgLlUImMgZumX7xrpM1TlloZ/dF03SKzFotHv5iXdT25dCz3wUnDA6eicckJ
lkKGr3LdP2XnkdhHE1V1rI8/z2HgDmEtxOD/mLjiAYDVzKXOVUOz7nZon3Lr
MO97Uonp8FpAty7N+p4W3MCrLJaGOFgE+WdBXbhL4SSRrA/BtiWtAl/1vJbF
ZnWtvmZ5/cafFTPtwSwtlD/Q0aayZO3PL61FM3l8reEwKmb4Fr/F7ZN3MldA
01FINieFA7bWn66fvoyqThiGH69Dq+iROVAJ9U+gnas3UEY2Y6nh5UbAbYBP
ZiSRQqbxm3PRU9um4CvNyGyud3g21LjO2m6TLYHCh6U1acQvk+GQR+9Lz+lI
x6qRR2jQikxr6yPTaggYxrD20/OFZY4malNOH1pPrATQvyWWvp4bXDt1vygI
yZXiMgi2AijOBEWo/cr7bsQJTHWGVblltIODdpO9/j3Dod/I6N4FCcAVtAe1
LlYIuxqtiVGi25LwgjWyG+GNkhEnTQ0TP5wxZuEDVj+4KH5F36571snuH/hP
wTXmHs32WucA5rZslR49C+Hhru2zaoozvaB2MKSSeBWweeewnCa6J36PJztO
6aFDX4/S5BzMfLkP3GliKI82gbi/5y0Sq0QBX0sIKOguXmK7uYTKx5V3VUHc
0D689tYY+iV+V2+SmRK0LZmwf+dcHU1gl1CAouddPRFtMExylmSSuNCClUxb
lbsgtcwwrnCbySWRbsO5a4psaWjngCb0BuJ5W+2C+6LMhPG9P6f+hW5HTHzn
mDLGGKnat8jCxE/NhwtZ2QVwILT057W/efNpqqLqBjNfRE1WDPqGtVj/IxUu
3JCktk1/6ZaPMnoNyTRlw2oGQsg3QZsMfVke0+LqB5Ka6+yHCTqCE9X1yocr
k2aif+wMOIuguNZHW+vD8pQY4P/2tZGAnCij22euc8zVXAFL8z7IkjLAPFVa
Kyoh88gSQIZX4br/vmuxn+W1yIIyptZg5IMXs6aw8rMEA/nhf15+p5p0/Olp
pEHmIEidRynOA8NbkZO3IwD1JIbis8Fdz+LoH+tB7oeyx2UXma7fGiGTPkVt
jOTV/Qu6b++1mE5Cw2g4OnArcVKp32r049CKp0AacDBAw47GUHAXYduEZWhN
QQqi9WfzCbh60fU6D8bRs1nQJzhrWy3Uj0yaEMLqf9HWvetxcReSvXUoioQo
e0RklJC/izjOq/WFUTe/PdvXtZo5gU2t+KyIGeWcEXXhYPOp5puJ5AwT7brp
iqLkcQYdcBGYhkP8gI9eJDgm9VwN5lqZUS4NO3VzwEkhpXOD6of9HsxSAsFL
h0pQieLNaqKIb+xW8ZDiVI3mjkx15axRodrZSgr2J72Nt9NJd2FceIj9vOyG
1rgWxfby91IyBtFr4nhT1oQeToOeDytKc4M0nsVpWb1Cm2l0jkkoQk1KpN5G
ETX41tBjhtNDfJDH/elWIsSa1JXA3Epj4kWiJcd4G/0X1fE0nquy6qponiDz
dDzYk7M+dAa85uZC1LIhTW9i7hGaHwUiz/GeOpQa3SxqGMY2EjO2WtM0a12P
G79CvQZwJpJD28JHVcHMhxyj2qDXhn0bwoCKPFfX+b/e9wrhCPEaokl4UnoM
Cmog0x4h8x/ixZrBbL8JP737Pr3fXuC4THV79uvSw0bjTWL4/gJe4O50DAkP
8NmNNmKfBzt4GKSN4TMOjRY+iVTsCZFgNlsowl6WIQ==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG2+MchBDS0pHuBl+y3STe9preN9w15hT3oYlMFUvoDspKIpQ91tpDu0ISTvT1DX7QoTOJeuUSF0SE2LNYSzzrqWW1m5RUgst0GQqD9bSHu/zFhs1fjQ9apgL6K3Kwnu0C+aXt3EVJbFI3Ez0RKT5Zuk0iwmnTOVoSiOkVCA0wfH3EIGq1WD4G6fTTtKpNpI1UhlI93+RX5XAVIG5MpJQOX4f5lA+L2QK734rPkptY9g2z9j9vesEvym+RzV985F2uP8hEm9prYxEHlUj0I3hbIWyBjHdikoxORyZ0+BhuPd0YcXYMQACeoKNSWZLsgR6quQd0UkpWg3wdoxRf5i/nvjd5VRmy3gYEAQ3hu4gT+DymM+QNOWHVV8DowYk834uoq0bYO3MzH5BA5dGJ+hjjLO5cG37tB1zAjG6oHG7220lrZ+eJUZbkHc77tZQU6TV85I495aVtiYrumnaaB8XBkYsjl5zysyCdz8p6A+ksRdwUGcsOJOt7GADp7aw4jsfJngSegP9xcwzrIKnWR3SpAaIDYgjraaPWvxiWkYZCFurNZZS/9OTpDyoLCt7bzyppE9iVOK7YslD7l/kiOj+PH0HBOhMLWBdxoG1/4PwgmSUtWW9uiP4Wgv1HBH4dShLbkmhk5htK6PBmDMv8LmWvnIkB/pKMox3dY81lQCk4J01zACs+1ICP2a6h6EeOoa6GWxrlmU+KdPG8gHYP3hd0Zz141NLyHe2eW+v8JBbb60GiS6HOcHwjmJkAxJSRhtw5ikicRAfLJynUBmIe4UA2Gy"
`endif