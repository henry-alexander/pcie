// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Xe02hQLGOVY03xtQAF3wNJMD0Q0KzU/U1zBkXRqCGMiKceATTe9hR+ssUNck
5MRhSC9msR5f/s0+Hpmy623ROH28PKqLuRLdFOfMVvuB3Yfztu2Mz1nr70RB
G537DL6KypnNlUiXfCtMRLSmZ4hRZvl25bELozFwgU4aOHnJ3S4UPZtm2xP6
XQFrdHLKImUQWe7XXG02soyWfPrqSCFuYpY7uM6qkiHnjypOkQwJCw5iqZmo
6OPiwUzKWj5PMiOzo0L8uFHjBXgiTuV+XfGXVh38rQuD84KgSWBgGZeMfGeY
H0LcDt+7CeAj8sUYJyL5PPIDohkEmdArG4aWZ57W7Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
l4L3UklySKb/ZQeA9ObDv/7xfLljZoyQ/Ee+q/f/zDSLQWX8IsIXoHvLpyzA
vEJGjB87el3XIV9cpEnTPeLp/B7iGO3CgH1A/yP86NUHaJJuaYPxs2WazDxI
i8CcnP292Pv3ouJDnw1LDNUJabjVeePiphN1Ttz/Vf0Mf7eYx3UeHsPXwNmE
hMk6JCd1wm81zVDcfvQyYSlymSWdxLU96vn4VlcEU2iX2cB5CEPgcGYAf3OB
2OMv4WHqCc+hi/DdGN4p2Tp71iTM3Znyii3zc/Vgiz3DpM20lTt/laJNtUuz
tixcrPuInL/Ah9+ZafSKDDnvSR+1MrQ4AHbu3lvukg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Og9bhMxJEwKmKrzkvNW7T0yWFzwT0N5jDuwIbVECeCvtiSjt++p3ncjydxUh
rUSxHBagkEZkuL/8xoHgWi6YjQTXfULrDpbgTv6A7ACmtZlpLhrdULAfes2a
XB++tj56tu7wOPoejOmIAXETxFAXjV0NlYHoDGwLA+VbkRl9fW5zM13JgZzf
Bn6d+rP9VFKHGd1yglm6u9ITlbEIWbXamxklgDqJgYARF5TsmItm3ZZYUBKT
XPs/RfnYkv5RUx5UoYeK/+eKTUwAVcypdzrPc4JnfvCAKcNQjaz7d9P064HK
AHje4vyeibAcSJwcUe2fl/LhWzImkAwIiJ02+p9JQw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VZWIuELFSJeuxNtNLIMPquTcKCV4rhtI0p6B7bGhAqs3CCKPm6whtRBoyY/S
vw2VO+yCTu+pajepuAa6rsj3wzCkcFrJ7DjaB0v9Ng9rHTdhhCs+X2usdIKJ
2ABuSpg9kwQtW6y8zfsp4JrFJHhuzhg68Mg6ArqWruiZ2wouSSo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Ph7Xt7hkJxq0pAGgm/km7Su4mlGKHMmXeGyq6mtkovevuKFB/whW7XwGuU3F
Lhvq2FuT8Kq/hc4CTSbDHxgj2hsUcpn+XCfMq7gBfingm2GPlG5widFVT0CE
p/PjP/v+TQdDf/9yRYbXuk50XahHspeYLavhxHlaZuXJudHyOQixQWBraGqB
toIamdy8L8m26mDrfnirjtoAe1ckr+s7kN5p/KrjQ3esuBpxH/g9zeyvTmWJ
jsHg9yfBy2TzlllECKg/rIGm53BkIWUAVpeyfyJSwm1+6lsNYjSWKm/BjHtQ
J9puoByKq4aI9CCW5w6VvSz/9Fy9QviSxJh3gRi7B6uGlv3T+FQZaLTOFhum
NkcNt9bK9piBQO51JuTDJeGoDb2/CPDUdW7ktl/lQQdsbzLKTO2xnCIyY19j
NCNrqEOBcp4CzDoRmIRx9jBsNE0AEnZ53jrnpDdlvk3n/bvZPfN1iWA6+JZg
i5vjD5ClAMLGZQLVKQwkEcWhF2tzm+xX


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MpDDrPdmkvZT9Dnd55F9kBxClLtjFrntb6tixD3/WEM6KGFHw1dbLhA5CqoC
BffHuCx3CsjxX7FyXflNNqcoZMiORGI9ZmutAumHlPpKtKJzr7BpJLgGlX5f
ETKx4uIa6NJN17Z935Xz5FFZorTwwvhQbmIo6NniU7TgSwLGGXk=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
UH9qQ5cmGUShkE7ewdMj1V305CD+x9g89aTIjKZikt39kay1ZVJA/tb4Tp+b
+2ADbsWgcAUW4jFPGVTJcSCyqfCVQbRzB0yTc/0sYkJYgHeWNJnHF2a+1tpo
mC0EHYZF8xMHuV0ae97onPCpH+6TWBaourx3F9TF4FlNAAEsdqE=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 9632)
`pragma protect data_block
xlUwraXeXRcbIpUAq9jAhBEJFZmKf3YRJLxAAue+wBnnu0e81btdm0OkGDhO
Za53ZuveL7OvE/dR7zUN9WNx12Ut/yUxat0kI67v8CbG+PYXC54iiLqqAmUv
8Hv/qKXt7IwnLUxdfEQjWkdG7OHIPZW9GdIgH30UWm3bqp4L+Iy5zy8BPg1q
cVBcTWSweVlngfWIxs826Qfi3tU8QBIStp/UyxMp3+R6LTBi35gM4Y0sgMvQ
1F2VD+vbz6IV5TARdc+blFdXC2kELagSx2yYcZ5EPanoJYazZ//EhxMvI2me
XpEuuo2vXrrA0O3lWGFtWaN2Nu1NN6Scs38oxoNkH2g/X+vWZ5F27nmOHNp9
rYBk12qur1CoX+HZzik5gGND43ueSGR8TgAA8J8N6CqGJa7xg6ggma+e//r3
xrQpfMlLaxdy1ST+MJNvPqk364aWowzcGWM2bhNWwAaEdrjV3tB+RBbT+stp
LyGEVOsI1u6mkOMV1A16IMDyb0cxN/8XbnKyESa+g03Goe8S+KaeqvyzFaVz
7zZ7G/lvUNfFs8AFUsb11Swi4+Oqu5mX52WbR66MYluGB1v7WHTvAf0pmYwH
+ikg3llHfzbjqMUSOqU4OFRWY+4JfwEKcsqkix85+bov2ZvXpXvDMm+6imAw
PZ5FYfBs9ogG1thI94UziU7SSyGld9DiDSSMkG6eztLo1Q+oreKIqsAgvCl0
nepISHwqwmvteUUjmZnSa5QGlq7XiNp1JpufjS/Q5jVbfZg3Rz38iYW1pnT2
pUElqhQ5QPJGqb4WMYm5niQ9NaSf1Qln7uGHASuMN1L9sQHTxfshfB9QySpJ
rj6I5+Ml0Y3wmPZcfqUKZPRPIrhsgJITL6hfELhlh8tDh5JVqQjEhOXila8u
AlbEfP9r4NZGVaAFjLvDWQeF6ebwLcHZooM+xQwVeVoMiCkeMNKs9aIe93Zl
Uk0t4Boc6t053lIhOA4ge9PDt2rsnM35/1SahzISwfDFHL6loGshd5yzH163
azlLiT1P92fryBiYlU3uSMJa1m9//HSJ5goloh3t8aa4B72gnaFFlRle7+Dm
9XMXpN9CtrXNFy+YXvBAgu2q1XNYHdgkDC/RcECicJz32EVXPRBXf1kP0m3S
rW6zIzUOsYjk2kCrgTPKq2ujkHIJ35tw4mQS0KCX1zMN2FrXqaa1yu1hcGUe
t/Tu87h982HYHXZA8Dvoz+Qr84WNLczeb5H5+GZ2XU2POOWtOXTrJAJkGUpS
yAvz5qETcFWvVk5zrZ5zm38XlndqkK3sCx2iZ/e3nKM9LZFm84by7tUaGwwB
iz+FkUJ035l3c0es/J/mqUeikzJn2Kp5kXPSK39fyC7OktVMeK/a1UU/Mbgz
QyKglocM9oox2FD4gE3nC3+ogiud33TQOCvUDWZXlIqx1F80aLw2tRdsKqhr
XmYJTgJRJgfYsRAxuFLC5Hs09ox2NZPKn+1Ez6ngjXmvZqTpjTpNs0HR9o9+
sUqziZeoPs8mhJp1iiMDP+nlwwFexs1XDf7O0OrjJ2VlfMlTo3fnb403Wl38
+mCrHFbHwtHoL3OA3IVcaGeQkU+cbrlBngr/uVyu/c0jAaqlK3+bvkBkclzc
vl9ZpThZZEZQXXTC8jfj09yon2zle7kmV/AsWg55fLBPf7n+MThvfrLbYNXu
wLEIc29WsKoU6EB444xVv2q5JTwJlhn60AFVsPdQKLN8/njMP0SWZu4x1n5x
RyqvyWS7IuLreE/VcR5P+VLM7IfaOWdOPHMsAC3vXJ8Xui6utymrqw5ibfxk
lS/WpWLHatwPBWosxu1o1DW1ck++makPtOc3xObXi48l92UFBi3o2KvBR23a
L2nEHXN/UJBgN8ODD5sGV+rYCt7NAum8HhECXFoCMomzjyE29cigYEMctR2A
a3Crw9fykUwZvOeAHP7U2w9C1bpftLG2y2SPBl+Qnd0ZPOBdKrFoacuI4+/P
Mt38MkVcA9GGEyzNVtHUEeuJu5RemFZzQmVCRJUjbxes2vLseZFjkb/VR3/9
BpUA43BZKCYq/v5Y19HMockN4zMUD904px5KH3VlMhuU0NjrIzZ+lbsKvi9r
2hX+G7c58N+PcpS2yHVF/eNYrJ1fYwI0qjebLWrOsTDGGgtLf3Dgid3fnoGu
C4vdqEWfDHdHPBasvU1fYOe9/ix0mYbImbT7+MRUgiJ6+N7CCM48p+AyxxvV
Pb/sSbDHnFw+kFl8rBln2t7oULs4SvhXz3eKM3JOGvAjnO4lJnRNuETooLJP
aLH674g1yvryIRp48iPuaqzFt9TvpDud3ZUm046BWqxDFbCWtlOsHqXUWqT/
08nwQ6qzqvMScJLFV09fa0WYD7t8sGKvqfHu49TRQS//OqTs1C+eSMLa85hM
zF3qXL4oWxCjU9pW7KQYFv7zHpThwZE+nJ9SJE5b7CJNX6+zMyU+jAVUoDFo
3z6hsI44W6sklnhmAWdpP5aarEgu0LxVRQiBNAGDPtLbmaBbyXZte24GNZ/K
mSfK6hoj74lGXgN4c0pgD0iQCsPLVq3dPAJ45asUa+gFHyEkGsEdWuFvb+vX
ZxoDp3Vz+FEXsRjyIoYnpcVLvEnmqs3uOnJx+HYYHOqLzDYuXx1pO4ACam6Z
vacang8Us7WbmOcugW4lbzPRNe5Q0YhK14A61rSjjmeF668tZfRd81wTt7wk
O6X5isiwa99Tr4AQit6BDGqXt9rayBp2hJ2XaNjzRuTFlQjZPcVLeF7gJ7iP
ZkV+Pv4ljBp5MwTt5EBqvprW8t441oPOIGeXAj3pXaiMgDOgok5VI/f6YA0j
tqWWOD9dVVxFmmpMDU9lWwUqBZfiy2oY5x0s+Bcz/kcUUoyMezvThS0tpSSv
hOU0WPWG/EcKDUXHlb7xTgYl+6SZqyngPMmZZTzsjb+7+2hpWOsvbRFjDEsO
Fa7goCt8I3ykEq/DAmdKhcMzHvYwR/CJEt0UsSw6+cg38zlIICf2UFRCHER9
NL9QV2QTh5Upd+o25fzbIFVTehjm8WgPG6xBcMT1UdlViODcjIN44HLiGQZU
HQPosi9pr7asOiey38PJUoIyVuQWU5s/pfQMEXVjibwUYTt1pUzssAkdwdxB
PjbL3UDbPKRM3YM0+PbCmaBA4mjMNpwoVbO1Z3P4hCdAlP6nCfehl+kOeoRm
1N+EhdlNCcMRgwFC/7LEyEvd3M0knZmzHdDlCRZnzZDwQIIB1irEdkrCl3WT
7xL3aLTbWlPVDLmBmm/k1Q2NTNnMKhG+p72L5PiK1IK8Uzbkqm7D6smlteRK
E3cqwXDTxRkZAHtnbqtXiW4+d1bzHi6swfVVLCBC0oHsDdueioWXXFWN4FB2
nlXpFQsVoyFoe24K/EKmBTm+UKChxpvABx8CzazI3eN9VM235dOHHb2Kb2Lr
a17pp3TdW3CTbNzipHy5pJK1y2SMUyoDAoL5XghwPjZeONPatVFKCR3W6ML3
/FiQSIwDgRtDPC6AhoaC1eJF8Z6mGadCburQ9R+anDZnBq5JBySthy6pahGu
6FGXnmP/kEQ8/64yYiORCktAK35+AiOg3nUZoDWiLUvLuxCanTS2MYOrEMJc
Tr8blA9cRxxflP6uOpgOH9NpDInX3s10AH2MBxom4zE7YR5ApVTaF9yD+W05
fsD/+tLstPXGXCObbEbfA8MljE0zEYwnSXgiiXGN95QQP4bF27dS/VTxqBEf
tL1ascraZk9M4CzgnSAZBIIKHUQtNPrGeNT2ADWTcv/M9KrZYTklpgzT22Pn
5Hjy3gqbjnnC6o1Ww0Ix4B2mbmtXjeS54Xd9X19shFl7/eUomdWX9pTVR08s
8jkKFlKTnMH0oThC8Z05Xdanag+P/k6da2FOka1MnVJqWCUDhiZA8GqqwusE
9kVNWH8Saq053l+e085c4zIZFpXv9ZvnpyHl1ZDvsseMQVNbXFgABm1vaPC4
Ro9tam6QA+9iVXYuIJo+ctzw6ouLiJCunlopaupFDQ4hKfsfChqrq4TZyxTA
29oi1AytXS4M3Kh396GHTbDlNCzNHWwWvKeoKVP2vtL8oGpED3oOFktvm6Ho
ZpVbbG7LRY71JPa7dbNsVnh9gU8iuIBqqqp5nskoBPPfIPEeYCRkkl9VeKGv
S9WWaPqJEqFKBaZivGuOnA817Eh06nzbU+IBJ8splLiS4ytxmNkgY4LtEPfL
FOoq3CZfdq/e+DgYoQWg+MJyXU93LcgG3sb998O7Z9UnOB/JfMqz+0rkSkO6
9Jssz0fXs0rumzk9lymfN+kZ/KKCm/3EpFo3iMdHu4ZBXVQzmXdJRU3ELcwG
Fmt38WpouVSs4B5yiBluLQpqQUNE+YOWPoeL7xQNF1xTTvtWTzg8s+pOXLWm
tifWvBMtBUXwuQmjUZB5cLmyQ7+HAiAP3vbu+s8hWz38jduYy2n6JAN9spMI
bY/gcdHZJYboD7gGdIugP07pFNhQRFzLYD/wxxpKLycrOZruYoigaTwbS707
VovnlKgf14rkUgtl0DtIyZH2+/CnVtt6AmJB1prCU2sE72WDDcMjMiRDE+Dw
/OByJebUSpm86PUIP8PgYfHbHhDfabnfQQcEMbLgfnS57jc73uW50MNyMli/
bMQ60+2HHKJYelh2h1HWwc3xBNucBStulZQWkNHowk0sTNEOB+KetPIRmiax
sP7vPxMGpUV+el7q97YXJ30CkF8NJ7pM5a/DEwY2Ovo7fk41QTaZLOyDc5Cx
6r871hBDmUQzzBTjK0BbjYZ057q0G+h82COR+WxcdC4787z+aPjp9Yyn1dyx
RasH1kcHokkpOVopSzXtLaY4JbLrrLWq9y/Jl5Ibg6b7I2ozEbKFdBfuWWts
KT7vUtgVD4LZHjZJ600Vg6uSxxwOAwEhHkHRPjU9o39VCA2/jwi6WA2xB0BU
qvLEXUUF4a6mgXL7jZKmajL8UZ6VKiY5BfJHtMuFYbaZ2sn02FbFa+zsvPiZ
wupE1Vz1ZqJdAHSKrs013dxrSuOFWYql9r1krewrpCSvMnOUTD33ViErEZ/e
toSfmH9889X4e8oF7TngLYECxacA73eP8iBldeONY9/2blhFgKYqD5HjLuWK
dBGa2G1EB2MqLmkphBVLsFrxuahlxL+/lNOv5ueESVSRL2ENBDwbEX4IUgl3
3OZnqTte5KdueXPld1i5ud126hr5WevaJsMnUzkH4QT6eGyYVvL2gJmDaPCP
0KTBVXreu0COUCo+vKoKg9R2ttP72w4Ow/x7lAw1ReOTKqGL6CbsmMEq6kRj
LEUC2hEyzcZixB/i4xokqcpIAbQRkUmfPXJsoCviqehljWqIj6C+kJjhrI9i
0VNLkiof0glHKUOg0uiC6RrQuYvRjOvdDpQlKlpU+dZFQF9yoAOweQtZKJ6u
wnE+e+xdM9gI2711ea9LPD5+3Nu63KlemUlQbjxoTaUUjRrZeWZ90MkBnitu
jr1SZPmNA+XcZlK9iCN/ojWbdVkB4M9LTT/1Cw/4V9pLqSbxMuw0cExJTqDO
wf1y6lBWiX97zAxW9kLVFOgTlyOscdJHzPFAzrCdPJzdSjLdsBm5OmiST3hv
OaAMVTwXf/o5NiVzrfGxLOckDpnjiFDh5yfcBLk5cPzWwi6j6rMUzMo8XoNM
KfQRP0ZLtrUjt9EJqHJrbbH7UbsEcwooPnSK4cPJ9mnGglXRlr+vR7olkku0
3CesCvTZJbqyv3oIfg5KTblRVSgoqFj66FImsTEFl+3tYB/4dMDVyPr2XtkG
xpY0xU5GVeJpcxqoWTU6aloH7XqrvgkoQNE6LFVLkFfih5prN4nIL2u2b+4v
34GX1n2Xyx2FGpbEAuli4rjs8BA/7KA8mx5LkaEtIL+DGIHRbQgETLKdfFT3
11Q87/N3IchmYR+k2m8vANUAAujlHQ7A/H+Sumf6W0X2JlsC+qB5bQYcpqiq
2XNpgLBXv46Md6BkhC1fMtEaYCs1b3TmILSXiv4XSY9Sp2gguiXDXE4LPP4f
JSz/0y00FZwsu9F2ZEqV2UJysOV1iJyxa9MXtGz2L/osXPtED9/kTifzb3+b
LLX8+M5coHVucaIsm55DnIBTSQfy9NYyhVSTUb3PN8AfxVpzezUsYdDHv59H
G6wcmVAFQvaEQrOAOeSJyYNOGmroVm3duqurNZSTADRmoMNK3AUXBFgoOsfF
sC1EsKaGxVLPuHc+abxgaahqSFwsxSf1ALF072oGol8aCoNhNYqqCd2jAQuB
oyl+XGLNq3g0+f4EhkY22MqdzeuYi01lNDq/VQxgk0bAaBeF5pKjs9zIMkU2
n7lNu0m81ayCQZ66/qSc16ZKaT18JD4gSzbvJ+kohzy794rjMYCmaj/1DoIl
GNQJYwD4jYUVWoLpZE926Uc5DaDj/zUOhksfDr5OioCcDLYgg7nlihZRHlPz
q2TvfAMsgOEcnd18oL5jLv1TpvZGH4GnUqPZ81yGt8d3Y9sMyzmKahMmYhL9
dbB/RI09ph5i/ps3XZaPyhh7PThCmuiC8oRga5w9LazNm7SB4cYtlRj1I+vT
jsWWA67IO0lx2q/wRipYfkiaL1pDHC9Li6rBS4NZAxLUSGGGBCQTNyo04Tkx
McAYEPTt7ak3BOMKWiKweVRzNDpOZILsfmsIbXhiLCFRGmkRbJybPLILHhR4
c7EatHawqEFnlMh+mNZjESECiPw0pu1lTfSoJz6N3ZexyVxE0bu5IpQX4GiO
fZhujj5RU+cGbtbv52+M7rBnVc6fSV8iVJduWONwxAplWa8bh9hX+ujFO5aa
7fZVWt2PzbjmTEGtKa2I9iaJLhGJX1fzJU3NUDelP2LKtk8I8iPlkwJfhkGQ
o+AcQiXHZjwIHN0KHHS7qd+kDldlLtAkehfsxyX0tEsNP+agmNrqbYCnAqTu
MwJPbmC5EPi5sOj4h+vRxYXAusu6481FFr0iuOZOwBb6+FFlQmZUrmAdU0ZF
SxP4k+77vUn0VH7DYnpoZ/404zoWhjwVtJwLSpFSvNoEzP011AtylDEChiKj
Yv3J8auqoMneWNBH1AdjIdxMh9xOx7DYQ+kA2sjJcmWby92c7nSe9y84DPlM
56LRbxROGGUIpveiaJBfFzjhH5uEZgS+w/m84Nrux3ueQH0ONlEbdraQOhz3
yl9evDs8EJG5mXYiGGogBziZfpHS6A/eOyViyOY+ycS4Hvt5lCzNAp8BvhKz
x7t7HLRE6mYXsiyZwtH2kpQi+6b71dSLSG0T4HB9rxeQFFmm5Yv5eL0sp83m
1sVwVl+do7owXLBB/6BNBa3tgqKT8dky7CgPF19jondhQOYmpWEZCbpdeO42
vTdrj5PDcAEPWWH4p8Y3vrQ7w2a0zbLff8x4YX+V++OsBKbHlee5mh4yijF7
/6pOro9pxOwUaHh9Q+BaQsExjdUCXW00al+Sxc6dg7yaNOSR8fTaTJSyliQi
v8PNm8/zU2cbLL/drT8C+JPWMEyxPqJFz5G9hZxwyJ/MxsKHalrEdRQwukmo
YcYN/dOU9mf7N0ZUVNOzktohXpCRxqGh8iO1A/DkTJBBCOPbggtIIZbW1c7l
eLCfEg3Uj971MuTx+xOfVbV7RvDb08DaNTTiQvyH8f4USA1K+lMAs9IIssB0
MyQs7g/HpqR96U5hg1LGq9+vWOpYVZ9d6XOAXhZtONeyuqGYHMUgDKuFX25w
J1mNL1wnhHc+QhPva4KLfCA6Sp8aIAkcUlu0yBFh2HeRzdgaikL+2BDW6b/r
moY1mLBgbxzhPbjLjbJL1LKge4cqsL79MVy89/bz9K39hDJ6fdKiVj0vzE7u
adjqIFy2usKeG0SSVScCwOdKDe09jaEIBSORYnWUFi54VHZrSryFOgLLX3fU
usqtTHcUt7vCTUjaw1jh7yxxc2xrQ58QFKTFOJb4N0UwLWBisbEVKFrxS/zm
fF7tkD9fCMASSTsU7z5hVGNm4CdXsqIeZKYmwSMyTpmS8hj2n0onwCnOdSKG
WrgVvFTzGQdXeG9jHaUhwokCsedCWJIb8QwOLEeKu5g1w9YXJMB6a4v6QwWb
0rgyfaHv1NIrh3vk0euGRApmDLAEJVwhAa24sRXOlv0SK7nC6KxtXKAes/d0
RMkUgrPuwgqwA72zl1SaD6y4slkOxiHJKLSamAkOvy6L9SNgAiRMfazSpKHM
/ogv6Xo1kLWGbSJ2wM/qWI1PKGId9LXLFAnHYalrva+YWVFyg8ki0mJbHCmm
jn3Hw3UEtR9ldxbEl/BR6WBK0hLC+pgZw9CfSAIHAyvq1kHWhqXIdaY/5FkG
3Nf07XeEc3TIYaPngb9r120fM92U7O7lFnTGN9zsmeY2OyfAZJNED1ZYpQRE
FmIl+XtpEm214gJGNtG6i+km5Qo7yCH4x1QNDCt41zX9yq3+b5meuZfIQ/Tt
P6yS4e4viQeVNNKAYBzQ92Ihmfs7GFdJpkxREZErsilU1iN52wTGAcd/Ujzk
+M9MLfouQzspx0nlPOnR2G9NoeHLi9hPrtnfUMGAU+Hs+6UmqJqaPldufjQS
9OJja1AyTILJipwqtD7W8cJneiUKXvhCY5LCc8YhIQBTfH7Kt4vnDD1Ez/RE
TY/heL6lWVvKDt/3A1RyY0cvaciXn1r6R5ew7abZZadhIxsBxCKSBFn9ZSa9
rnJMp7l9wLw5BVLbLsDGtmPylG1DZ2/5uDZDXWN+Q6btDqEwETrdjoQ2+MZX
c3qj/hClYtmCxOTZhTn6a24dc7SzLGYyKp2Y3l1cOB0xs5nm0EGaFjMjNdEW
H7NqZ06FKihQ/O/E9grp5KQLNb6SSBEt9F6dHLOTk2DaznFTjMZ4rRxViYv0
LuggnoUdBKwvR5Ij61r3ezKnK2pq/7ZHyAvZvarqQcb2FaF+ffvGYqEeufOI
TIqeh5U6Blhp7AGOGUAX+BGjHUsIw3LhbLGfLMrPRbGbzWmD8A8j2Lbmzjm+
ct+DYOuukYVnKTaL9M9dqk3CFz0U8zRQ1FCRPB7wAROVvdBXzXrlODt6VfyE
yVrYHPJdgOD1yJo+bYaBKO4ygDd81PYeT4VHF7Z2sjqcRdn70XXjqjbWfw96
sEMGoPUDpfom2CB3WTGyKWwe200W7YMXJOlkFQamxoVxig4ekOP6OjiHODyr
6ik/JUXbTfWwyUSRarELrqFZVl7oJBcvnS7Ja4uAcYG4XKRKejD2MLC2HG1Z
z+b1bFzfcBIIow/HCJrSIn0e15ZMWF4wOhwnOAYqmitvM8rW1yCJAKPPYJZN
/KQyqeeEDlIX8F7I+EGO96L1D9nEtzWWgLovpACKU5Hb9ZXhr/nuClH7KHQu
aCLJme2+fNlfRLDLaPpOpDQyuTD0JnzIp7/3SaeWYUy1SWtEFceWHxkOy/Er
ksy91g5QCISKenbCMAwR1JYEfu6DOkFfUinJhxx0Jn2rQVbEZFEpMgo3tajZ
4rrziKUFqcCrR51N4Dn5pPJMlkFXmF+PeXFGpFh7TCnhMTFQOt6uqu14Ab8l
CEvAjSOMFf2SoavRVLBUw27LzfFkZ/AZ+1NmKFxbObxg4xfkIa2wAf+0OPkh
JqtDrv72VfOkFow3s/5MTtYxYfNy6fYjZzTMoSz8rCiD7xXJWR+HUBGG17UV
7kKBC8i30RwgL3XRfDj0wRieHs8jatvPmJMRTmyhR4aLP9lpZaig7bOGPI7D
adRK4zedUcBd7w19iB6naiqYKI0X0wck9uyC+uZjeVomPl2vOJRwxkpv1Hx6
uFB0QcinHMNFqiwflfXNoF93IYW/OFnmXq5jOS+xgJKAvTIY8dlORittpAJr
4GBbfEGRLU7pm+4r2356zJ02mot+eH8fCQUnUMjYaN1QtCFpMvhmm63fmsVf
4NeciegtJ+ujAnkWcOHD2M/OIGdYlgknY1T1b533UMXIsUF14ofa04i1KErd
l0MQF+XvU2ZlYVI2VmvCgpWJk/c+THRao6CH29QEBOFQPFa+WvhfbTluhCVo
6ogT3tAYFMHdzjMUH/gXn6yA12boBudCc0jzjCmXzIK3fhp+Z79j+lND4SVb
Xgh08rAN+fRAKW8jd0387425rWEZNheixmT9ljzkg8x3z3wCyZ8aKdXFagLq
MxKT+yjwGAhHVYPt2X7e42aOyKyqi/PhU/3335MnYCPMACrGElOZAm4pwv+0
bUtR99KBrL3twNfl11EE74zKVkx+f1lu6ocQFOYKMurgGYW7RTxTz9J3Q+fm
fYKryq/25+OKGahAQRyz6NY3DS6zOxeFwE5DU0Ao2zE/zJ2JE+/zjEKvnbvU
lCEbz5Qlos8koa+dOaEfTKoUu9W3358G1E0vvT1gi1esyfsa2vrYGTipmbMg
VP2YYoctFvwqiFjU4KJZP61FM2zf0NEiMKYD5IpnDJFUtOLn6rkUIzMQcz+g
tqkDENLgHFIfcC6jf1zAFX4CNrv31TJA2fvfNgCZ54WKGady2675ZHaucdYz
caS2wLFc5/YN/llycl5RoRKDtnOj/OO7wRMje1RQArK5vz2DPxET2HLuMkoF
Yu/v1PSHpwOSGM0tymDL9gH4Y54kpJqTBOCDp38tNQ+BAGIn2XHWM+gtvtSa
mQxkXViVNiq34qEI0mHUoAhuWQEItylSxBVRnjG6V1hM3vZyvgxBsFfpr5b5
WVNe0OhnfhL9eVtspdUES4+QrDyX0EUH8+Yq0eqqIVoMabP95+WT8gGHG9Zb
EzmAaOWH1QICWKq81uQvXbfLasTAls9AWEaYZc22wH0XofuMGDCaycftJTzf
IB41jFYbkop352v7UZL6K5XDRKBrw//NjE5HhN/nvFzYXaXFKCmZSIya4VzO
6WgmeSZpjhtO1rGJVimdAT3uRttV6OpJ4YGqpmi8EAWgLZPtUyWB/Pnl2o4h
LAwSvHFC3I8mPccWwHyVYcKrdv8kijaVlKjZ3DN/Zw3AytonjUWbKo/U9n05
xXSxgBNxhp7RGoxGEyt4PmCh2VMBVzRU+z1hGLqZAIfi4S1vVBG91DwF7TwF
4yNbBPsmMf6eYPV5eu0HTbfu7OtnIpPB7/KE21EL8JQ1joyZfrANHx1XVZOn
oEOl7QjK/3AAnnnrW8bhcl1CaVS/cGPW1KqVw5WOzITPVOMAa2CfpT8D6dIY
FXu8dWxgnwtZnxUto9TjYhc3UFmJU+VsnFe0eeq3bOEjmW691l1S08k9vOhk
LyoIi+UZT5kIWNEndI+ihuUODoRVakwLMFfG1nbXmeePeNUTTX2sH/1hQf6T
VdgZFzppw+6bS6vAvxGwz8p5+hsOim+L16BrQnzlzdHSKOVtPZ52dPyT9U+4
vC/hnHr1zAlQadUjizmAEJex/w+F5a+OXRMnp/eVkwQD6hr0eKDXhAZ+nD1K
CCzMWCJrMWNzOx6qlZMQX2Y0ut4tdG6J3zbljsSigWk5WzJUtdwhDNnE213o
BitZDfgoCXjHDPMDFOo8uuqJYgAe9EsC6Lyxl44I+Qj8W5Er1/rnSWMKtq0V
fsdFCboDOy1l2XaVq/YTHTUQuUYfCAxLO6R7xStayWN7hX8L3Pa377lTC6zp
GUUrnRPJUFw5mJYi5BXTaTZ4qykXWITpF3uXkavG5ctvq36NFiApk1ThCTga
TohWLJtcOE+4558C/602t6XqwAFua/pBsqQaPjkEOydk58ki2Nzf+OBZJ+yK
Xe469mJGs6xtNbgXjNOZKJVC1E8360/zLkmK3XW/vKeF9RMIiYLuXUlAkwHi
hdSIQFMz554kLTINKr3aFKUgboC0Fe3oVIRsDpZHhQzEi15qJzpIRO7Xhjka
SMDPlkj1ZHWWDc+F7a6gVhhI46N6iY/DxV/4GLPHvqrakojE5MhrQ/HFSGBW
FlXszCzM2qp32Tjj39nzh1qa8gjNIwtW5EkOsD4RmbgXhQEIGE4wxRzcijzN
p+prGNazyS4lz+wI98mV87qQr6k/jzg1GVhYQbPhJ3x61UDYp42vNGP98K3m
r02hdL+bLnbDtKlP/sG3Qm5j+GWdsRMgG3G4CHQgi6FGuCqgjMNGRkaDnmTv
wfuzftWbMUAnqHi7IF/kHt3qIA99ZKT4agMmEv5Sw2J1jyRFHtG6yuJqkdgV
dUDs6BGWKiAHG1nlWMlA346ae8eI3RPhd3AE0W2f0aitWiiXyw/HgqHYroJB
5kfYTUDEahrS84bSSe4wFEPScUXxPv/Ak7b1ddk2z6t+vVAVWNEpWRlKJ4SH
i5nVPvkzfrADipMUF8Mv4uRiSIKuV0E3/jBt3dikCA3m0qwI7B1qG0W/IiNN
dm7/C761RrEJVSLfxVaz+829XOeWD5dC1ll3LGkr1SxwnwYg8TEIja4gwTJw
DpPpBdPm1FrhktSndnjnbG8P4MK4Lspf2R3dxNOmf1juSU9VbqA45+prRX9c
yTgJf0ebVRFiQYO41BUlM/f3yg+FUun/9BCdUdXeMU/ShIpnGC/9zwO3/GQs
S+LuU9dmLmTZTjKSKiOdVr5NRYQNp6DZHOfz5i2SHsap2ft3EGc+9/qnflq2
cNIqMXNipXDTxXrx8W0HbfKxgWmc5/WBLoWngJ7hFigPkHLNly+YlWZ3CLWA
/wrjHcvKIrD5NjFmp5JvV7obGXPUDFPospTExZpoACnFohJ6M+jhTbr2UZHs
Q2lY/oSwRE6KQKTrrosXjKA3eB07Dmbq/py7jIU2BOd5/6CjBe8BwEhp69gZ
+0u4GDn7PgFJ409zdK+TKLVndCFn8rnEd5mQGWdB9FdZxAFUNiqmkgu8oAvc
q2MS3oe9vtq7JhwQw81VtYUaZ9HpqXJFzjcgJrNv1WY5P5ZijtK5cKbdb/Tl
+OwNhVc2PnOJQNSdZGheBKTv/IKWjL4zPve/T3QPQqFPSnT8iUbK05N/f1jw
N0s=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfTNqB6t6M5ys5ML0ysHOYO8Y7dNIRwNWNy+LobthCphuG2cwf2+fpQIx4Bl0kzdUdBhVwkiEYxXvZyseZPdLG1dP+KNFLQIYFBho8G/vgI1hLvhPri/Sfs0/iZ9mDx9HLwzVB1MigR+lzxiLRT527WYJWlvRsDbyzbFzeqa3sp7KmMNr3NwJgDsw65DyH9I0c/F88dja9z/jcnGLtFiBzr63cXC7ptnEuI1Eh44RHOYpa1Qxebjy790kMALosuyCvH+KYUS3nIG+E9GXeWXIyYsOcGWmgsc47QxS+ludl4PPC+odoSddxMXFYWETj/TWhKnzWNJV3zuaYKxqormOJ/XQI+CZQg9z/TJPSOtxQj7dPTtDLbfBfQ/B16YlHUSASIb2MUJ8/VAwfpxMs7r2GoVBmoo3qN26MzLh8H4liyocK5XGSvMANe1HZL/YC2tP032RYLEfc5/tHx3BUKWxoC6ydueawashKaajEe/ppkWa3lsyA+/Dk6xvP3UjcimaYW1NGdk49YLBv9m0b/woy6dTfgVgRry46R5/3BXzbCnFYOfpAKufGNelPz1O71KDXWhN45mzQw87OArIS+m+q2owppDL9JuIlfFmsGXkW+Anaae/iQFzYBcefvDFEkNRIqNIyUqzd9tJeS3BB/DZPtYW0FkA5tTt/iRr+kby7rvdINDbYn/jQBzqQoRqOp/OBbHSSan+BBoEDS0liGEFCt/Igs1lRoyK5v7fTH7hreYF0oWToKMJLamNa7/H4FGGF3o9dccwbvz3jfCJSR68nZc"
`endif