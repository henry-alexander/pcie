// system_intel_pcie_gts_0_pcie_hal_top_one_lane_pcie_hal_2100_ssolv5i.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_intel_pcie_gts_0_pcie_hal_top_one_lane_pcie_hal_2100_ssolv5i #(
		parameter ch_tx_channel_mode            = "FECD",
		parameter ch_rx_channel_mode            = "PMAD",
		parameter ch_mac_sf_en                  = "DISABLED",
		parameter ch_pldif_sf_en                = "DISABLED",
		parameter ch_pcs_sf_en                  = "DISABLED",
		parameter ch_fec_sf_en                  = "DISABLED",
		parameter ch_SF_PCS_TXMUX_EN            = "ENABLED",
		parameter ch_SF_PCS_RXMUX_EN            = "ENABLED",
		parameter ch_SF_FEC_TXMUX_EN            = "ENABLED",
		parameter ch_SF_FEC_INGRESS_EN          = "ENABLED",
		parameter ch_SF_FEC_EGRESS_EN           = "ENABLED",
		parameter ch_SF_PLDCH_TX_USER1_MUX_EN   = "ENABLED",
		parameter ch_SF_PLDCH_TX_USER2_MUX_EN   = "ENABLED",
		parameter ch_SF_PLDCH_RX_USER1_MUX_EN   = "ENABLED",
		parameter ch_SF_PLDCH_RX_USER2_MUX_EN   = "ENABLED",
		parameter ch_SF_DESKEW_EN               = "ENABLED",
		parameter ch_SF_DESKEW_RXMUX_EN         = "ENABLED",
		parameter ch_SF_PTP_INGRESS_EN          = "ENABLED",
		parameter ch_SF_PTP_EGRESS_EN           = "ENABLED",
		parameter ch_SF_PTP_S_EN                = "ENABLED",
		parameter ch_SF_PTP_EN                  = "ENABLED",
		parameter ch_SF_UX_EN                   = "ENABLED",
		parameter ch_SF_FLUX_GLOBAL_MEM_EN      = "ENABLED",
		parameter ch_SF_FLUX_S_EN               = "ENABLED",
		parameter ch_SF_FLUX_TXUSER_CLK1_MUX_EN = "ENABLED",
		parameter ch_SF_FLUX_TXUSER_CLK2_MUX_EN = "ENABLED",
		parameter ch_SF_FLUX_RXUSER_CLK1_MUX_EN = "ENABLED",
		parameter ch_SF_FLUX_RXUSER_CLK2_MUX_EN = "ENABLED",
		parameter ch_SF_FLUX_I_EN               = "ENABLED",
		parameter ch_SF_UX_TOOLBOX_EN           = "ENABLED",
		parameter ch_SF_FLUX_CORE_EN            = "ENABLED",
		parameter ch_SF_XCVRIF_1CH_EN           = "ENABLED",
		parameter ch_SF_XCVRIF_TXMUX_EN         = "ENABLED",
		parameter ch_SF_XCRIF_TX_RST_MUX_EN     = "ENABLED",
		parameter ch_SF_XCRIF_TX_WREN_MUX_EN    = "ENABLED",
		parameter ch_SF_XCRIF_TX_RDEN_MUX_EN    = "ENABLED",
		parameter ch_SF_XCRIF_TXWORD_CLK_MUX_EN = "ENABLED",
		parameter ch_SF_XCRIF_RXWORD_CLK_MUX_EN = "ENABLED"
	) (
		input  wire [79:0]  i_hio_txdata,                                //                           i_hio_txdata.data,         Stats Snapshot
		input  wire [9:0]   i_hio_txdata_extra,                          //                     i_hio_txdata_extra.data,         RX PFC
		input  wire         i_hio_txdata_fifo_wr_en,                     //                i_hio_txdata_fifo_wr_en.data,         CSR access address
		input  wire         i_hio_rxdata_fifo_rd_en,                     //                i_hio_rxdata_fifo_rd_en.data,         RX error bits asserted on the EOP cycle
		input  wire         i_hio_ptp_rst_n,                             //                        i_hio_ptp_rst_n.reset,        Stats Snapshot
		input  wire         i_hio_ehip_rx_rst_n,                         //                    i_hio_ehip_rx_rst_n.reset,        RX PFC
		input  wire         i_hio_ehip_tx_rst_n,                         //                    i_hio_ehip_tx_rst_n.reset,        CSR access address
		input  wire         i_hio_ehip_signal_ok,                        //                   i_hio_ehip_signal_ok.reset,        RX error bits asserted on the EOP cycle
		input  wire         i_hio_sfreeze_2_r03f_rx_mac_srfz_n,          //     i_hio_sfreeze_2_r03f_rx_mac_srfz_n.reset,        Stats Snapshot
		input  wire         i_hio_sfreeze_3_c2f_tx_deskew_srfz_n,        //   i_hio_sfreeze_3_c2f_tx_deskew_srfz_n.reset,        RX PFC
		input  wire         i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n,          //     i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n.reset,        CSR access address
		input  wire         i_hio_rstfec_fec_rx_rst_n,                   //              i_hio_rstfec_fec_rx_rst_n.reset,        RX error bits asserted on the EOP cycle
		input  wire         i_hio_rstfec_fec_tx_rst_n,                   //              i_hio_rstfec_fec_tx_rst_n.reset,        RX error bits asserted on the EOP cycle
		input  wire         i_hio_rstfec_fec_csr_ret,                    //               i_hio_rstfec_fec_csr_ret.reset,        Stats Snapshot
		input  wire         i_hio_rstfec_rx_fec_sfrz_n,                  //             i_hio_rstfec_rx_fec_sfrz_n.reset,        RX PFC
		input  wire         i_hio_rstfec_tx_fec_sfrz_n,                  //             i_hio_rstfec_tx_fec_sfrz_n.reset,        CSR access address
		input  wire         i_hio_rstxcvrif_xcvrif_rx_rst_n,             //        i_hio_rstxcvrif_xcvrif_rx_rst_n.reset
		input  wire         i_hio_rstxcvrif_xcvrif_tx_rst_n,             //        i_hio_rstxcvrif_xcvrif_tx_rst_n.reset,        Stats Snapshot
		input  wire         i_hio_rstxcvrif_xcvrif_signal_ok,            //       i_hio_rstxcvrif_xcvrif_signal_ok.reset,        RX PFC
		input  wire         i_hio_rstxcvrif_rx_xcvrif_sfrz_n,            //       i_hio_rstxcvrif_rx_xcvrif_sfrz_n.reset,        CSR access address
		input  wire         i_hio_rstxcvrif_tx_xcvrif_sfrz_n,            //       i_hio_rstxcvrif_tx_xcvrif_sfrz_n.reset
		input  wire         i_hio_rst_pld_clrhip,                        //                   i_hio_rst_pld_clrhip.reset,        Stats Snapshot
		input  wire         i_hio_rst_pld_clrpcs,                        //                   i_hio_rst_pld_clrpcs.reset
		input  wire         i_hio_rst_pld_perstn,                        //                   i_hio_rst_pld_perstn.reset,        CSR access address
		input  wire         i_hio_rst_pld_ready,                         //                    i_hio_rst_pld_ready.reset
		input  wire         i_hio_rst_pld_adapter_rx_pld_rst_n,          //     i_hio_rst_pld_adapter_rx_pld_rst_n.reset
		input  wire         i_hio_rst_pld_adapter_tx_pld_rst_n,          //     i_hio_rst_pld_adapter_tx_pld_rst_n.reset
		input  wire         i_hio_rst_ux_rx_pma_rst_n,                   //              i_hio_rst_ux_rx_pma_rst_n.reset
		input  wire         i_hio_rst_ux_rx_sfrz,                        //                   i_hio_rst_ux_rx_sfrz.reset
		input  wire         i_hio_rst_ux_tx_pma_rst_n,                   //              i_hio_rst_ux_tx_pma_rst_n.reset
		input  wire         i_hio_pld_reset_clk_row,                     //                i_hio_pld_reset_clk_row.reset
		input  wire [79:0]  i_hio_uxquad_async,                          //                     i_hio_uxquad_async.data
		input  wire [79:0]  i_hio_uxquad_async_pcie_mux,                 //            i_hio_uxquad_async_pcie_mux.data
		input  wire [20:0]  i_hio_lavmm_addr,                            //                               reconfig.address
		input  wire [3:0]   i_hio_lavmm_be,                              //                                       .byteenable
		input  wire         i_hio_lavmm_read,                            //                                       .read
		input  wire [31:0]  i_hio_lavmm_wdata,                           //                                       .writedata
		input  wire         i_hio_lavmm_write,                           //                                       .write,        RX error bits asserted on the EOP cycle
		output wire [31:0]  o_hio_lavmm_rdata,                           //                                       .readdata
		output wire         o_hio_lavmm_rdata_valid,                     //                                       .readdatavalid
		output wire         o_hio_lavmm_waitreq,                         //                                       .waitrequest
		input  wire         i_hio_lavmm_clk,                             //                           reconfig_clk.clk
		input  wire         i_hio_lavmm_rstn,                            //                           reconfig_rst.reset
		output wire [16:0]  o_ss_lavmm_pcie_addr,                        //                          reconfig_phip.address
		output wire [3:0]   o_ss_lavmm_pcie_be,                          //                                       .byteenable
		output wire         o_ss_lavmm_pcie_read,                        //                                       .read
		output wire [31:0]  o_ss_lavmm_pcie_wdata,                       //                                       .writedata
		output wire         o_ss_lavmm_pcie_write,                       //                                       .write,        RX error bits asserted on the EOP cycle
		input  wire [31:0]  i_ss_lavmm_pcie_rdata,                       //                                       .readdata
		input  wire         i_ss_lavmm_pcie_rdata_valid,                 //                                       .readdatavalid
		input  wire         i_ss_lavmm_pcie_waitreq,                     //                                       .waitrequest
		output wire         o_ss_lavmm_pcie_clk,                         //                      reconfig_clk_phip.clk
		output wire         o_ss_lavmm_pcie_rstn,                        //                      reconfig_rst_phip.reset
		output wire [79:0]  sm_pld_tx_demux_0_o_pcie,                    //               sm_pld_tx_demux_0_o_pcie.data
		input  wire [79:0]  sm_pld_rx_mux_0_i_pcie,                      //                 sm_pld_rx_mux_0_i_pcie.data
		input  wire         o_pld_pcie_clk_4,                            //                       o_pld_pcie_clk_4.clk
		output wire         o_pcie_rxword_clk,                           //                      o_pcie_rxword_clk.clk
		output wire         o_pcie_txword_clk,                           //                      o_pcie_txword_clk.clk
		output wire         ss_rst_ux_rxcdrlock2data,                    //               ss_rst_ux_rxcdrlock2data.data
		output wire [13:0]  o_rxeq_best_eye_vala,                        //                   o_rxeq_best_eye_vala.data
		output wire         o_rxeq_donea,                                //                           o_rxeq_donea.data
		output wire         o_rxmargin_nacka,                            //                       o_rxmargin_nacka.data
		output wire         o_rxmargin_statusa,                          //                     o_rxmargin_statusa.data
		output wire         o_rxsignaldetect_lfpsa,                      //                 o_rxsignaldetect_lfpsa.data
		output wire         o_rxsignaldetecta,                           //                      o_rxsignaldetecta.data
		output wire [1:0]   o_rxmargin_status_gray,                      //                 o_rxmargin_status_gray.data
		output wire         rxstatusa,                                   //                              rxstatusa.data
		output wire [39:0]  o_pcie_pcs,                                  //                             o_pcie_pcs.data
		input  wire [39:0]  i_pcie_pcs,                                  //                             i_pcie_pcs.data
		output wire         o_synthlcfast_postdiv,                       //                  o_synthlcfast_postdiv.data
		output wire         o_synthlcmed_postdiv,                        //                   o_synthlcmed_postdiv.data
		output wire         o_synthlcslow_postdiv,                       //                  o_synthlcslow_postdiv.data
		output wire         o_txdetectrx_acka,                           //                      o_txdetectrx_acka.data
		output wire         o_txdetectrx_statct,                         //                    o_txdetectrx_statct.data
		output wire         txstatusa,                                   //                              txstatusa.data
		input  wire         i_pcs_pipe_rstn,                             //                        i_pcs_pipe_rstn.data
		input  wire         i_ux_ock_pma_clk,                            //                       i_ux_ock_pma_clk.data
		input  wire         i_lfps_ennt,                                 //                            i_lfps_ennt.data
		input  wire [1:0]   i_pcie_l1ctrla,                              //                         i_pcie_l1ctrla.data
		input  wire         i_pma_cmn_ctrl,                              //                         i_pma_cmn_ctrl.data
		input  wire         i_pma_ctrl,                                  //                             i_pma_ctrl.data
		input  wire         i_pcie_pcs_rx_rst,                           //                      i_pcie_pcs_rx_rst.data
		input  wire         i_pcie_pcs_tx_rst,                           //                      i_pcie_pcs_tx_rst.data
		input  wire         i_rxeiosdetectstata,                         //                    i_rxeiosdetectstata.data
		input  wire [2:0]   i_rxeq_precal_code_selnt,                    //               i_rxeq_precal_code_selnt.data
		input  wire         i_rxeq_starta,                               //                          i_rxeq_starta.data
		input  wire         i_rxeq_static_ena,                           //                      i_rxeq_static_ena.data
		input  wire         i_rxmargin_direction_nt,                     //                i_rxmargin_direction_nt.data
		input  wire         i_rxmargin_mode_nt,                          //                     i_rxmargin_mode_nt.data
		input  wire         i_rxmargin_offset_change_a,                  //             i_rxmargin_offset_change_a.data
		input  wire [6:0]   i_rxmargin_offset_nt,                        //                   i_rxmargin_offset_nt.data
		input  wire         i_rxmargin_start_a,                          //                     i_rxmargin_start_a.data
		input  wire [2:0]   i_rxpstate,                                  //                             i_rxpstate.data
		input  wire [3:0]   i_rxrate,                                    //                               i_rxrate.data
		input  wire         i_rxterm_hiz_ena,                            //                       i_rxterm_hiz_ena.data
		input  wire [2:0]   i_rxwidth,                                   //                              i_rxwidth.data
		input  wire         i_tstbus_lane,                               //                          i_tstbus_lane.data
		input  wire         i_txbeacona,                                 //                            i_txbeacona.data
		input  wire [2:0]   i_txclkdivrate,                              //                         i_txclkdivrate.data
		input  wire         i_txdetectrx_reqa,                           //                      i_txdetectrx_reqa.data
		input  wire [5:0]   i_txdrv_levn,                                //                           i_txdrv_levn.data
		input  wire [4:0]   i_txdrv_levnm1,                              //                         i_txdrv_levnm1.data
		input  wire [2:0]   i_txdrv_levnm2,                              //                         i_txdrv_levnm2.data
		input  wire [4:0]   i_txdrv_levnp1,                              //                         i_txdrv_levnp1.data
		input  wire [3:0]   i_txdrv_slew,                                //                           i_txdrv_slew.data
		input  wire [3:0]   i_txelecidle,                                //                           i_txelecidle.data
		input  wire [2:0]   i_txpstate,                                  //                             i_txpstate.data
		input  wire [3:0]   i_txrate,                                    //                               i_txrate.data
		input  wire [2:0]   i_txwidth,                                   //                              i_txwidth.data
		input  wire         i_hio_pld_rx_clk_in_row_clk,                 //            i_hio_pld_rx_clk_in_row_clk.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_pld_tx_clk_in_row_clk,                 //            i_hio_pld_tx_clk_in_row_clk.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_det_lat_rx_dl_clk,                     //                i_hio_det_lat_rx_dl_clk.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_det_lat_rx_mux_select,                 //            i_hio_det_lat_rx_mux_select.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_det_lat_rx_sclk_flop,                  //             i_hio_det_lat_rx_sclk_flop.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_det_lat_rx_sclk_gen_clk,               //          i_hio_det_lat_rx_sclk_gen_clk.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_det_lat_rx_trig_flop,                  //             i_hio_det_lat_rx_trig_flop.clk,          RX error bits asserted on the EOP cycle
		input  wire         i_hio_det_lat_sampling_clk,                  //             i_hio_det_lat_sampling_clk.clk
		input  wire         i_hio_det_lat_tx_dl_clk,                     //                i_hio_det_lat_tx_dl_clk.clk
		input  wire         i_hio_det_lat_tx_mux_select,                 //            i_hio_det_lat_tx_mux_select.clk
		input  wire         i_hio_det_lat_tx_sclk_flop,                  //             i_hio_det_lat_tx_sclk_flop.clk
		input  wire         i_hio_det_lat_tx_sclk_gen_clk,               //          i_hio_det_lat_tx_sclk_gen_clk.clk
		input  wire         i_hio_det_lat_tx_trig_flop,                  //             i_hio_det_lat_tx_trig_flop.clk
		input  wire         rx_serial_n,                                 //                            rx_serial_n.data
		input  wire         rx_serial_p,                                 //                            rx_serial_p.data
		output wire         o_hio_txdata_fifo_wr_empty,                  //             o_hio_txdata_fifo_wr_empty.data
		output wire         o_hio_txdata_fifo_wr_pempty,                 //            o_hio_txdata_fifo_wr_pempty.data
		output wire         o_hio_txdata_fifo_wr_full,                   //              o_hio_txdata_fifo_wr_full.data
		output wire         o_hio_txdata_fifo_wr_pfull,                  //             o_hio_txdata_fifo_wr_pfull.data
		output wire [79:0]  o_hio_rxdata,                                //                           o_hio_rxdata.data
		output wire [9:0]   o_hio_rxdata_extra,                          //                     o_hio_rxdata_extra.data
		output wire         o_hio_rxdata_fifo_rd_empty,                  //             o_hio_rxdata_fifo_rd_empty.data
		output wire         o_hio_rxdata_fifo_rd_pempty,                 //            o_hio_rxdata_fifo_rd_pempty.data
		output wire         o_hio_rxdata_fifo_rd_full,                   //              o_hio_rxdata_fifo_rd_full.data
		output wire         o_hio_rxdata_fifo_rd_pfull,                  //             o_hio_rxdata_fifo_rd_pfull.data
		output wire         o_hio_rstepcs_rx_pcs_fully_aligned,          //     o_hio_rstepcs_rx_pcs_fully_aligned.reset
		output wire         o_hio_rstfec_fec_rx_rdy_n,                   //              o_hio_rstfec_fec_rx_rdy_n.reset
		output wire         o_hio_rst_flux0_cpi_cmn_busy,                //           o_hio_rst_flux0_cpi_cmn_busy.reset
		output wire         o_hio_rst_oflux_rx_srds_rdy,                 //            o_hio_rst_oflux_rx_srds_rdy.reset
		output wire         o_hio_rst_ux_all_synthlockstatus,            //       o_hio_rst_ux_all_synthlockstatus.reset
		output wire         o_hio_rst_ux_octl_pcs_rxstatus,              //         o_hio_rst_ux_octl_pcs_rxstatus.reset
		output wire         o_hio_rst_ux_octl_pcs_txstatus,              //         o_hio_rst_ux_octl_pcs_txstatus.reset
		output wire         o_hio_rst_ux_rxcdrlock2data,                 //            o_hio_rst_ux_rxcdrlock2data.reset
		output wire         o_hio_rst_ux_rxcdrlockstatus,                //           o_hio_rst_ux_rxcdrlockstatus.reset
		output wire [49:0]  o_hio_uxquad_async,                          //                     o_hio_uxquad_async.data
		output wire         o_hio_user_rx_clk1_clk,                      //                 o_hio_user_rx_clk1_clk.clk
		output wire         o_hio_user_rx_clk2_clk,                      //                 o_hio_user_rx_clk2_clk.clk
		output wire         o_hio_user_tx_clk1_clk,                      //                 o_hio_user_tx_clk1_clk.clk
		output wire         o_hio_user_tx_clk2_clk,                      //                 o_hio_user_tx_clk2_clk.clk
		output wire         o_hio_ux_chnl_refclk_mux,                    //               o_hio_ux_chnl_refclk_mux.clk
		output wire         o_hio_det_lat_rx_async_dl_sync,              //         o_hio_det_lat_rx_async_dl_sync.clk
		output wire         o_hio_det_lat_rx_async_pulse,                //           o_hio_det_lat_rx_async_pulse.clk
		output wire         o_hio_det_lat_rx_async_sample_sync,          //     o_hio_det_lat_rx_async_sample_sync.clk
		output wire         o_hio_det_lat_rx_sclk_sample_sync,           //      o_hio_det_lat_rx_sclk_sample_sync.clk
		output wire         o_hio_det_lat_rx_trig_sample_sync,           //      o_hio_det_lat_rx_trig_sample_sync.clk
		output wire         o_hio_det_lat_tx_async_dl_sync,              //         o_hio_det_lat_tx_async_dl_sync.clk
		output wire         o_hio_det_lat_tx_async_pulse,                //           o_hio_det_lat_tx_async_pulse.clk
		output wire         o_hio_det_lat_tx_async_sample_sync,          //     o_hio_det_lat_tx_async_sample_sync.clk
		output wire         o_hio_det_lat_tx_sclk_sample_sync,           //      o_hio_det_lat_tx_sclk_sample_sync.clk
		output wire         o_hio_det_lat_tx_trig_sample_sync,           //      o_hio_det_lat_tx_trig_sample_sync.clk
		output wire         o_hio_xcvrif_rx_latency_pulse,               //          o_hio_xcvrif_rx_latency_pulse.clk
		output wire         o_hio_xcvrif_tx_latency_pulse,               //          o_hio_xcvrif_tx_latency_pulse.clk
		output wire         tx_serial_p,                                 //                            tx_serial_p.data
		output wire         tx_serial_n,                                 //                            tx_serial_n.data
		input  wire [99:0]  i_hio_txdata_async,                          //                     i_hio_txdata_async.data
		input  wire [9:0]   i_hio_txdata_direct,                         //                    i_hio_txdata_direct.data
		output wire [99:0]  o_hio_rxdata_async,                          //                     o_hio_rxdata_async.data
		output wire [9:0]   o_hio_rxdata_direct,                         //                    o_hio_rxdata_direct.data
		input  wire [767:0] i_uxwrap_bus_in_phy_shared,                  //                          uxwrap_bus_in.data
		output wire [703:0] o_uxwrap_bus_out_phy_shared,                 //                         uxwrap_bus_out.data
		output wire [19:0]  o_lavmm_addr_phy_shared,                     //                    reconfig_phy_shared.address
		output wire [3:0]   o_lavmm_be_phy_shared,                       //                                       .byteenable
		output wire         o_lavmm_read_phy_shared,                     //                                       .read
		output wire [31:0]  o_lavmm_wdata_phy_shared,                    //                                       .writedata
		output wire         o_lavmm_write_phy_shared,                    //                                       .write
		input  wire [31:0]  i_lavmm_rdata_phy_shared,                    //                                       .readdata
		input  wire         i_lavmm_rdata_valid_phy_shared,              //                                       .readdatavalid
		input  wire         i_lavmm_waitreq_phy_shared,                  //                                       .waitrequest
		output wire         o_lavmm_clk_phy_shared,                      //                reconfig_clk_phy_shared.clk
		output wire         o_lavmm_rstn_phy_shared,                     //                reconfig_rst_phy_shared.reset
		output wire         o_sclk_return_sel_rx_phy_shared,             //                   o_sclk_return_sel_rx.data
		output wire         o_sclk_return_sel_tx_phy_shared,             //                   o_sclk_return_sel_tx.data
		output wire         o_ick_sclk_rx_phy_shared,                    //                          o_ick_sclk_rx.clk
		input  wire [4:0]   i_sync_common_control_phy_shared,            //                  i_sync_common_control.data
		output wire         o_ft_rx_sclk_sync_ch_phy_shared,             //                   o_ft_rx_sclk_sync_ch.data
		output wire         o_ft_tx_sclk_sync_ch_phy_shared,             //                   o_ft_tx_sclk_sync_ch.data
		output wire         o_rst_ux_rx_pma_rst_n_phy_shared,            //                  o_rst_ux_rx_pma_rst_n.reset
		output wire         o_rst_ux_tx_pma_rst_n_phy_shared,            //                  o_rst_ux_tx_pma_rst_n.reset
		output wire         o_ick_pcs_txword_phy_shared,                 //                       o_ick_pcs_txword.data
		output wire         o_tx_dl_ch_bit_phy_shared,                   //                         o_tx_dl_ch_bit.data
		input  wire         i_dat_pcs_measlatbit_phy_shared,             //                   i_dat_pcs_measlatbit.data
		input  wire         i_ft_rx_async_pulse_ch_phy_shared,           //                 i_ft_rx_async_pulse_ch.data
		input  wire         i_ft_tx_async_pulse_ch_phy_shared,           //                 i_ft_tx_async_pulse_ch.data
		input  wire         i_rx_dl_ch_bit_phy_shared,                   //                         i_rx_dl_ch_bit.data
		input  wire [1:0]   i_ux_rxuser1_sel_phy_shared,                 //                       i_ux_rxuser1_sel.data
		input  wire [1:0]   i_ux_rxuser2_sel_phy_shared,                 //                       i_ux_rxuser2_sel.data
		input  wire [1:0]   i_ux_txuser1_sel_phy_shared,                 //                       i_ux_txuser1_sel.data
		input  wire [1:0]   i_ux_txuser2_sel_phy_shared,                 //                       i_ux_txuser2_sel.data
		output wire         o_octl_pcs_txstatus_a_phy_shared,            //                  o_octl_pcs_txstatus_a.data
		input  wire         i_ictl_pcs_txenable_a_phy_shared,            //                  i_ictl_pcs_txenable_a.data
		input  wire [124:0] i_sync_cfg_data_phy_shared,                  //                        i_sync_cfg_data.data
		input  wire [249:0] i_sync_interface_control_phy_shared,         //               i_sync_interface_control.data
		output wire [79:0]  o_tx_data_phy_shared,                        //                              o_tx_data.data
		input  wire [79:0]  i_rx_data_phy_shared,                        //                              i_rx_data.data
		output wire [319:0] o_sm_flux_ingress_phy_shared,                //                      o_sm_flux_ingress.data
		input  wire [256:0] i_sm_flux_egress_phy_shared,                 //                       i_sm_flux_egress.data
		input  wire         i_flux_cpi_int_phy_shared,                   //                         i_flux_cpi_int.data
		input  wire         i_flux_int_phy_shared,                       //                             i_flux_int.data
		input  wire         i_oflux_octl_pcs_txptr_smpl_lane_phy_shared, //       i_oflux_octl_pcs_txptr_smpl_lane.data
		output wire         o_ick_sclk_tx_phy_shared,                    //                          o_ick_sclk_tx.clk
		input  wire         i_flux_srds_rdy_phy_shared,                  //                        i_flux_srds_rdy.data
		input  wire         i_pcs_rxword_phy_shared,                     //                           i_pcs_rxword.data
		input  wire         i_pcs_rxpostdiv_phy_shared,                  //                        i_pcs_rxpostdiv.data
		input  wire         i_ock_pcs_txword_phy_shared,                 //                       i_ock_pcs_txword.data
		output wire         o_dat_pcs_measlatrndtripbit_phy_shared,      // o_dat_pcs_measlatrndtripbit_phy_shared.data
		input  wire [11:0]  i_ch_eth_fec_rx_async_fec_wrap,              //                            asyncdata_4.data
		input  wire         i_ch_eth_fec_rx_direct_fec_wrap,             //                            asyncdata_5.data
		input  wire         i_fec_rx_rdy_n_fec_wrap,                     //                i_fec_rx_rdy_n_fec_wrap.data
		input  wire         i_fec_tx_data_mux_sel_fec_wrap,              //         i_fec_tx_data_mux_sel_fec_wrap.muxsel
		input  wire [42:0]  i_fec_rx_data_fec_wrap,                      //                 i_fec_rx_data_fec_wrap.data
		input  wire [42:0]  i_xcvr_tx_data,                              //                         i_xcvr_tx_data.data
		output wire         ss_rst_flux0_cpi_cmn_busy,                   //              ss_rst_flux0_cpi_cmn_busy.data
		output wire         o_pma_rx_sf,                                 //                            o_pma_rx_sf.data
		input  wire         i_refclk_tx_p,                               //                          i_refclk_tx_p.clk
		input  wire         i_syspll_c0_clk,                             //                        i_syspll_c0_clk.clk
		input  wire         i_syspll_c1_clk,                             //                        i_syspll_c1_clk.clk
		input  wire         i_syspll_c2_clk,                             //                        i_syspll_c2_clk.clk
		input  wire         i_flux_clk,                                  //                             i_flux_clk.clk
		input  wire         i_refclk_rx_p,                               //                          i_refclk_rx_p.clk
		input  wire         i_ux_chnl_refclk_mux_phy_shared,             //        i_ux_chnl_refclk_mux_phy_shared.clk
		output wire         o_xcvrif_tx_fifo_rd_en_mux_x1,               //          o_xcvrif_tx_fifo_rd_en_mux_x1.clk
		input  wire         i_xcvrif_tx_fifo_rd_en_mux_x2,               //          i_xcvrif_tx_fifo_rd_en_mux_x2.clk
		input  wire         i_xcvrif_tx_fifo_rd_en_mux_x4,               //          i_xcvrif_tx_fifo_rd_en_mux_x4.clk
		input  wire         i_xcvrif_tx_fifo_rd_en_mux_x6_bot,           //      i_xcvrif_tx_fifo_rd_en_mux_x6_bot.clk
		input  wire         i_xcvrif_tx_fifo_rd_en_mux_x6_top,           //      i_xcvrif_tx_fifo_rd_en_mux_x6_top.clk
		input  wire         i_xcvrif_tx_fifo_rd_en_mux_x8_bot,           //      i_xcvrif_tx_fifo_rd_en_mux_x8_bot.clk
		input  wire         i_xcvrif_tx_fifo_rd_en_mux_x8_top,           //      i_xcvrif_tx_fifo_rd_en_mux_x8_top.clk
		output wire         o_xcvrif_tx_rst_mux_x1,                      //                 o_xcvrif_tx_rst_mux_x1.clk
		input  wire         i_xcvrif_tx_rst_mux_x2,                      //                 i_xcvrif_tx_rst_mux_x2.clk
		input  wire         i_xcvrif_tx_rst_mux_x4,                      //                 i_xcvrif_tx_rst_mux_x4.clk
		input  wire         i_xcvrif_tx_rst_mux_x6_bot,                  //             i_xcvrif_tx_rst_mux_x6_bot.clk
		input  wire         i_xcvrif_tx_rst_mux_x6_top,                  //             i_xcvrif_tx_rst_mux_x6_top.clk
		input  wire         i_xcvrif_tx_rst_mux_x8_bot,                  //             i_xcvrif_tx_rst_mux_x8_bot.clk
		input  wire         i_xcvrif_tx_rst_mux_x8_top,                  //             i_xcvrif_tx_rst_mux_x8_top.clk
		output wire         o_xcvrif_tx_word_clk_mux_x1,                 //            o_xcvrif_tx_word_clk_mux_x1.clk
		input  wire         i_xcvrif_tx_word_clk_mux_x2,                 //            i_xcvrif_tx_word_clk_mux_x2.clk
		input  wire         i_xcvrif_tx_word_clk_mux_x4,                 //            i_xcvrif_tx_word_clk_mux_x4.clk
		input  wire         i_xcvrif_tx_word_clk_mux_x6_bot,             //        i_xcvrif_tx_word_clk_mux_x6_bot.clk
		input  wire         i_xcvrif_tx_word_clk_mux_x6_top,             //        i_xcvrif_tx_word_clk_mux_x6_top.clk
		input  wire         i_xcvrif_tx_word_clk_mux_x8_bot,             //        i_xcvrif_tx_word_clk_mux_x8_bot.clk
		input  wire         i_xcvrif_tx_word_clk_mux_x8_top,             //        i_xcvrif_tx_word_clk_mux_x8_top.clk
		input  wire         ioack_cdrdiv_left_ux_bidir_in,               //          ioack_cdrdiv_left_ux_bidir_in.clk
		input  wire         ioack_synthdiv1_left_ux_bidir_in,            //       ioack_synthdiv1_left_ux_bidir_in.clk
		input  wire         ioack_synthdiv2_left_ux_bidir_in,            //       ioack_synthdiv2_left_ux_bidir_in.clk
		output wire         ioack_cdrdiv_left_ux_bidir_out,              //         ioack_cdrdiv_left_ux_bidir_out.clk
		output wire         ioack_synthdiv1_left_ux_bidir_out,           //      ioack_synthdiv1_left_ux_bidir_out.clk
		output wire         ioack_synthdiv2_left_ux_bidir_out,           //      ioack_synthdiv2_left_ux_bidir_out.clk
		output wire         o_xcvrif_tx_rst_wr_sync_mux_x1,              //         o_xcvrif_tx_rst_wr_sync_mux_x1.clk
		input  wire         i_xcvrif_tx_rst_wr_sync_mux_x2,              //         i_xcvrif_tx_rst_wr_sync_mux_x2.clk
		input  wire         i_xcvrif_tx_rst_wr_sync_mux_x4,              //         i_xcvrif_tx_rst_wr_sync_mux_x4.clk
		input  wire         i_xcvrif_tx_rst_wr_sync_mux_x6_bot,          //     i_xcvrif_tx_rst_wr_sync_mux_x6_bot.clk
		input  wire         i_xcvrif_tx_rst_wr_sync_mux_x6_top,          //     i_xcvrif_tx_rst_wr_sync_mux_x6_top.clk
		input  wire         i_xcvrif_tx_rst_wr_sync_mux_x8_bot,          //     i_xcvrif_tx_rst_wr_sync_mux_x8_bot.clk
		input  wire         i_xcvrif_tx_rst_wr_sync_mux_x8_top,          //     i_xcvrif_tx_rst_wr_sync_mux_x8_top.clk
		output wire         ss_user_rx_clk1_clk,                         //                    ss_user_rx_clk1_clk.clk
		output wire         ss_user_rx_clk2_clk,                         //                    ss_user_rx_clk2_clk.clk
		output wire         ss_user_tx_clk1_clk,                         //                    ss_user_tx_clk1_clk.clk
		output wire         ss_user_tx_clk2_clk,                         //                    ss_user_tx_clk2_clk.clk
		output wire         ss_user_rx_clk1_clk_w,                       //                  ss_user_rx_clk1_clk_w.clk
		output wire         ss_user_rx_clk2_clk_w,                       //                  ss_user_rx_clk2_clk_w.clk
		output wire         ss_user_tx_clk1_clk_w,                       //                  ss_user_tx_clk1_clk_w.clk
		output wire         ss_user_tx_clk2_clk_w,                       //                  ss_user_tx_clk2_clk_w.clk
		output wire         o_hio_ux_tx_ch_ptr_smpl                      //                o_hio_ux_tx_ch_ptr_smpl.data
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (ch_tx_channel_mode != "FECD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_tx_channel_mode_check ( .error(1'b1) );
		end
		if (ch_rx_channel_mode != "PMAD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_rx_channel_mode_check ( .error(1'b1) );
		end
		if (ch_mac_sf_en != "DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_mac_sf_en_check ( .error(1'b1) );
		end
		if (ch_pldif_sf_en != "DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_sf_en_check ( .error(1'b1) );
		end
		if (ch_pcs_sf_en != "DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pcs_sf_en_check ( .error(1'b1) );
		end
		if (ch_fec_sf_en != "DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_fec_sf_en_check ( .error(1'b1) );
		end
		if (ch_SF_PCS_TXMUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_pcs_txmux_en_check ( .error(1'b1) );
		end
		if (ch_SF_PCS_RXMUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_pcs_rxmux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FEC_TXMUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_fec_txmux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FEC_INGRESS_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_fec_ingress_en_check ( .error(1'b1) );
		end
		if (ch_SF_FEC_EGRESS_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_fec_egress_en_check ( .error(1'b1) );
		end
		if (ch_SF_PLDCH_TX_USER1_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_pldch_tx_user1_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_PLDCH_TX_USER2_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_pldch_tx_user2_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_PLDCH_RX_USER1_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_pldch_rx_user1_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_PLDCH_RX_USER2_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_pldch_rx_user2_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_DESKEW_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_deskew_en_check ( .error(1'b1) );
		end
		if (ch_SF_DESKEW_RXMUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_deskew_rxmux_en_check ( .error(1'b1) );
		end
		if (ch_SF_PTP_INGRESS_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_ptp_ingress_en_check ( .error(1'b1) );
		end
		if (ch_SF_PTP_EGRESS_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_ptp_egress_en_check ( .error(1'b1) );
		end
		if (ch_SF_PTP_S_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_ptp_s_en_check ( .error(1'b1) );
		end
		if (ch_SF_PTP_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_ptp_en_check ( .error(1'b1) );
		end
		if (ch_SF_UX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_ux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_GLOBAL_MEM_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_global_mem_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_S_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_s_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_TXUSER_CLK1_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_txuser_clk1_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_TXUSER_CLK2_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_txuser_clk2_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_RXUSER_CLK1_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_rxuser_clk1_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_RXUSER_CLK2_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_rxuser_clk2_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_I_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_i_en_check ( .error(1'b1) );
		end
		if (ch_SF_UX_TOOLBOX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_ux_toolbox_en_check ( .error(1'b1) );
		end
		if (ch_SF_FLUX_CORE_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_flux_core_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCVRIF_1CH_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcvrif_1ch_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCVRIF_TXMUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcvrif_txmux_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCRIF_TX_RST_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcrif_tx_rst_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCRIF_TX_WREN_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcrif_tx_wren_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCRIF_TX_RDEN_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcrif_tx_rden_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCRIF_TXWORD_CLK_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcrif_txword_clk_mux_en_check ( .error(1'b1) );
		end
		if (ch_SF_XCRIF_RXWORD_CLK_MUX_EN != "ENABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_sf_xcrif_rxword_clk_mux_en_check ( .error(1'b1) );
		end
	endgenerate

	system_intel_pcie_gts_0_one_lane_pcie_hal_2100_5iub4oy #(
		.ch_tx_channel_mode            ("FECD"),
		.ch_rx_channel_mode            ("PMAD"),
		.ch_mac_sf_en                  ("DISABLED"),
		.ch_pldif_sf_en                ("DISABLED"),
		.ch_pcs_sf_en                  ("DISABLED"),
		.ch_fec_sf_en                  ("DISABLED"),
		.ch_SF_PCS_TXMUX_EN            ("ENABLED"),
		.ch_SF_PCS_RXMUX_EN            ("ENABLED"),
		.ch_SF_FEC_TXMUX_EN            ("ENABLED"),
		.ch_SF_FEC_INGRESS_EN          ("ENABLED"),
		.ch_SF_FEC_EGRESS_EN           ("ENABLED"),
		.ch_SF_PLDCH_TX_USER1_MUX_EN   ("ENABLED"),
		.ch_SF_PLDCH_TX_USER2_MUX_EN   ("ENABLED"),
		.ch_SF_PLDCH_RX_USER1_MUX_EN   ("ENABLED"),
		.ch_SF_PLDCH_RX_USER2_MUX_EN   ("ENABLED"),
		.ch_SF_DESKEW_EN               ("ENABLED"),
		.ch_SF_DESKEW_RXMUX_EN         ("ENABLED"),
		.ch_SF_PTP_INGRESS_EN          ("ENABLED"),
		.ch_SF_PTP_EGRESS_EN           ("ENABLED"),
		.ch_SF_PTP_S_EN                ("ENABLED"),
		.ch_SF_PTP_EN                  ("ENABLED"),
		.ch_SF_UX_EN                   ("ENABLED"),
		.ch_SF_FLUX_GLOBAL_MEM_EN      ("ENABLED"),
		.ch_SF_FLUX_S_EN               ("ENABLED"),
		.ch_SF_FLUX_TXUSER_CLK1_MUX_EN ("ENABLED"),
		.ch_SF_FLUX_TXUSER_CLK2_MUX_EN ("ENABLED"),
		.ch_SF_FLUX_RXUSER_CLK1_MUX_EN ("ENABLED"),
		.ch_SF_FLUX_RXUSER_CLK2_MUX_EN ("ENABLED"),
		.ch_SF_FLUX_I_EN               ("ENABLED"),
		.ch_SF_UX_TOOLBOX_EN           ("ENABLED"),
		.ch_SF_FLUX_CORE_EN            ("ENABLED"),
		.ch_SF_XCVRIF_1CH_EN           ("ENABLED"),
		.ch_SF_XCVRIF_TXMUX_EN         ("ENABLED"),
		.ch_SF_XCRIF_TX_RST_MUX_EN     ("ENABLED"),
		.ch_SF_XCRIF_TX_WREN_MUX_EN    ("ENABLED"),
		.ch_SF_XCRIF_TX_RDEN_MUX_EN    ("ENABLED"),
		.ch_SF_XCRIF_TXWORD_CLK_MUX_EN ("ENABLED"),
		.ch_SF_XCRIF_RXWORD_CLK_MUX_EN ("ENABLED")
	) one_lane_pcie_hal_top_p1 (
		.i_hio_txdata                                (i_hio_txdata),                                //   input,   width = 80,                           i_hio_txdata.data
		.i_hio_txdata_extra                          (i_hio_txdata_extra),                          //   input,   width = 10,                     i_hio_txdata_extra.data
		.i_hio_txdata_fifo_wr_en                     (i_hio_txdata_fifo_wr_en),                     //   input,    width = 1,                i_hio_txdata_fifo_wr_en.data
		.i_hio_rxdata_fifo_rd_en                     (i_hio_rxdata_fifo_rd_en),                     //   input,    width = 1,                i_hio_rxdata_fifo_rd_en.data
		.i_hio_ptp_rst_n                             (i_hio_ptp_rst_n),                             //   input,    width = 1,                        i_hio_ptp_rst_n.reset
		.i_hio_ehip_rx_rst_n                         (i_hio_ehip_rx_rst_n),                         //   input,    width = 1,                    i_hio_ehip_rx_rst_n.reset
		.i_hio_ehip_tx_rst_n                         (i_hio_ehip_tx_rst_n),                         //   input,    width = 1,                    i_hio_ehip_tx_rst_n.reset
		.i_hio_ehip_signal_ok                        (i_hio_ehip_signal_ok),                        //   input,    width = 1,                   i_hio_ehip_signal_ok.reset
		.i_hio_sfreeze_2_r03f_rx_mac_srfz_n          (i_hio_sfreeze_2_r03f_rx_mac_srfz_n),          //   input,    width = 1,     i_hio_sfreeze_2_r03f_rx_mac_srfz_n.reset
		.i_hio_sfreeze_3_c2f_tx_deskew_srfz_n        (i_hio_sfreeze_3_c2f_tx_deskew_srfz_n),        //   input,    width = 1,   i_hio_sfreeze_3_c2f_tx_deskew_srfz_n.reset
		.i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n          (i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n),          //   input,    width = 1,     i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n.reset
		.i_hio_rstfec_fec_rx_rst_n                   (i_hio_rstfec_fec_rx_rst_n),                   //   input,    width = 1,              i_hio_rstfec_fec_rx_rst_n.reset
		.i_hio_rstfec_fec_tx_rst_n                   (i_hio_rstfec_fec_tx_rst_n),                   //   input,    width = 1,              i_hio_rstfec_fec_tx_rst_n.reset
		.i_hio_rstfec_fec_csr_ret                    (i_hio_rstfec_fec_csr_ret),                    //   input,    width = 1,               i_hio_rstfec_fec_csr_ret.reset
		.i_hio_rstfec_rx_fec_sfrz_n                  (i_hio_rstfec_rx_fec_sfrz_n),                  //   input,    width = 1,             i_hio_rstfec_rx_fec_sfrz_n.reset
		.i_hio_rstfec_tx_fec_sfrz_n                  (i_hio_rstfec_tx_fec_sfrz_n),                  //   input,    width = 1,             i_hio_rstfec_tx_fec_sfrz_n.reset
		.i_hio_rstxcvrif_xcvrif_rx_rst_n             (i_hio_rstxcvrif_xcvrif_rx_rst_n),             //   input,    width = 1,        i_hio_rstxcvrif_xcvrif_rx_rst_n.reset
		.i_hio_rstxcvrif_xcvrif_tx_rst_n             (i_hio_rstxcvrif_xcvrif_tx_rst_n),             //   input,    width = 1,        i_hio_rstxcvrif_xcvrif_tx_rst_n.reset
		.i_hio_rstxcvrif_xcvrif_signal_ok            (i_hio_rstxcvrif_xcvrif_signal_ok),            //   input,    width = 1,       i_hio_rstxcvrif_xcvrif_signal_ok.reset
		.i_hio_rstxcvrif_rx_xcvrif_sfrz_n            (i_hio_rstxcvrif_rx_xcvrif_sfrz_n),            //   input,    width = 1,       i_hio_rstxcvrif_rx_xcvrif_sfrz_n.reset
		.i_hio_rstxcvrif_tx_xcvrif_sfrz_n            (i_hio_rstxcvrif_tx_xcvrif_sfrz_n),            //   input,    width = 1,       i_hio_rstxcvrif_tx_xcvrif_sfrz_n.reset
		.i_hio_rst_pld_clrhip                        (i_hio_rst_pld_clrhip),                        //   input,    width = 1,                   i_hio_rst_pld_clrhip.reset
		.i_hio_rst_pld_clrpcs                        (i_hio_rst_pld_clrpcs),                        //   input,    width = 1,                   i_hio_rst_pld_clrpcs.reset
		.i_hio_rst_pld_perstn                        (i_hio_rst_pld_perstn),                        //   input,    width = 1,                   i_hio_rst_pld_perstn.reset
		.i_hio_rst_pld_ready                         (i_hio_rst_pld_ready),                         //   input,    width = 1,                    i_hio_rst_pld_ready.reset
		.i_hio_rst_pld_adapter_rx_pld_rst_n          (i_hio_rst_pld_adapter_rx_pld_rst_n),          //   input,    width = 1,     i_hio_rst_pld_adapter_rx_pld_rst_n.reset
		.i_hio_rst_pld_adapter_tx_pld_rst_n          (i_hio_rst_pld_adapter_tx_pld_rst_n),          //   input,    width = 1,     i_hio_rst_pld_adapter_tx_pld_rst_n.reset
		.i_hio_rst_ux_rx_pma_rst_n                   (i_hio_rst_ux_rx_pma_rst_n),                   //   input,    width = 1,              i_hio_rst_ux_rx_pma_rst_n.reset
		.i_hio_rst_ux_rx_sfrz                        (i_hio_rst_ux_rx_sfrz),                        //   input,    width = 1,                   i_hio_rst_ux_rx_sfrz.reset
		.i_hio_rst_ux_tx_pma_rst_n                   (i_hio_rst_ux_tx_pma_rst_n),                   //   input,    width = 1,              i_hio_rst_ux_tx_pma_rst_n.reset
		.i_hio_pld_reset_clk_row                     (i_hio_pld_reset_clk_row),                     //   input,    width = 1,                i_hio_pld_reset_clk_row.reset
		.i_hio_uxquad_async                          (i_hio_uxquad_async),                          //   input,   width = 80,                     i_hio_uxquad_async.data
		.i_hio_uxquad_async_pcie_mux                 (i_hio_uxquad_async_pcie_mux),                 //   input,   width = 80,            i_hio_uxquad_async_pcie_mux.data
		.i_hio_lavmm_addr                            (i_hio_lavmm_addr),                            //   input,   width = 21,                               reconfig.address
		.i_hio_lavmm_be                              (i_hio_lavmm_be),                              //   input,    width = 4,                                       .byteenable
		.i_hio_lavmm_read                            (i_hio_lavmm_read),                            //   input,    width = 1,                                       .read
		.i_hio_lavmm_wdata                           (i_hio_lavmm_wdata),                           //   input,   width = 32,                                       .writedata
		.i_hio_lavmm_write                           (i_hio_lavmm_write),                           //   input,    width = 1,                                       .write
		.o_hio_lavmm_rdata                           (o_hio_lavmm_rdata),                           //  output,   width = 32,                                       .readdata
		.o_hio_lavmm_rdata_valid                     (o_hio_lavmm_rdata_valid),                     //  output,    width = 1,                                       .readdatavalid
		.o_hio_lavmm_waitreq                         (o_hio_lavmm_waitreq),                         //  output,    width = 1,                                       .waitrequest
		.i_hio_lavmm_clk                             (i_hio_lavmm_clk),                             //   input,    width = 1,                           reconfig_clk.clk
		.i_hio_lavmm_rstn                            (i_hio_lavmm_rstn),                            //   input,    width = 1,                           reconfig_rst.reset
		.o_ss_lavmm_pcie_addr                        (o_ss_lavmm_pcie_addr),                        //  output,   width = 17,                          reconfig_phip.address
		.o_ss_lavmm_pcie_be                          (o_ss_lavmm_pcie_be),                          //  output,    width = 4,                                       .byteenable
		.o_ss_lavmm_pcie_read                        (o_ss_lavmm_pcie_read),                        //  output,    width = 1,                                       .read
		.o_ss_lavmm_pcie_wdata                       (o_ss_lavmm_pcie_wdata),                       //  output,   width = 32,                                       .writedata
		.o_ss_lavmm_pcie_write                       (o_ss_lavmm_pcie_write),                       //  output,    width = 1,                                       .write
		.i_ss_lavmm_pcie_rdata                       (i_ss_lavmm_pcie_rdata),                       //   input,   width = 32,                                       .readdata
		.i_ss_lavmm_pcie_rdata_valid                 (i_ss_lavmm_pcie_rdata_valid),                 //   input,    width = 1,                                       .readdatavalid
		.i_ss_lavmm_pcie_waitreq                     (i_ss_lavmm_pcie_waitreq),                     //   input,    width = 1,                                       .waitrequest
		.o_ss_lavmm_pcie_clk                         (o_ss_lavmm_pcie_clk),                         //  output,    width = 1,                      reconfig_clk_phip.clk
		.o_ss_lavmm_pcie_rstn                        (o_ss_lavmm_pcie_rstn),                        //  output,    width = 1,                      reconfig_rst_phip.reset
		.sm_pld_tx_demux_0_o_pcie                    (sm_pld_tx_demux_0_o_pcie),                    //  output,   width = 80,               sm_pld_tx_demux_0_o_pcie.data
		.sm_pld_rx_mux_0_i_pcie                      (sm_pld_rx_mux_0_i_pcie),                      //   input,   width = 80,                 sm_pld_rx_mux_0_i_pcie.data
		.o_pld_pcie_clk_4                            (o_pld_pcie_clk_4),                            //   input,    width = 1,                       o_pld_pcie_clk_4.clk
		.o_pcie_rxword_clk                           (o_pcie_rxword_clk),                           //  output,    width = 1,                      o_pcie_rxword_clk.clk
		.o_pcie_txword_clk                           (o_pcie_txword_clk),                           //  output,    width = 1,                      o_pcie_txword_clk.clk
		.ss_rst_ux_rxcdrlock2data                    (ss_rst_ux_rxcdrlock2data),                    //  output,    width = 1,               ss_rst_ux_rxcdrlock2data.data
		.o_rxeq_best_eye_vala                        (o_rxeq_best_eye_vala),                        //  output,   width = 14,                   o_rxeq_best_eye_vala.data
		.o_rxeq_donea                                (o_rxeq_donea),                                //  output,    width = 1,                           o_rxeq_donea.data
		.o_rxmargin_nacka                            (o_rxmargin_nacka),                            //  output,    width = 1,                       o_rxmargin_nacka.data
		.o_rxmargin_statusa                          (o_rxmargin_statusa),                          //  output,    width = 1,                     o_rxmargin_statusa.data
		.o_rxsignaldetect_lfpsa                      (o_rxsignaldetect_lfpsa),                      //  output,    width = 1,                 o_rxsignaldetect_lfpsa.data
		.o_rxsignaldetecta                           (o_rxsignaldetecta),                           //  output,    width = 1,                      o_rxsignaldetecta.data
		.o_rxmargin_status_gray                      (o_rxmargin_status_gray),                      //  output,    width = 2,                 o_rxmargin_status_gray.data
		.rxstatusa                                   (rxstatusa),                                   //  output,    width = 1,                              rxstatusa.data
		.o_pcie_pcs                                  (o_pcie_pcs),                                  //  output,   width = 40,                             o_pcie_pcs.data
		.i_pcie_pcs                                  (i_pcie_pcs),                                  //   input,   width = 40,                             i_pcie_pcs.data
		.o_synthlcfast_postdiv                       (o_synthlcfast_postdiv),                       //  output,    width = 1,                  o_synthlcfast_postdiv.data
		.o_synthlcmed_postdiv                        (o_synthlcmed_postdiv),                        //  output,    width = 1,                   o_synthlcmed_postdiv.data
		.o_synthlcslow_postdiv                       (o_synthlcslow_postdiv),                       //  output,    width = 1,                  o_synthlcslow_postdiv.data
		.o_txdetectrx_acka                           (o_txdetectrx_acka),                           //  output,    width = 1,                      o_txdetectrx_acka.data
		.o_txdetectrx_statct                         (o_txdetectrx_statct),                         //  output,    width = 1,                    o_txdetectrx_statct.data
		.txstatusa                                   (txstatusa),                                   //  output,    width = 1,                              txstatusa.data
		.i_pcs_pipe_rstn                             (i_pcs_pipe_rstn),                             //   input,    width = 1,                        i_pcs_pipe_rstn.data
		.i_ux_ock_pma_clk                            (i_ux_ock_pma_clk),                            //   input,    width = 1,                       i_ux_ock_pma_clk.data
		.i_lfps_ennt                                 (i_lfps_ennt),                                 //   input,    width = 1,                            i_lfps_ennt.data
		.i_pcie_l1ctrla                              (i_pcie_l1ctrla),                              //   input,    width = 2,                         i_pcie_l1ctrla.data
		.i_pma_cmn_ctrl                              (i_pma_cmn_ctrl),                              //   input,    width = 1,                         i_pma_cmn_ctrl.data
		.i_pma_ctrl                                  (i_pma_ctrl),                                  //   input,    width = 1,                             i_pma_ctrl.data
		.i_pcie_pcs_rx_rst                           (i_pcie_pcs_rx_rst),                           //   input,    width = 1,                      i_pcie_pcs_rx_rst.data
		.i_pcie_pcs_tx_rst                           (i_pcie_pcs_tx_rst),                           //   input,    width = 1,                      i_pcie_pcs_tx_rst.data
		.i_rxeiosdetectstata                         (i_rxeiosdetectstata),                         //   input,    width = 1,                    i_rxeiosdetectstata.data
		.i_rxeq_precal_code_selnt                    (i_rxeq_precal_code_selnt),                    //   input,    width = 3,               i_rxeq_precal_code_selnt.data
		.i_rxeq_starta                               (i_rxeq_starta),                               //   input,    width = 1,                          i_rxeq_starta.data
		.i_rxeq_static_ena                           (i_rxeq_static_ena),                           //   input,    width = 1,                      i_rxeq_static_ena.data
		.i_rxmargin_direction_nt                     (i_rxmargin_direction_nt),                     //   input,    width = 1,                i_rxmargin_direction_nt.data
		.i_rxmargin_mode_nt                          (i_rxmargin_mode_nt),                          //   input,    width = 1,                     i_rxmargin_mode_nt.data
		.i_rxmargin_offset_change_a                  (i_rxmargin_offset_change_a),                  //   input,    width = 1,             i_rxmargin_offset_change_a.data
		.i_rxmargin_offset_nt                        (i_rxmargin_offset_nt),                        //   input,    width = 7,                   i_rxmargin_offset_nt.data
		.i_rxmargin_start_a                          (i_rxmargin_start_a),                          //   input,    width = 1,                     i_rxmargin_start_a.data
		.i_rxpstate                                  (i_rxpstate),                                  //   input,    width = 3,                             i_rxpstate.data
		.i_rxrate                                    (i_rxrate),                                    //   input,    width = 4,                               i_rxrate.data
		.i_rxterm_hiz_ena                            (i_rxterm_hiz_ena),                            //   input,    width = 1,                       i_rxterm_hiz_ena.data
		.i_rxwidth                                   (i_rxwidth),                                   //   input,    width = 3,                              i_rxwidth.data
		.i_tstbus_lane                               (i_tstbus_lane),                               //   input,    width = 1,                          i_tstbus_lane.data
		.i_txbeacona                                 (i_txbeacona),                                 //   input,    width = 1,                            i_txbeacona.data
		.i_txclkdivrate                              (i_txclkdivrate),                              //   input,    width = 3,                         i_txclkdivrate.data
		.i_txdetectrx_reqa                           (i_txdetectrx_reqa),                           //   input,    width = 1,                      i_txdetectrx_reqa.data
		.i_txdrv_levn                                (i_txdrv_levn),                                //   input,    width = 6,                           i_txdrv_levn.data
		.i_txdrv_levnm1                              (i_txdrv_levnm1),                              //   input,    width = 5,                         i_txdrv_levnm1.data
		.i_txdrv_levnm2                              (i_txdrv_levnm2),                              //   input,    width = 3,                         i_txdrv_levnm2.data
		.i_txdrv_levnp1                              (i_txdrv_levnp1),                              //   input,    width = 5,                         i_txdrv_levnp1.data
		.i_txdrv_slew                                (i_txdrv_slew),                                //   input,    width = 4,                           i_txdrv_slew.data
		.i_txelecidle                                (i_txelecidle),                                //   input,    width = 4,                           i_txelecidle.data
		.i_txpstate                                  (i_txpstate),                                  //   input,    width = 3,                             i_txpstate.data
		.i_txrate                                    (i_txrate),                                    //   input,    width = 4,                               i_txrate.data
		.i_txwidth                                   (i_txwidth),                                   //   input,    width = 3,                              i_txwidth.data
		.i_hio_pld_rx_clk_in_row_clk                 (i_hio_pld_rx_clk_in_row_clk),                 //   input,    width = 1,            i_hio_pld_rx_clk_in_row_clk.clk
		.i_hio_pld_tx_clk_in_row_clk                 (i_hio_pld_tx_clk_in_row_clk),                 //   input,    width = 1,            i_hio_pld_tx_clk_in_row_clk.clk
		.i_hio_det_lat_rx_dl_clk                     (i_hio_det_lat_rx_dl_clk),                     //   input,    width = 1,                i_hio_det_lat_rx_dl_clk.clk
		.i_hio_det_lat_rx_mux_select                 (i_hio_det_lat_rx_mux_select),                 //   input,    width = 1,            i_hio_det_lat_rx_mux_select.clk
		.i_hio_det_lat_rx_sclk_flop                  (i_hio_det_lat_rx_sclk_flop),                  //   input,    width = 1,             i_hio_det_lat_rx_sclk_flop.clk
		.i_hio_det_lat_rx_sclk_gen_clk               (i_hio_det_lat_rx_sclk_gen_clk),               //   input,    width = 1,          i_hio_det_lat_rx_sclk_gen_clk.clk
		.i_hio_det_lat_rx_trig_flop                  (i_hio_det_lat_rx_trig_flop),                  //   input,    width = 1,             i_hio_det_lat_rx_trig_flop.clk
		.i_hio_det_lat_sampling_clk                  (i_hio_det_lat_sampling_clk),                  //   input,    width = 1,             i_hio_det_lat_sampling_clk.clk
		.i_hio_det_lat_tx_dl_clk                     (i_hio_det_lat_tx_dl_clk),                     //   input,    width = 1,                i_hio_det_lat_tx_dl_clk.clk
		.i_hio_det_lat_tx_mux_select                 (i_hio_det_lat_tx_mux_select),                 //   input,    width = 1,            i_hio_det_lat_tx_mux_select.clk
		.i_hio_det_lat_tx_sclk_flop                  (i_hio_det_lat_tx_sclk_flop),                  //   input,    width = 1,             i_hio_det_lat_tx_sclk_flop.clk
		.i_hio_det_lat_tx_sclk_gen_clk               (i_hio_det_lat_tx_sclk_gen_clk),               //   input,    width = 1,          i_hio_det_lat_tx_sclk_gen_clk.clk
		.i_hio_det_lat_tx_trig_flop                  (i_hio_det_lat_tx_trig_flop),                  //   input,    width = 1,             i_hio_det_lat_tx_trig_flop.clk
		.rx_serial_n                                 (rx_serial_n),                                 //   input,    width = 1,                            rx_serial_n.data
		.rx_serial_p                                 (rx_serial_p),                                 //   input,    width = 1,                            rx_serial_p.data
		.o_hio_txdata_fifo_wr_empty                  (o_hio_txdata_fifo_wr_empty),                  //  output,    width = 1,             o_hio_txdata_fifo_wr_empty.data
		.o_hio_txdata_fifo_wr_pempty                 (o_hio_txdata_fifo_wr_pempty),                 //  output,    width = 1,            o_hio_txdata_fifo_wr_pempty.data
		.o_hio_txdata_fifo_wr_full                   (o_hio_txdata_fifo_wr_full),                   //  output,    width = 1,              o_hio_txdata_fifo_wr_full.data
		.o_hio_txdata_fifo_wr_pfull                  (o_hio_txdata_fifo_wr_pfull),                  //  output,    width = 1,             o_hio_txdata_fifo_wr_pfull.data
		.o_hio_rxdata                                (o_hio_rxdata),                                //  output,   width = 80,                           o_hio_rxdata.data
		.o_hio_rxdata_extra                          (o_hio_rxdata_extra),                          //  output,   width = 10,                     o_hio_rxdata_extra.data
		.o_hio_rxdata_fifo_rd_empty                  (o_hio_rxdata_fifo_rd_empty),                  //  output,    width = 1,             o_hio_rxdata_fifo_rd_empty.data
		.o_hio_rxdata_fifo_rd_pempty                 (o_hio_rxdata_fifo_rd_pempty),                 //  output,    width = 1,            o_hio_rxdata_fifo_rd_pempty.data
		.o_hio_rxdata_fifo_rd_full                   (o_hio_rxdata_fifo_rd_full),                   //  output,    width = 1,              o_hio_rxdata_fifo_rd_full.data
		.o_hio_rxdata_fifo_rd_pfull                  (o_hio_rxdata_fifo_rd_pfull),                  //  output,    width = 1,             o_hio_rxdata_fifo_rd_pfull.data
		.o_hio_rstepcs_rx_pcs_fully_aligned          (o_hio_rstepcs_rx_pcs_fully_aligned),          //  output,    width = 1,     o_hio_rstepcs_rx_pcs_fully_aligned.reset
		.o_hio_rstfec_fec_rx_rdy_n                   (o_hio_rstfec_fec_rx_rdy_n),                   //  output,    width = 1,              o_hio_rstfec_fec_rx_rdy_n.reset
		.o_hio_rst_flux0_cpi_cmn_busy                (o_hio_rst_flux0_cpi_cmn_busy),                //  output,    width = 1,           o_hio_rst_flux0_cpi_cmn_busy.reset
		.o_hio_rst_oflux_rx_srds_rdy                 (o_hio_rst_oflux_rx_srds_rdy),                 //  output,    width = 1,            o_hio_rst_oflux_rx_srds_rdy.reset
		.o_hio_rst_ux_all_synthlockstatus            (o_hio_rst_ux_all_synthlockstatus),            //  output,    width = 1,       o_hio_rst_ux_all_synthlockstatus.reset
		.o_hio_rst_ux_octl_pcs_rxstatus              (o_hio_rst_ux_octl_pcs_rxstatus),              //  output,    width = 1,         o_hio_rst_ux_octl_pcs_rxstatus.reset
		.o_hio_rst_ux_octl_pcs_txstatus              (o_hio_rst_ux_octl_pcs_txstatus),              //  output,    width = 1,         o_hio_rst_ux_octl_pcs_txstatus.reset
		.o_hio_rst_ux_rxcdrlock2data                 (o_hio_rst_ux_rxcdrlock2data),                 //  output,    width = 1,            o_hio_rst_ux_rxcdrlock2data.reset
		.o_hio_rst_ux_rxcdrlockstatus                (o_hio_rst_ux_rxcdrlockstatus),                //  output,    width = 1,           o_hio_rst_ux_rxcdrlockstatus.reset
		.o_hio_uxquad_async                          (o_hio_uxquad_async),                          //  output,   width = 50,                     o_hio_uxquad_async.data
		.o_hio_user_rx_clk1_clk                      (o_hio_user_rx_clk1_clk),                      //  output,    width = 1,                 o_hio_user_rx_clk1_clk.clk
		.o_hio_user_rx_clk2_clk                      (o_hio_user_rx_clk2_clk),                      //  output,    width = 1,                 o_hio_user_rx_clk2_clk.clk
		.o_hio_user_tx_clk1_clk                      (o_hio_user_tx_clk1_clk),                      //  output,    width = 1,                 o_hio_user_tx_clk1_clk.clk
		.o_hio_user_tx_clk2_clk                      (o_hio_user_tx_clk2_clk),                      //  output,    width = 1,                 o_hio_user_tx_clk2_clk.clk
		.o_hio_ux_chnl_refclk_mux                    (o_hio_ux_chnl_refclk_mux),                    //  output,    width = 1,               o_hio_ux_chnl_refclk_mux.clk
		.o_hio_det_lat_rx_async_dl_sync              (o_hio_det_lat_rx_async_dl_sync),              //  output,    width = 1,         o_hio_det_lat_rx_async_dl_sync.clk
		.o_hio_det_lat_rx_async_pulse                (o_hio_det_lat_rx_async_pulse),                //  output,    width = 1,           o_hio_det_lat_rx_async_pulse.clk
		.o_hio_det_lat_rx_async_sample_sync          (o_hio_det_lat_rx_async_sample_sync),          //  output,    width = 1,     o_hio_det_lat_rx_async_sample_sync.clk
		.o_hio_det_lat_rx_sclk_sample_sync           (o_hio_det_lat_rx_sclk_sample_sync),           //  output,    width = 1,      o_hio_det_lat_rx_sclk_sample_sync.clk
		.o_hio_det_lat_rx_trig_sample_sync           (o_hio_det_lat_rx_trig_sample_sync),           //  output,    width = 1,      o_hio_det_lat_rx_trig_sample_sync.clk
		.o_hio_det_lat_tx_async_dl_sync              (o_hio_det_lat_tx_async_dl_sync),              //  output,    width = 1,         o_hio_det_lat_tx_async_dl_sync.clk
		.o_hio_det_lat_tx_async_pulse                (o_hio_det_lat_tx_async_pulse),                //  output,    width = 1,           o_hio_det_lat_tx_async_pulse.clk
		.o_hio_det_lat_tx_async_sample_sync          (o_hio_det_lat_tx_async_sample_sync),          //  output,    width = 1,     o_hio_det_lat_tx_async_sample_sync.clk
		.o_hio_det_lat_tx_sclk_sample_sync           (o_hio_det_lat_tx_sclk_sample_sync),           //  output,    width = 1,      o_hio_det_lat_tx_sclk_sample_sync.clk
		.o_hio_det_lat_tx_trig_sample_sync           (o_hio_det_lat_tx_trig_sample_sync),           //  output,    width = 1,      o_hio_det_lat_tx_trig_sample_sync.clk
		.o_hio_xcvrif_rx_latency_pulse               (o_hio_xcvrif_rx_latency_pulse),               //  output,    width = 1,          o_hio_xcvrif_rx_latency_pulse.clk
		.o_hio_xcvrif_tx_latency_pulse               (o_hio_xcvrif_tx_latency_pulse),               //  output,    width = 1,          o_hio_xcvrif_tx_latency_pulse.clk
		.tx_serial_p                                 (tx_serial_p),                                 //  output,    width = 1,                            tx_serial_p.data
		.tx_serial_n                                 (tx_serial_n),                                 //  output,    width = 1,                            tx_serial_n.data
		.i_hio_txdata_async                          (i_hio_txdata_async),                          //   input,  width = 100,                     i_hio_txdata_async.data
		.i_hio_txdata_direct                         (i_hio_txdata_direct),                         //   input,   width = 10,                    i_hio_txdata_direct.data
		.o_hio_rxdata_async                          (o_hio_rxdata_async),                          //  output,  width = 100,                     o_hio_rxdata_async.data
		.o_hio_rxdata_direct                         (o_hio_rxdata_direct),                         //  output,   width = 10,                    o_hio_rxdata_direct.data
		.i_uxwrap_bus_in_phy_shared                  (i_uxwrap_bus_in_phy_shared),                  //   input,  width = 768,                          uxwrap_bus_in.data
		.o_uxwrap_bus_out_phy_shared                 (o_uxwrap_bus_out_phy_shared),                 //  output,  width = 704,                         uxwrap_bus_out.data
		.o_lavmm_addr_phy_shared                     (o_lavmm_addr_phy_shared),                     //  output,   width = 20,                    reconfig_phy_shared.address
		.o_lavmm_be_phy_shared                       (o_lavmm_be_phy_shared),                       //  output,    width = 4,                                       .byteenable
		.o_lavmm_read_phy_shared                     (o_lavmm_read_phy_shared),                     //  output,    width = 1,                                       .read
		.o_lavmm_wdata_phy_shared                    (o_lavmm_wdata_phy_shared),                    //  output,   width = 32,                                       .writedata
		.o_lavmm_write_phy_shared                    (o_lavmm_write_phy_shared),                    //  output,    width = 1,                                       .write
		.i_lavmm_rdata_phy_shared                    (i_lavmm_rdata_phy_shared),                    //   input,   width = 32,                                       .readdata
		.i_lavmm_rdata_valid_phy_shared              (i_lavmm_rdata_valid_phy_shared),              //   input,    width = 1,                                       .readdatavalid
		.i_lavmm_waitreq_phy_shared                  (i_lavmm_waitreq_phy_shared),                  //   input,    width = 1,                                       .waitrequest
		.o_lavmm_clk_phy_shared                      (o_lavmm_clk_phy_shared),                      //  output,    width = 1,                reconfig_clk_phy_shared.clk
		.o_lavmm_rstn_phy_shared                     (o_lavmm_rstn_phy_shared),                     //  output,    width = 1,                reconfig_rst_phy_shared.reset
		.o_sclk_return_sel_rx_phy_shared             (o_sclk_return_sel_rx_phy_shared),             //  output,    width = 1,                   o_sclk_return_sel_rx.data
		.o_sclk_return_sel_tx_phy_shared             (o_sclk_return_sel_tx_phy_shared),             //  output,    width = 1,                   o_sclk_return_sel_tx.data
		.o_ick_sclk_rx_phy_shared                    (o_ick_sclk_rx_phy_shared),                    //  output,    width = 1,                          o_ick_sclk_rx.clk
		.i_sync_common_control_phy_shared            (i_sync_common_control_phy_shared),            //   input,    width = 5,                  i_sync_common_control.data
		.o_ft_rx_sclk_sync_ch_phy_shared             (o_ft_rx_sclk_sync_ch_phy_shared),             //  output,    width = 1,                   o_ft_rx_sclk_sync_ch.data
		.o_ft_tx_sclk_sync_ch_phy_shared             (o_ft_tx_sclk_sync_ch_phy_shared),             //  output,    width = 1,                   o_ft_tx_sclk_sync_ch.data
		.o_rst_ux_rx_pma_rst_n_phy_shared            (o_rst_ux_rx_pma_rst_n_phy_shared),            //  output,    width = 1,                  o_rst_ux_rx_pma_rst_n.reset
		.o_rst_ux_tx_pma_rst_n_phy_shared            (o_rst_ux_tx_pma_rst_n_phy_shared),            //  output,    width = 1,                  o_rst_ux_tx_pma_rst_n.reset
		.o_ick_pcs_txword_phy_shared                 (o_ick_pcs_txword_phy_shared),                 //  output,    width = 1,                       o_ick_pcs_txword.data
		.o_tx_dl_ch_bit_phy_shared                   (o_tx_dl_ch_bit_phy_shared),                   //  output,    width = 1,                         o_tx_dl_ch_bit.data
		.i_dat_pcs_measlatbit_phy_shared             (i_dat_pcs_measlatbit_phy_shared),             //   input,    width = 1,                   i_dat_pcs_measlatbit.data
		.i_ft_rx_async_pulse_ch_phy_shared           (i_ft_rx_async_pulse_ch_phy_shared),           //   input,    width = 1,                 i_ft_rx_async_pulse_ch.data
		.i_ft_tx_async_pulse_ch_phy_shared           (i_ft_tx_async_pulse_ch_phy_shared),           //   input,    width = 1,                 i_ft_tx_async_pulse_ch.data
		.i_rx_dl_ch_bit_phy_shared                   (i_rx_dl_ch_bit_phy_shared),                   //   input,    width = 1,                         i_rx_dl_ch_bit.data
		.i_ux_rxuser1_sel_phy_shared                 (i_ux_rxuser1_sel_phy_shared),                 //   input,    width = 2,                       i_ux_rxuser1_sel.data
		.i_ux_rxuser2_sel_phy_shared                 (i_ux_rxuser2_sel_phy_shared),                 //   input,    width = 2,                       i_ux_rxuser2_sel.data
		.i_ux_txuser1_sel_phy_shared                 (i_ux_txuser1_sel_phy_shared),                 //   input,    width = 2,                       i_ux_txuser1_sel.data
		.i_ux_txuser2_sel_phy_shared                 (i_ux_txuser2_sel_phy_shared),                 //   input,    width = 2,                       i_ux_txuser2_sel.data
		.o_octl_pcs_txstatus_a_phy_shared            (o_octl_pcs_txstatus_a_phy_shared),            //  output,    width = 1,                  o_octl_pcs_txstatus_a.data
		.i_ictl_pcs_txenable_a_phy_shared            (i_ictl_pcs_txenable_a_phy_shared),            //   input,    width = 1,                  i_ictl_pcs_txenable_a.data
		.i_sync_cfg_data_phy_shared                  (i_sync_cfg_data_phy_shared),                  //   input,  width = 125,                        i_sync_cfg_data.data
		.i_sync_interface_control_phy_shared         (i_sync_interface_control_phy_shared),         //   input,  width = 250,               i_sync_interface_control.data
		.o_tx_data_phy_shared                        (o_tx_data_phy_shared),                        //  output,   width = 80,                              o_tx_data.data
		.i_rx_data_phy_shared                        (i_rx_data_phy_shared),                        //   input,   width = 80,                              i_rx_data.data
		.o_sm_flux_ingress_phy_shared                (o_sm_flux_ingress_phy_shared),                //  output,  width = 320,                      o_sm_flux_ingress.data
		.i_sm_flux_egress_phy_shared                 (i_sm_flux_egress_phy_shared),                 //   input,  width = 257,                       i_sm_flux_egress.data
		.i_flux_cpi_int_phy_shared                   (i_flux_cpi_int_phy_shared),                   //   input,    width = 1,                         i_flux_cpi_int.data
		.i_flux_int_phy_shared                       (i_flux_int_phy_shared),                       //   input,    width = 1,                             i_flux_int.data
		.i_oflux_octl_pcs_txptr_smpl_lane_phy_shared (i_oflux_octl_pcs_txptr_smpl_lane_phy_shared), //   input,    width = 1,       i_oflux_octl_pcs_txptr_smpl_lane.data
		.o_ick_sclk_tx_phy_shared                    (o_ick_sclk_tx_phy_shared),                    //  output,    width = 1,                          o_ick_sclk_tx.clk
		.i_flux_srds_rdy_phy_shared                  (i_flux_srds_rdy_phy_shared),                  //   input,    width = 1,                        i_flux_srds_rdy.data
		.i_pcs_rxword_phy_shared                     (i_pcs_rxword_phy_shared),                     //   input,    width = 1,                           i_pcs_rxword.data
		.i_pcs_rxpostdiv_phy_shared                  (i_pcs_rxpostdiv_phy_shared),                  //   input,    width = 1,                        i_pcs_rxpostdiv.data
		.i_ock_pcs_txword_phy_shared                 (i_ock_pcs_txword_phy_shared),                 //   input,    width = 1,                       i_ock_pcs_txword.data
		.o_dat_pcs_measlatrndtripbit_phy_shared      (o_dat_pcs_measlatrndtripbit_phy_shared),      //  output,    width = 1, o_dat_pcs_measlatrndtripbit_phy_shared.data
		.i_ch_eth_fec_rx_async_fec_wrap              (i_ch_eth_fec_rx_async_fec_wrap),              //   input,   width = 12,                            asyncdata_4.data
		.i_ch_eth_fec_rx_direct_fec_wrap             (i_ch_eth_fec_rx_direct_fec_wrap),             //   input,    width = 1,                            asyncdata_5.data
		.i_fec_rx_rdy_n_fec_wrap                     (i_fec_rx_rdy_n_fec_wrap),                     //   input,    width = 1,                i_fec_rx_rdy_n_fec_wrap.data
		.i_fec_tx_data_mux_sel_fec_wrap              (i_fec_tx_data_mux_sel_fec_wrap),              //   input,    width = 1,         i_fec_tx_data_mux_sel_fec_wrap.muxsel
		.i_fec_rx_data_fec_wrap                      (i_fec_rx_data_fec_wrap),                      //   input,   width = 43,                 i_fec_rx_data_fec_wrap.data
		.i_xcvr_tx_data                              (i_xcvr_tx_data),                              //   input,   width = 43,                         i_xcvr_tx_data.data
		.ss_rst_flux0_cpi_cmn_busy                   (ss_rst_flux0_cpi_cmn_busy),                   //  output,    width = 1,              ss_rst_flux0_cpi_cmn_busy.data
		.o_pma_rx_sf                                 (o_pma_rx_sf),                                 //  output,    width = 1,                            o_pma_rx_sf.data
		.i_refclk_tx_p                               (i_refclk_tx_p),                               //   input,    width = 1,                          i_refclk_tx_p.clk
		.i_syspll_c0_clk                             (i_syspll_c0_clk),                             //   input,    width = 1,                        i_syspll_c0_clk.clk
		.i_syspll_c1_clk                             (i_syspll_c1_clk),                             //   input,    width = 1,                        i_syspll_c1_clk.clk
		.i_syspll_c2_clk                             (i_syspll_c2_clk),                             //   input,    width = 1,                        i_syspll_c2_clk.clk
		.i_flux_clk                                  (i_flux_clk),                                  //   input,    width = 1,                             i_flux_clk.clk
		.i_refclk_rx_p                               (i_refclk_rx_p),                               //   input,    width = 1,                          i_refclk_rx_p.clk
		.i_ux_chnl_refclk_mux_phy_shared             (i_ux_chnl_refclk_mux_phy_shared),             //   input,    width = 1,        i_ux_chnl_refclk_mux_phy_shared.clk
		.o_xcvrif_tx_fifo_rd_en_mux_x1               (o_xcvrif_tx_fifo_rd_en_mux_x1),               //  output,    width = 1,          o_xcvrif_tx_fifo_rd_en_mux_x1.clk
		.i_xcvrif_tx_fifo_rd_en_mux_x2               (i_xcvrif_tx_fifo_rd_en_mux_x2),               //   input,    width = 1,          i_xcvrif_tx_fifo_rd_en_mux_x2.clk
		.i_xcvrif_tx_fifo_rd_en_mux_x4               (i_xcvrif_tx_fifo_rd_en_mux_x4),               //   input,    width = 1,          i_xcvrif_tx_fifo_rd_en_mux_x4.clk
		.i_xcvrif_tx_fifo_rd_en_mux_x6_bot           (i_xcvrif_tx_fifo_rd_en_mux_x6_bot),           //   input,    width = 1,      i_xcvrif_tx_fifo_rd_en_mux_x6_bot.clk
		.i_xcvrif_tx_fifo_rd_en_mux_x6_top           (i_xcvrif_tx_fifo_rd_en_mux_x6_top),           //   input,    width = 1,      i_xcvrif_tx_fifo_rd_en_mux_x6_top.clk
		.i_xcvrif_tx_fifo_rd_en_mux_x8_bot           (i_xcvrif_tx_fifo_rd_en_mux_x8_bot),           //   input,    width = 1,      i_xcvrif_tx_fifo_rd_en_mux_x8_bot.clk
		.i_xcvrif_tx_fifo_rd_en_mux_x8_top           (i_xcvrif_tx_fifo_rd_en_mux_x8_top),           //   input,    width = 1,      i_xcvrif_tx_fifo_rd_en_mux_x8_top.clk
		.o_xcvrif_tx_rst_mux_x1                      (o_xcvrif_tx_rst_mux_x1),                      //  output,    width = 1,                 o_xcvrif_tx_rst_mux_x1.clk
		.i_xcvrif_tx_rst_mux_x2                      (i_xcvrif_tx_rst_mux_x2),                      //   input,    width = 1,                 i_xcvrif_tx_rst_mux_x2.clk
		.i_xcvrif_tx_rst_mux_x4                      (i_xcvrif_tx_rst_mux_x4),                      //   input,    width = 1,                 i_xcvrif_tx_rst_mux_x4.clk
		.i_xcvrif_tx_rst_mux_x6_bot                  (i_xcvrif_tx_rst_mux_x6_bot),                  //   input,    width = 1,             i_xcvrif_tx_rst_mux_x6_bot.clk
		.i_xcvrif_tx_rst_mux_x6_top                  (i_xcvrif_tx_rst_mux_x6_top),                  //   input,    width = 1,             i_xcvrif_tx_rst_mux_x6_top.clk
		.i_xcvrif_tx_rst_mux_x8_bot                  (i_xcvrif_tx_rst_mux_x8_bot),                  //   input,    width = 1,             i_xcvrif_tx_rst_mux_x8_bot.clk
		.i_xcvrif_tx_rst_mux_x8_top                  (i_xcvrif_tx_rst_mux_x8_top),                  //   input,    width = 1,             i_xcvrif_tx_rst_mux_x8_top.clk
		.o_xcvrif_tx_word_clk_mux_x1                 (o_xcvrif_tx_word_clk_mux_x1),                 //  output,    width = 1,            o_xcvrif_tx_word_clk_mux_x1.clk
		.i_xcvrif_tx_word_clk_mux_x2                 (i_xcvrif_tx_word_clk_mux_x2),                 //   input,    width = 1,            i_xcvrif_tx_word_clk_mux_x2.clk
		.i_xcvrif_tx_word_clk_mux_x4                 (i_xcvrif_tx_word_clk_mux_x4),                 //   input,    width = 1,            i_xcvrif_tx_word_clk_mux_x4.clk
		.i_xcvrif_tx_word_clk_mux_x6_bot             (i_xcvrif_tx_word_clk_mux_x6_bot),             //   input,    width = 1,        i_xcvrif_tx_word_clk_mux_x6_bot.clk
		.i_xcvrif_tx_word_clk_mux_x6_top             (i_xcvrif_tx_word_clk_mux_x6_top),             //   input,    width = 1,        i_xcvrif_tx_word_clk_mux_x6_top.clk
		.i_xcvrif_tx_word_clk_mux_x8_bot             (i_xcvrif_tx_word_clk_mux_x8_bot),             //   input,    width = 1,        i_xcvrif_tx_word_clk_mux_x8_bot.clk
		.i_xcvrif_tx_word_clk_mux_x8_top             (i_xcvrif_tx_word_clk_mux_x8_top),             //   input,    width = 1,        i_xcvrif_tx_word_clk_mux_x8_top.clk
		.ioack_cdrdiv_left_ux_bidir_in               (ioack_cdrdiv_left_ux_bidir_in),               //   input,    width = 1,          ioack_cdrdiv_left_ux_bidir_in.clk
		.ioack_synthdiv1_left_ux_bidir_in            (ioack_synthdiv1_left_ux_bidir_in),            //   input,    width = 1,       ioack_synthdiv1_left_ux_bidir_in.clk
		.ioack_synthdiv2_left_ux_bidir_in            (ioack_synthdiv2_left_ux_bidir_in),            //   input,    width = 1,       ioack_synthdiv2_left_ux_bidir_in.clk
		.ioack_cdrdiv_left_ux_bidir_out              (ioack_cdrdiv_left_ux_bidir_out),              //  output,    width = 1,         ioack_cdrdiv_left_ux_bidir_out.clk
		.ioack_synthdiv1_left_ux_bidir_out           (ioack_synthdiv1_left_ux_bidir_out),           //  output,    width = 1,      ioack_synthdiv1_left_ux_bidir_out.clk
		.ioack_synthdiv2_left_ux_bidir_out           (ioack_synthdiv2_left_ux_bidir_out),           //  output,    width = 1,      ioack_synthdiv2_left_ux_bidir_out.clk
		.o_xcvrif_tx_rst_wr_sync_mux_x1              (o_xcvrif_tx_rst_wr_sync_mux_x1),              //  output,    width = 1,         o_xcvrif_tx_rst_wr_sync_mux_x1.clk
		.i_xcvrif_tx_rst_wr_sync_mux_x2              (i_xcvrif_tx_rst_wr_sync_mux_x2),              //   input,    width = 1,         i_xcvrif_tx_rst_wr_sync_mux_x2.clk
		.i_xcvrif_tx_rst_wr_sync_mux_x4              (i_xcvrif_tx_rst_wr_sync_mux_x4),              //   input,    width = 1,         i_xcvrif_tx_rst_wr_sync_mux_x4.clk
		.i_xcvrif_tx_rst_wr_sync_mux_x6_bot          (i_xcvrif_tx_rst_wr_sync_mux_x6_bot),          //   input,    width = 1,     i_xcvrif_tx_rst_wr_sync_mux_x6_bot.clk
		.i_xcvrif_tx_rst_wr_sync_mux_x6_top          (i_xcvrif_tx_rst_wr_sync_mux_x6_top),          //   input,    width = 1,     i_xcvrif_tx_rst_wr_sync_mux_x6_top.clk
		.i_xcvrif_tx_rst_wr_sync_mux_x8_bot          (i_xcvrif_tx_rst_wr_sync_mux_x8_bot),          //   input,    width = 1,     i_xcvrif_tx_rst_wr_sync_mux_x8_bot.clk
		.i_xcvrif_tx_rst_wr_sync_mux_x8_top          (i_xcvrif_tx_rst_wr_sync_mux_x8_top),          //   input,    width = 1,     i_xcvrif_tx_rst_wr_sync_mux_x8_top.clk
		.ss_user_rx_clk1_clk                         (ss_user_rx_clk1_clk),                         //  output,    width = 1,                    ss_user_rx_clk1_clk.clk
		.ss_user_rx_clk2_clk                         (ss_user_rx_clk2_clk),                         //  output,    width = 1,                    ss_user_rx_clk2_clk.clk
		.ss_user_tx_clk1_clk                         (ss_user_tx_clk1_clk),                         //  output,    width = 1,                    ss_user_tx_clk1_clk.clk
		.ss_user_tx_clk2_clk                         (ss_user_tx_clk2_clk),                         //  output,    width = 1,                    ss_user_tx_clk2_clk.clk
		.ss_user_rx_clk1_clk_w                       (ss_user_rx_clk1_clk_w),                       //  output,    width = 1,                  ss_user_rx_clk1_clk_w.clk
		.ss_user_rx_clk2_clk_w                       (ss_user_rx_clk2_clk_w),                       //  output,    width = 1,                  ss_user_rx_clk2_clk_w.clk
		.ss_user_tx_clk1_clk_w                       (ss_user_tx_clk1_clk_w),                       //  output,    width = 1,                  ss_user_tx_clk1_clk_w.clk
		.ss_user_tx_clk2_clk_w                       (ss_user_tx_clk2_clk_w),                       //  output,    width = 1,                  ss_user_tx_clk2_clk_w.clk
		.o_hio_ux_tx_ch_ptr_smpl                     (o_hio_ux_tx_ch_ptr_smpl)                      //  output,    width = 1,                o_hio_ux_tx_ch_ptr_smpl.data
	);

endmodule
