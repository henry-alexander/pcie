//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pspY1WcG/b5Bwv7r7UUGPRQ4yBHRQ9WHaYIXYYJwuXcqE1G46HMlgnzhMAXW
NgRLxpOONlZC87U/Y3qBzkF2udXFprUyWG4yoYitCEvPFyJ+DpgqzJueAI+a
xTUU78O2iebl5WDulrVXNGl6TssrmrijD76ZLd7gs9PKnPO5BTqFsmqSJGlJ
GdJ+RhCKZOTTTe8cftfIBCshgFOeR2rlOYxQIkySZexyZqjC6nri3yWs/LLj
G1lpUSvoVKx2cHmLcPYZklYsc8KM6EcuQjw/0KVEXxwdrYpvMWxeTXzojwye
ol0uURgnt89J8Yx4exsA8hbEvfz4MOsOl5fnV0pj6Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
DpDilrVWZZeVzGtUXYvzP+BiVerHaWoxCUGf0uWuJ3PkQhdK2zXtXAVlpGXD
HnfpCL/6SPfYDaBsYNvgFg6e3GiXseD8h80QKKFvpr41fDz6zzps0p7f7kFN
KAe64fsrWLZHm5/FkRjjNp3dgW0DN3eYSWbNvpn1lAa0oaMBjEmsqPMru/vx
/4gRevn14KPTJHeS33wi5AGKDVp9jD32x1mKy1hHjCXiwqc7dbPFUNWzlU3v
A3InQAmG4esnWwBBzCht+KjzSkkHpiU4hPIyX0Qmr1fgnWIcSRRFS6961h7W
FZ6TLY+8DZtq1yfJpIPtxQxFeg0uukS31lDipqdm1Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
kGrPV4QkAcPJfjPE9xU3t7xTUmLsFsCZXj9UVv3NdJr0I2pdJ9XzMxA7IUhf
kUJUuaOy+ZAAHJaV1nEqM7F70/hqiybpqWHGdFKMk2mYaUDcj8/SvAkB4Fjx
tQJFq8LwBeJlmA+oxVYzGlKRW7nlmVDvy5KxJLmutI/hGCI96FI9IgsS7ly2
l+EGpn7eRkmAgODbqVg04AVCQxwz+32+m3Q5ebNsyrrv2yUWg+znbXWlf5Oi
ssgqbQJBlK/LATT1Y/bsXGOmM3bfK5R+BLO0wFifHlkGoVp24/ZuyIWebWON
Wt0uNEAJ7gaUoaMBCJekCxVXMB1zc9D3b+jOsEH+ZA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FwcLZc0rlimofXXTW9qO91/+9dLojKjaKGhh0Vl03+311L1Lp0f/TnJoHt0E
zg1WYOaxA0DiMtLr9hHFvHJFJ7IVN1DFQc286WHZfy+Ej6rSfe/40Kka2v2u
BE/Aq/0DnLVWMCaYYuEmHkw1mYsZXujZTTT6m03yUUYFMc2LK0c=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
GIoFpypjC8jY4Bmka2s3BQ2wThW/4W4UggR9VWkKcWzE+kKxB/Vh+nLu8Dd2
FwNfyOpU+CJk95PJcGn/TBUobtBMzFqFpCbSAzh8UjYMCXJS4fP6RMFquXVj
NZ2/6fKD3Cv51c4q/w4KaQgDjrYSlAFe4HDj0BJKApFHEwcNLs9gQUL1uz3C
yBSBBBy/2q548fWxeb9Ibp0JNTSmgx2FB1eCT44dNJjGMTjgBJhByaHQUn74
nrSPK9wkEqVV2Q60Dy6h+ZdVLu2xIuwkMd6LlLZJL9KLvndiqRr413aCKS4a
/s1sG/yBitz06Xhrr8Z4OXgVFd0RekwUpUNZrudmjuVnl8CIaUWvssTm79EZ
HdcMAnx4ucomzWg2JKsa42LjphruXMxDWN4vacYuNBD32WbO0Iav83bm/45J
5CJh66FruTNACbV1lPkgGrC3mzw42NqTGQv9Du2Okec3x2ZoT3YhJ70+5/Q4
o7vttvRFI/WG2A6d+wLrNMFhqqGxgre7


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
foNthM1opp6ZBhubltimT/lhlhLKEG0z4F40gmn3bE3+gKS6Ywuwtc1b6DCT
6rXKGdWoYegTQ7yaEpT/7tNcYgKi52UZckuyF7DqmgfRCRhhw9unfgTmZD/N
kzTNAcOhAS0UVXcVdVOD5+TZNnwwlddoNpAvfRuDcuqzmDPWwZI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
fuPxPx2Blm0qC7edlmm2w4ROhxR/2po+6ZFbksLowoCsjhmYiRb2q93xRpad
DYCTxCjC9c/KIKL1i+D09eF90/j9sFUP8CfzR3UndfYVV9d+WKx6TzEoeLf5
HaO8+AzZzIOu4zttyxzP9kkx3RoeoG1amQdm3b537iBW7OWW9L8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 43072)
`pragma protect data_block
YKEwsSVpqohs7YnkQBkzPoD3drZhoEO0fJipq24W5CchkdPHJs4/EJvorjfr
pcUZsORhyB5Vd1MBP9EbSU+pOQNTrUiaVI2eU72ul5oW8vop4Wba9wUjt2W7
/2QnpWpcwt34PsfAQ0QdBYCuzL8b++T4lv3I8hUFZD8J+kRWd4RTgAtD6qjH
K9u1fZ4LTy6DpKP7+8hLE60ietedX6M6oarrfn2Jf+Hh7MBK+hq20m0zUx5V
WBrfMux9Tydc5A9iRNYMQfn9YrNB3NS7VEAYX0CH3ovuBWyRd+zCBEN5s7sD
QJ304IwlRQhmrLvAtFT/E58YZNPtaz7OV2oYbVZ6jGCRpHsiMd/LB5DwJUsd
vdHq0xmcd4o48DCnAB+4LFjjFs/giK63KHPwoTLiF609T6X0KTr8rtf/5Ge9
Egqo1bIpqRz/D1wTSV42i9ZlC22TxTiqiQretG6FaGuL2zx4mIgyIVNPjm+G
+j6NdE/yJCrqeKO4MLqxZhR9BnFA5g1RoQwaafN2qiRe/gBB3a/V4hMpPU+A
mOu3S2NlNLQ4eJLkBBpNQ7VxC3XX7kjWAapW2K0q/asFjwKYB0gsGKd005Mb
NHb2IDxZzdZkptlVZXvhosLUhmYsPPByI0bjKqdCqC3mM2iuuAW8nt3c7voI
jr6K13tj5CqdDYUgCJtfrSlt5SpNvMiZ4PjwZ3EaZi9k4QmWGzQ6YtbFnRRV
ipb7pMVzZTKspThSCD2laC/oUw8n5S6I7n+1e4Wpi5M7R3phMGPe6zYnYFc0
lfNb0hTbPOoFeEnUy8pxUCY4LO4OyjrfEuA5UgrHKIvx2/X6KwK2aPxL0kYO
EjXE5xo/G7D8NaanEv5SGV3Nxd1TfaCWDWGIpo0Zbsmiu5qwCZANCq5ng1BM
xHyenE75Ujo+TUxyGnPIzf9aQTjlRnoQYQE8zIZgvUmxbMdKVXCdA5vcQBGB
ZeffMZ6EEMYzhWFNR5EGW/VBkTqywFAEdWNcgvpB9BWJcslucfmM7WSHZtEX
3+O1yXBaFNtK378C6umLHc2Z0IiWa7vZKE2KRDK1s8QBPeJ4n5DXUY0xXQ7T
6c26MY1OZgDXR81Tmg7oz1Exz+VYaINVi/Cty404nxhorEwYytgCB4cNAhJC
EEkUcwG2Kdkah7V66vBVH8oiwrnJ03MDck+uIngF7Mr6Qu4uIO6pn/Y1/PW0
oqVcGM85DRJCofAnu5hG8Cy9VjYxU+2ZL0BeuSRBQzANKhb6nOPKO4T1ZYj8
+dkk/2mlz+5rKARtmihG+DFnB1uFYnkcEuQm4oMKzJbkAVoGg7jBF4Vj+LKw
eE4Uq/SDhwUk2eafI3PfGqMg11f6tH1s5WPSMYGdoBm3WlrK0+FWUa0b9xLk
Mo78D1i0d2EXzLwHIg4lw2v8QWSuj+i7K4zvPWqdwFvm9Erg0Hzw7N6UEvkB
TRbMesoZuSdvRXgb1lpxb2hRvm9n1+WwojZ491eoWj9fnTVeGKkJ4dvnTvl4
4EXHBP39rcrjpUzxZfim1iAHWc85hr+WmZ0lPJKNelQjzovcEQpG5C/1zYef
Nk1XVgr4qlWyhq7kWxZV5nS5xdiPuDnHy7KGauqaVHUxMZMMmlABJB3Ronx4
XFoI2/kn10GjXbAP0PGzSD+KkmTzgiqRvtWU8wj9u25Nmk5pgcao6Rejf5tL
dP2ONcK5Xv9PF8aGoMh0+ZmdOH66GlNHBVnkJPRTG4F9WCHqLRwnAPBL35AW
Xzk3C5IwyAHkTynIvGVHbfmeLozGQynOmKzCtXn2N5s2EXDUWA8BzEJ72INl
LOujd3e/MHrxHkkzwSwdUCbVyfCCkNEYU8kEQRSF9bnl6qpMntyXae3fYVe5
PHbDRHXB9+sehmn0xnigkJ+qOIRdXSA2Ubk6/x5I7JCni8IYP9ETPJzSCzmI
l2gNWc3cevdU/aBo/9PbS3pNPUAcYwV7GDLvf88+Z+9L+yjYEaiJTqkgEcLT
ToYJADy52pY7Ut+N4rVmBLDShn7YsekLO9wMDS78f9iJZeUBlN5aI0RTguOw
XqKY79PQe3ebm2kWoZ5XjjiVChC55Ra/xTfA9kb0GFfSUQNtWRudfv1lPSaO
sYVfaygrIW1v2hbFH9DZecAPOnRvILAyU+0AHYU9V7zJNWc4on0fIlwxtHb8
0k/PR3RYQE3Q5PJuxyqoPl5J8jk7U4WHmpJlWt75UA77Kc35Y/5TBp1oucQ/
5mr4gIWRm4IEaf2jUDWSP2RZEDqcOo7tuKHpHEaC24zNtupwBvUPRgbe8pDy
AXUtF26tOgFy3TVGlZe8eVdX8l1KryHrUjEOtxmlfmzegeEzeoD62/YLNbMW
Yu3swGCJMmd+F6ACPXBaVHX87HGNyhT+lIXJSqErDKqANdVkhtPnGAdBqBVW
45dn5QgZ5jslrv3PBGYCufFrtz9uDKPeoQKzSGUt5paiUXeMEK3dKnaz1OQe
T7wK8yIsBt23PY9obO32QZSWhQE2WC4JBFaOT6Dkd95SwtTNWvKje8qlZs5B
MFnTjko6J6G/sKJPJ2OQpXNDRrZBn5C5lbqSAWjSzW682MXoSxrui9UOyqpz
gb6pa7gA03Gkf2h/H66xMLRUxAcaqsNKAOI742U0yQOhNdkZg4lBV/2fWAzs
BaQgxhOaNnhPV5E7ivNWcXgJuvzIHi7/Gc694urwTQzvyKGzIXZuDafgAuuz
xjhF44HaaHqG0gkAPQRf0DhgApZgZXezohJwzAUp7h5f0CWTHCYehnTt2PDd
VgQSC4m8dbCYV7C5YIlHWE51DktT3OgsBxRD2mpZDJatngalZb1ODVi2TPNR
+ivJU1Gpaa8spBeQYYbcF1PFpcMPteZhggcpKzJyZrrAd9QeiBlM2rYVdbFw
zGAOHNDASeef7vLhHMGciBlkQN3u6mP4KuEVIYrR1aTLeztLqJA5QvJ+qzBz
NEXBzzOdsANQ75yGfFOSe8/1b76EiBzvExBXceUsCQrM7kRSP/6iEt7vGITk
mc9/tM8kmqRL5FPlvhYIo/ATQObrpTmKRYmt9FUQ8auIj8M3r8r0ndZqMpnk
wODDraD104+LUqadGAlOlfOjhrjaR4uzrs0l4XoDTBqLr8TGnvD5bqBvInsK
YN/A/ZitKm0CkrwaerUBf6yc1TPGdj6wokr20HMgoLosaUtnag2utyy8WZ1V
6c+/Pf9Ibw6QCV526FFIYKIk6oDbgvmK1GJVmtnxWhUhad/AoFsBFTpc73X5
rFm61BHbVI/iZggRHONHoP2SWgLbULqyhmvQwAQQ7/QohUTtrIJ1Qwn+1/MO
XK6c5sn4NtQBYjE8eZ0MlFP7PZgztMvLDWSj9VT1EjJr4z+AcxJEZzs7gHHR
9n2gY55+ZtpYI08HcRjbZ7wXC8rerB0qnFX5xnYhkhT/xZQlN3toUqbCZPC5
v/MmIWDCq647oJ0kgxfxCV3Q9vKXJLwwqgJmaDkaEA2907RR5w6KSBA0P624
9p/YAqkr+2EsxjhO+XN56xOB7ydB90CrEZr30j6JP7uVl03KwcZ68QQANfJY
Gn8BDbWCxTj9KJIhqjjk3wEqhk9TPcY77WLVdyuWtdwx++QKgGWtp5RB4Pz1
7rGhSjDf2Gl8pWZj/RI7jRHdDcqfGhf9T3RKW5eHz8vRhQbquUt6Yv7KAn81
P9pBVrfTRLKvqqCtreIXwwQSxPE8jJW0O2J8BJSSvFQNA/TO672zwphhCSIy
W0eF/kc6MmzIoxztVv0oZ4xmOlXvjRaEX8AUr23AxlW44rhMrXmT/UAfq54O
52w3iVWISreJXB7XIp1BPQ1sGSZ2CV6yC9TxY8N6597nNSpnIgTYTd9m3eRp
PmXz1T/XlrRUCtfc4p8Pb5jsHOhtXzC8KSvF4jqMJjSc7GHprtAmY1svHte8
yumtKAJx4r9K/0IXebavhdHhKGpTDGTO9kdbSLcFl3kDQp0fp0MjrWMpZHjc
XGF3LpK/xjjM76a/JX3WK9tuTmmS8lS7lpvGEJPkfSIGs33zFgh7hIwePNxs
5mTWCNQ/8o2B4bd0v2HkTYjn2Sz0126YT7fPH/8+wpe3hp3M1NFSncVed8hj
3yYMYq79WYYPq7G5I7mHfn73OhZ/3iYApphZjZHKinWw2Swwbou1wjP6Cki5
p19wADAc27UdMRBVMtMs/N5kI1OubXjqzsOZSger7M2Cn4bxbxOvbTNswJj7
wpY90zPs69qsqg9yws6jFPJ+4xUTki6+yHD036NA+oE8svxpeuqn4Ykgq1RZ
QEzQAm0KllqtH1JglaKeQ7H/IqZ6+n2LfVJugEASby26YgRiGDdNlLHLN3Ev
P9W+9fkg48Rg+VfNX384js4oV1/1XYl88dnJbRTVwC3/rGOeotjLKajcIdkZ
xErgyTYMAnblX/NjRC356QH0yB0ikyLTNAuEWFuKZeGcQvKjCt2rsuCyZo13
An9LvNJB4pLPbfqPAFUJOguibszB65kUhqJDExY3aNdR+lX/K3Lf8SbbuN1v
qj5TOUsUusYfy3Ar9/eTrCW9ljUK0rml3UbXD2F8AZSitxzqYxLMO+5JUvPf
t4g56IlnxLbQHweMIfPFJ9wgriLRORcCNT3ga+tZVlNPIMIwjhFBkrdq18ta
hVcDST5TUvRrCohscntydE56Pua8kXW7uRJS+4dOEc9ecLf24ceQgGoySl2h
B7f5D3pHd2/OPXZQtwr8Zw2Ai+/60rgprjYJlZHl4C9yEq2ijdct/dQzDRqO
9YgycfERK/7D7QWRhHHeBaGqQTBFzmdrpRWgvfNae6xIfbgDThDNkHfpZC4l
J6wMRaXiuViiB/9hmGMvwnJm1ltUrQBfPN2XEaIt0ytfxKnjcUR/aPd91Jrn
vGdsht/QTXsO6F9SIBaB/MldQdQ9CWSILRSt+qyOAMrhNFJscZhHZAH7RJUZ
SGdDbGZUwwP1+dQY4SsoBGipOVlnQBVppfFdB7WxXeMwfwMbm5tOejARoPK5
4wHtFTxhX8XdSxnkL7x2MW/FXf0ArEgfx5oj3LPYXh9z8vWtt0X8w/SCmzka
FzZOQ5BfqgI8sDcNTbAidacfVFvek4mdosiXMkf7uSezR+lbow3n8nV3CHLf
T2HD7el2Gt0v8YGKp8qDhOJQ8xREaWy5m9fCwCzfcteeCX6VafsDLc5JmOXC
z4HAJGsrH6GdeIpQfdoWm4JuLhDJ+LgI+awYhXFSNzbhKmZ8ffeD7rZ20Bh/
UVKT1PHbU5S9Ww/C9WJ790+jf/91EtwETDVACWGPMKQxEQt+Fru0UgoEmzNz
R8JZUOqul1hslPiwzOv7lfzs6SlfjE5dNKZ2ldhHwtn7AFth23Qvla9L0Rql
HHtEPLlInICrM7cHawKRzy5f0NSE3uCPKgw+08hah1wSLRWpZhrLuGOmDcMw
YMQtctP21ynU5m8Qjs+SUtGG+iJsgWto/qBKemSS1RzJKSsgJLrOU1yR+xC8
Rbt3UCQwdg0IQ3kdLhXbJFL2Yl1zNVtkPb2R5+I51OIDs9cHDZx3sm1yea0M
hc6gFgzDAnd13eqtw7Bqa0cLFm8HuE6C6NgabrKKWD1e4CWDgQKZEjRboVKs
WK+36dlpDeLV05QpW8sigb3Iwr2gg8XOwNqLkZUOE/SV8vA9vhPqRieD1sEa
3TO7h73xHRQVqeRXrByW8UoJkFjapxa1yxlTQsT2wLSxRcsGIFlaBm9i4hsh
NuZ0YenrPGu5sDyZqorlCiVJuhDWoQs5nb46o95XETrUS3ixIsZZFCRCNZyz
kldxgFGd1CbPSnacoxQafnFQMNBPPg5zBRAy5BU8dUBIbbOqzBeJuPBd/sCc
W5dSqbNtiko2AEHcOh56aNY7ImtSHB+Hn0vxq4iJjbeAsUNFiPlYGYO2NiRh
WARX9s1eFAN0gd158+W1aCH89PeDwdIls1GTrWtEDbWiazvdPl8ngOPCFa2C
7I4JpFxjGEdx33XMcBlibUCp2AJX9mZXY7XHjmkK3oOgJHSSRqIjyYAc3gZx
T9hohupHanzEiZugpQcdrd0tlEQE2q4qXjHXz1Q6x9gLhX4iLLCy+TmFUWFW
h0OgtNcerxNXLcxyUG18OdHA3USCdwLi6T5w4pt4E+vx8n//wHWA2IWyxOBA
2djn9qrawCXV79Lj3LlzHGG/+DSzAzmXknagBDDULVDHGLFNzz21cE67xrGt
GVuZx123QdxkIIL8fEPdYLBwByJxkLaVZcmVhmPHJID7Ma76I+M1NqqthXev
Xe2A7sNse/H2Btkc6g8nT5+ZLR5n87x8QWotUkqM1E9/rFl91gyB4r6x/UDZ
uRNPX3mqmmjsDOLxPB1ggrqabu+QG2chfaLW84SQQmzZPMA/WnY2Day0zVFV
nu6KKyeyLaQe+lFt8Q9AVI1Wv7dkZp+NHv0ltxPAsmwDMDgDhrHUwwxt0rg+
ivTCvhlxp3rWq4gMPLTb1qAR/R3H9BTYSADKeuhjYPUsWSri8YTLlTJBwQUL
PQTQDQp6IWm9SdQ1d0+yHHzjPmwIDOCNR67iL1i+/pegXugUWWMI8HnPbMwU
g/1AjfootyNdHHBnJgyOtiuypDrralWvj5So5Solp6rkrGgAbAStGUPZ0H0y
DfEmkdPhPvbr1vQXua5gMONW4+FlleHeMKG50LHP8sgjI73kiNacE/58YBHz
8nJ8YAodQMzQdCbUY/bib6vKHX6r69EnknqIxDppRG3KxlLXzKujL0GZysSX
mdbt2mMILth0mY2MAQ5T2CY85h9yWHrXMxeZDCQcyB/bbRhTPJBoh7u6QykG
iKW+1cgbAR0Dnlx52rTVBJybRs0M5qOBrKXlEpv4WQhtu4AuL5yOIUfVsTv8
gndP72tJ2pEbw8L2MJsRyN2siXOsJ6v2Pt8MqXDTLW+LSRTzTCdai4be0b1y
O+JoqNrY8C4/KycnEW4h/iy0TjcP4UFF3hTGK2Brh/D9zzvony+szX8pyJAE
Xhp8DjQC0acc9jB7WoUaItDOjNI67Md4dqKl0Hj9AteLAddRtPeIazIOh8Or
sKua7p4vg/wfUYUvk578Ar29smSVUdMa2/XLm/wg+s+GdXcmjNvkLkIQ0hFb
mk+99uOOQPFqSwJ03WlR4vDw4cNQ8QOuMwCTso1pFg3m6LceBuDrAsEJjNQR
6EUCTR9eO0zTZePm2ltb6wjhVvm4Tg7nKkJ4V4SwxNOKwcQg5mpbns1hpEC9
AB3bCpP3qrwvGzBWLb7omW9rvTdHcPZAbCHu6YWqJCFIqOu4Clti2ygWKJcu
o0c6PAjBrnJoreaKt7Z7jVcQTza9ZGxmZo2rvAys0QroK4xrhtiAVaOCI+PP
AeRYnTCKR2d5UE7eifPB/BFI4Lnh7Qg4zMh3itS7yg216czVgEAUNnim2wJ5
/sTuMX9hn9b4zyFuDaUwUNMDi0g1g00V/cdoJO7UfRxPRVYwA7KXIfNK7uXn
1iQZ3s6a0uKNa6C37k4QZx92G7/M+IXQye0i1awmcgZCZs3QPXTmvt15QQWl
SibFijbKAznchhJpakSS6M17IvudkY0HRGslfSkfeX04Pa/1PKlJ/NvtdUD+
W+LNQoBgPR9yPe+4CSdVBNJx3xBixHpK644raLCUs2XoyofgcYPPZIRRo0M0
HmgfjO6Ir+g90jVQwtBMY3HXYPW+EFk/UJx0F+GbsBh7T54x240khoj6tJe8
9+nO18anAfQmKouIMZf8KGbPf5eexYEXdclTSF77TkSDmDZBra8uMpnX2ryp
VSeBzljlUU6TjxaZwLY3/6BdmIKqETxDbrR4kppPKvkg3wYMXW9epFS++uiZ
4CQ/+VY6wiUCWArUbOLJhVvR4RV8DLCF3FoqU16CNUz/RoagMZh5yiRgOyzG
kbKo/EXqMKLXoku5YCNjncgsgSzyssOrqo/xPmbAv2Dvhan7DU2pBygoGEp+
x2CYAI24R5UxQL99FHRAOZ82lpNEBCwmnL32E794wDiurCO7V2S3pghbll88
hUEi1SbtGU7ZhEv2pUeoKWK+dQoHvJTpqjSW7c6tiud0WyykDkfT8yvCmOG0
cJZxmaXV+31SNarpFhJxYBNYUjTHax7Sj/C6znPWqyptND0MUKjqB6EE6FqU
PeRqVmDqTZVkRxPHW8SsT3drYlgObecRw/qQj8CJsjWr3HE916RTPqlQxwNw
e9Kl13pGTVkjiXn1R0ywYYnap4k+i/dBC+lxh3mLH640EhEYyEBkclG6VfKx
0e7+Xb+XhAWSkQZ67oW/QXCuJyBOihWyBx58sOHJM4N7eW+uQ4H2sYLbug9+
ow894sXLtTx2TmjLpJB8OZgCkCBxxCV5bSIZNl0jkUlluJmWicCjIPAkFdOR
WJLCUiYdCPAtVYJ9JXJEVKYT7NLjutbVc4VJnfaxV11FvdAEc5p+oCQWCdh8
4LBxuKbXtyYztynNp6sY4FBMmdB9QsVRs6hpkQIHhaSJW6Y4DzN/lNjHRvcX
F96ofORl8g0KK2chfsnNJcRuk6367vip13PQZ7WHX3rGfD/mmeErEtlXnBq8
RoNioXn6YzW5hMsQ9TK6yPGVhY3cJW+MSeldYZZdUbzxndJIorrr7c4xkdnM
acwZbpOTLjfQIRshe+LVp6s/jZWuXA2DfSBhzonswsH5EhLsv4RmlfcDSk0m
H5r4B1z5oDSeXBnB3qyOJyWHGdtBVwUMorCJ+kzTQOgBZLhfZlkHtTSVh2hs
8S5XFU54iRy0lwRlIWcAB8u5RFIK8SfuCxzNH5IiRpWXC6iE6qlGGP+V1+Vo
SVHLB9SSnfkOPLDSEtTz+tiOmFaWWt03DNrIoh4+D237Ylx4FfsGSiuOchNS
091HbSgCNGEkSMSRuRs+UIc6NiKWqZB0WidAnHQNaLwX1vY+p9AmwcBu59CT
WObBdmWNptVIyuTnCFBeu10E2b6PeaHG90wZkE3rsrXBTrarGPJSv3L7LSLH
GAjJOElBDq1YQtxW33hHvlNiT25TdPl4s4Hl1q71vruQTcf8WZyUdY3VPV8U
kKkiXa//zi6kq4AZ8dpJp7MgTOnN8Xl9y0NwjvSl82+PiC2s0cxXXA477dyb
iyAmoF7A6i55BT/sb+IuUwKT0Oxp6zUtkFbfDOCOibOlmgu3APe9LAYMZ3O6
9LsY6ytVW83F0YtkgBVg2sTbUo2IYWjiHPxckiEvMUhpsCdX4XePEiTmDuFY
RW30WQ1AIB257LGHh630zM5uPUqpWcNpG5UktuHSKNF56GrS6oZ9O47hKbnu
3m6acrW+0eeleaWvx8yw+/whN5tww4ZitR62xwIgij7qHUi8fahGn/wO3GbZ
xtxNFR/VgHWeq1dGoYKnXR9kcc9UsFcM34m7wECButFBJJso3lAMKY8iJQnM
Kl/5ukEiQbXdu93qz3rgE744/A8AbFYCdvKIE7ItqlVQLxiA7WLsHV2kDn7+
da2d/f+8Pr688PrC6KcFLZ24zV0OpEoS50PxZdVi7yBotO3iJp/wjDQ3nuIK
89NFEyYK65OjYb4Vahh86rq+PNiekkbIUOgmWgBMCES/n/tJcuCEaTybayF8
eWpvSC42r9C/W7OEfuNSfJv0iqt/Twp53wgXPxq3JQq1ebO6Gd/Tk6hMh6Kj
sD7DV9JTdcY97jpzXjdShkecNSZVdW43uttsCqntH4moFwBqoARNDI3tGyd6
VZ5z3utXx/O8N+TghHS/AeALjOeCWKGOG6EoW0xdt4ylbow82NrH0fzRfcQI
3aZtfVtyFzVdC7112DPCY/ztTXPhRzg4mfPMOjYmRzolJ+deAilP+EsJJ771
KycLvpj52qBBFaJiA1rCP11IgAnvwPbXNL+W0tT+n0eOHf/QQicZj+6W19hf
wfM3x+03/lQXLdXcWY8ACUpIRP3+LHmg4UAdUCzsj+/kkAkcj1RlN8y+yjTY
gBcqQVjE5tWwyA6mAxO9FlDDAwWDF0aj+sBL3OvhGPK6tP2Hv7iXfUS05VWI
hSWZ5A7IfsYYSX9B/GwF+1WqM4lc07J/NbdIQeAuRYyY9MiRYYpJgT6Vg3iO
FFn6pflAoOpsjVVhNCuJrOGUGVhW7NlUZg6pOYXWeaVhm6gIADe/wrcGVyLt
/Z8FaHfftQX6UCNQdVGkOeAvhJVeZjwlqi0RQ3LTGAycSXRSekCv7dah+ZKu
Nbfpq6yaCS/2NDx6SAo0jXY8WHcEFVlAWKLdIj6LjuSY16g59YIyHyvnzful
/hSRGSKODehMUfIyZTNoyBuOgDvnqdpstRkLu+GpugXoC20zmi0LQzQx/wYq
lG9QrI9nizLX36MJR77e8VDOvv6Sfv/u0w64bInX1/lVVNyGVQpvzgdG71/1
D7n27xCqHwDDxrGjmjCO0BpGC2wvGx1HioHEWhQJVxybxX8W5LreQQm6NDP5
etZuqz8u4DJV2WLpbYq/HnylHTJ1T8XoLo6DqeB/BwXWrQ1bEgx/FSfCJ3c2
Ze3DSS/ukpZjJIXVuGStSVAE1aQwU7j2Y2nZ/7RLXQEyzUdrDR70PuM7rEXQ
/h2eRQJtWOluatbTOBifmmqY4+FWH8N51iaIzKdllZnXu65JiHbOpZm1mM4e
yuuJTau8M+HV/WNTOXLo3TTFsW0aiHU3bdlKMoqZlNnHky9bxfKfqbYCD9MJ
PmDWSebTVKbuVtsZ+ZTx9tF6B4voixc8d62h3MlBG4+OuZq2aELHOBMEPrZl
Ys7DVPkgbLgppvvIOY8b3LPGx118iunPLRfHh4er/A3rqr5T722FXDIRWyjX
tOVX4OwTS5/mz8raGIVl3+m0mFSl90dcwFT6/97KGpkkm0njvnT4sS1ymCmy
pdG3oCo9BtksmZIixGLMwaNDAqJbj9/ANBZCNyl9QqNoEYg4DNWR4b6ibgEF
2UnW8zPcrQ2i0yE/AnXEHzUh6T17R3MwfQnMi8oJBI8M5d1Rt5na07MeRLjC
iZTZOghmdYO103xJ/+vm4SjxZHrtaFTtGF5dfk3tsuc0MIrZu7bL5wblo+tc
QbpjiGmdkyFNwRdKFNHkYKqqcADcqIiKAFIKuSW631H5kF5hPKpEqaa+08U7
brJ0jAvH4dfgexjVkq3wiLUKFSDvy3yy++gFBpCgikmAhOWvefy7GWeAnXFc
vADL5+uRmNh1nln94ca8x/skNDJgzllVGlrUcSsq9c8wL/mANpDqF8tqD+dr
8wUYDIjz4tgyeYtB4MNeC+Sn0zJOrcwHCH8DE0w0PgIVE86EZstzAPRhSF3I
swQkClOsTPurZ99xhKs0LKKRX3izMBkczWol/5AxZ5ySGaa9k4fUSwTy9ChW
bKaQUHFLKnWXBhnOi8UMAP3dMGTElBsbDpWwqVZ8MU4ExFPd1sGxJfQywE4v
OORAAhkvriPrmGuhbATBAsX+2NQ7GL/C883gJsFQ4aATvBT3Vf4zXFhkk2Ah
73VWlePZlEX2UmmqzUq4vpWzZJLjDlg2V7fGpwgt2ENsC+ej6HzjiLHOSL2Z
Ayt4PUXv2osSHKg4yAODeZI3m6IlhvVineytCoeG8MqwYQW9LkSfgPH8XKtD
HstRTP6AXOx1K4OFqt7H72x3sjDkrTFojhB+H3BfWzpp0cr6TwEPq077c+ke
ZfccUVp8OJJX5eCtCpW4SuT6DWY0/0RH5PrfCXu/ObX+YRtMqfFGzRjBhk9J
Bsr6LkCSkhm2JdVWjh/jZbFW0xmWsc5GCjZTBaqc74hqC5bfjmqpZJwjhcku
7qcLdjYFxQit1G+DKAL+5mF+5PRQTdnMAwUXRB17Raj5h8Wxjz+f1uA42Cbn
zgeEDKqVYJPOm3PQ9ohKtcR95NePZknO9icMQvjj6neSr12cvlmLEjFCVt4N
6zYwBJben95Fbaz0acMla/l2hhQWLpBGa17VLFEpv+n/5JhjnDpcK6zeMS2l
OJWJMnl8EABTqzbFszBP6hotaDXXpdnxpDIBFUbWacAAC1FWZmvg3FhkNPiG
/UOm7doRkNj48TyD8X3VnlXZlEZlzzLZ18gpwF16ldqpU7SBsK99rbaEFBf8
c+DVae6gXx5QlcHWaHN0ltzzfuYClyS/P2GetYKcUMdfttVFAmc0i8S/67DZ
JASedHxAyzSnaDkF13/O9uNEx/bdu6g5BrB9sDc0wSR9p0RkWzxskP7UB4m8
62S6D8k+mFq/Djy3XcLiuEU6EO7vCSX19hmTjQt+Rx06xVJgYl/ZJwpNn85w
GxjKzEn6P5n3yQbdVglyNLgRYCnTOxXHa4oWfElKazly0I8KJ+ACbL+zrWDQ
7+hR5TFJvLqjDmqIuRJArtL4kvR5EWjjhBgWwi5dNU0qmoL1I6Emi+TW9iRt
w88f2vdpMvxunpdb4FjkXKsxJMxp03jXC9b/rKxhmFxs39iZ96zWhsBVKjos
/rGQWwdjFmW5mtP/ogKtGwNQtY7/Hd05tdFDbag9duahqRkFq4CiqQ6+6mbG
yGi8TQEnXr8EtH1bzWXyvijkCXIu3ojBCojELen4998WeXemCRgbvLYGribO
SM9hfYmftEtahI8fLNLURbCig4rOwe4eQZbIYUoRWOdLSDRxE8ux0GdDYHNb
hYoUrGDv5GTc347Ht4RBxfOxGS0B+r73aaGoNN95oVhfcLgcjL1RoeZVbyt9
zB6FMQkSlmNEEPMvoI/gSvgu9A+8X+naDe0grOK4sr9R7J/4iHhIAl7S1lC1
N7t6bQ+oBQDe38SC9G2506/jxBsjgSy9rqV1kgNB+bULqLcmzLIgUOXbNH89
NfgVwS6R6ZrBuwdBEabcQUO0ZRTnUuBp+8I4nL4t8rK1V0O7emfaiimRmQXc
QjwqWZh3ZTR+E21FQejFLgxNUfcqb3j7RqWxL6kukEluj2tTKT3GpiOXoAk8
HYGdfLoUnedoIuUhaRur8TQLaYqzng7Zq+aKDYaxXw3l4JisZNS0vfsxSJ2P
Q/AUygCpvklja/OnLvhZ6R4I3cqYiQwukzuKQRaTHv4ZobEJJ0KvkpFdsNa6
vvqBVeHyF0oGN8DcO9X20rZuDQoNOfPsUZYfAC0P6FHhRTYTIJCuQi5F+Jc5
KkfPc4k/MyJ04B61nbvzZKrsQrStlTMN4f8dCGM1vmFdsp1uf0VthEsgp+cM
5ByCiBvSSxD3BOP5xPiK13EZFC0ITv1ejk/5nF0H0SZkEEgJH2jOeHoQviEs
h+RVcnYPRGkDywD/ixv0lBbVkH6aLZPTsfGxlS2GMCYMDNt554YAt4OETTSr
raOXm4fcv4+1m75zAcmqWNZQHvdMz5P3MRrXXBiyHCPLOw2Jy8dCVHf0Hudr
KpS2hoDu3dQGW07z7ZMveEOsxij0iSC58wyF2ZZC4oP11Zltng1T3jYbX3fs
H7P2XP5wRIcvClFHYav/KDJ5Ox8ZLBhcUI3XqLbVcUeibWZRJBhsBnNNGkNO
V1GB3F4IrZ3G/m8TeoWQB/TjApymF3YOTPi7Ckjj0tcXkj0qTup5qsGRhRjG
kN2sQPHwcJheiYnmafx9IsjC1M7jRNKM4YhtA9Wg0iI29pJ72heQ6bBMWa8I
lci3RYLJ+/P9l1u3DIxtoqK+KcT2s23ixe+xmRkv6OUdbXG8t5Twj/ZZCXrr
rDJaMMRuhSrk5QfuYV06BD5xnAxYFhYL+ZXqBhQ05ygCxalA+hKoECMHTJL9
Yh5FVq9+RuW8jeFWrxCUNj6Z04PanTwN0Li+HQdEHtO/ptqZhy0C5dynP4BS
J0tnoxa0HEgEPC/kpXjYPx0GEapRZEDByJE2QIAfPXRd1gYhQTNFIJ2wtSBB
9RTMD7BKrfQY1HDSwdfhE74Ojjs8HbyYrLy93b/DOsJYxVnwUShGr8MBQwfl
q8ZlKiJn9L0jsSJldZK+bh1T2R/GoN8jK7rl3tZ+qUWGWLz3k1bNmz1Z3AZQ
WhmCyygNhmt/2dNXb/94N8YNZKgxpYOLEdQKslkNc77N7D/p2xmn46NTKiyD
eK+qFcbSdilhJ92nxL5N4MdzOFucwimziZkJIR3oOdjnRelC2bsQDfyrvlZK
Aag5gFRnEmeFXa8moWj1RQozGO1uH53IztvwC5BNqgH5koFmfRbfoqN7xMZU
suIonEbyHRUgLW83C/wpFz66rjw9B3ynqO1QVKfXkGkwOu5TeKXlwOLhemJC
k1cSiKVEQi7245f/F+4hRtXh6X2Jb3AUaSfgvETq6O9XHWML020nglgfpXwm
1SOuGUU9zvPupHTQSuVBDS98hLwzcg9cPPkbCcLSbtBFVxxhyxMe/aVO9pYY
gvdNDRAA2dP8iQ5JrSmlQQjLC/ZHHzoaUofwgjuRdC+jCoK9bru8vcqGPdlY
6fIBHFCSjRF6llLi19+78/5QQeqAdjgwNzvFIblWV+pzHzisd0DPErlez9he
ANFCxN8/gmWki5q2rGuwSCaIEBSsjnJw3FHHOWCOcixXndxmJZxxLFNObiBg
e4Gf0uwpO2o1rDhAZXtNUPTGF1umEXEGRUJ9qDl6ecrgOxFzv4CHU3b0eyV9
mWLng0VVVzfWs+wWkNTybrv4+Yig2A2fV2hdC5fupPdsrqzR7b1hfh+45B4K
QEzfljvzy3I2Ia5UZtyZKXUXK2zYnil62XZMiUXkSu4WwsFYX4yZE7Esv7fY
yRK6oyvQ2yz9tmoCCqcX+pRa7HK9kQAl3k/8OFSbGO51ArtCVYH31KtPJQEZ
JXOU2lQRA9C2+biNwJTw8DRuqlo1TfYZDhjFSlMar3GmRlvVPT60Us44EBUv
tUHcpJG2OEVtxB8oFb9pvGvQIQksjvTE6/A91Rg8ZLM6P5pyHMEXANX0n7SC
Noeiu+lGnepak5JtkAHTXFKXN+YsBWBdNg8Rjy6jiStWxiaBDGGjWbI6/OKP
GMlxjhZYHHEk1Ul+zE8i4bV5Ddob94jFntYWW1RRiBj6JDy/rhKVqWZUCZJT
kslSmP6MGY9Yb0Zhxcm6uoCwL0TsbIuJRkr8QLywQFtR1xBIUzdFT8j31+DT
Z/N4JDTQkAThci30r03DrvQ91eyFrmMsbIyNhwdNHVFKViJBF5r5goQQtN5d
lEMpLCxUPfNnm3s+DzGvfSHT66zHNUK3cv/hryb/xe2FG6ANCUoRazcgLstO
YjQSSOh9Azu0JPhgEMT89bX2Tn81HZ6iqHTyrnCtgZ6q0Gvwrbs78c0fr6R+
a+ikgLazJ1QvFaq2ePWWn8UXZChXQMIYnVdFleSp6ijIOWf2MKkjUlgGxQpk
K36zGKne7cgU1rshsr+vQmO4PTlc2W4KYXORkRsee/vJvPIGUu8WAFfzGI8/
XP1JfmkTMM7P1jahWTRCYHZYVb8OEoPqXJ8Ga3TlcGdVDGiug/pRZiDbWufk
2RZ1jU5X4iAYSDgEjLG0XFVVeE+MlC+yFDSMOTrePDgJeL+oLe/hpMV9CEeO
5+VjmmM7K/J1x5JfpVn9s5aLcAVn1XoVmB0UhtQk5PXCGu9DpNHtFOSBBXym
Cvck3abu1ifKEpwD6dDlWQmmNMKtfZkZFE5Xoat6wKgIUPqclUnOHATeCdyS
R7ugU6fUNGknQLNPVM5LuwAnkoJK53D3B5bnOduwJ9+NkSiT9VOtD/RXPQf9
lNwFX8+hijrfLtP2CT/U9PqyG1QFaA9NGt8py//uLNx8bP/sXKOZ+zTjx9Ac
mijRe4tkDOHkYmntiumhjQESVXIWiUw0NEjGr1xeiYqhsfVng008Yq46+SVk
4383xCbc6gac8yGZrcy+2D/5ned0x9aeVuherUgG/MVxe8TvYMMlW7R6Xpjc
LyWfQGrAvLJe7ai6YxGRZT9GYDtMvEBSMppfJx5NUf2JQ5un42iWey+sJcy1
IIDQyrnCq1jq+t17Pffs07eFa8H6YIicCHjAuUjl6mJ19XTzcKDhFwyXHSsf
rXqbjI3reXpXSEg28LD/qpOvCLvjWnCBxnTODkaoBRuusBzp3AS9pqRp0H9/
IMA/gww4hSCVdKKMw6dnLjPhFSPX5+fxXTbRPz1t5AFDLMBzk0EPpbZ0NOBn
eGZ0szaV9YZvgHlg6pX9CIdPn3XPo6uzHEh7nVrtsHNB5PuLdzrUljTv2oCC
jTEFXHaeAkRLu61LeNUHbqQzSoIyD1gPMCKxC96W6GVmXvqrFDIiPBQ9o0f6
ZLizl3Z+TQRdhkvkyOY+sUvurOWDiFLa5vcTqXc8VsgjPN1dwlT+LOpaj9I5
nK+sdH6CtmV0v6l+/91JwIf/gMfsB3ky3TKw2sfAqpZbF6EwxKzVHvmyqYz0
wBwn/mm2sTOTuIn5ELempjY+cXCARKQ3oaheNezmgx8WMGf0dBW+b1NMmX6q
OhkMjs+uJn00SvV+k8Bp5tWUs3TCufZ0MjPZtGqNSc33emgfriHUtFZjRgUQ
7u8vtmDiK2SgVblLCF3V6xxXGOXkEEXlc5itmANerV0PMCgaiRs730Ph1fAo
Gdk89UNokbL38hU5Y8DV3371GBEi9Z4weG+ilTvk0ybSGVSEZJ7cdsf3c1bw
rYDXsBvzV5g7gq1sORc3COWWC7OU1J7L5YjEj/UShCmdkdOQ6gdphdcGrQG9
v6EjWPxEXcWgv14h2GU5WV5RZSOrSVdJSxx+2Yf2XYIh42mxKBNuNdgByO9f
lw+FVQ2Pk7iWL56h17dvOZPB2tMk/TUFBV52exHkenHqng9NfT5Bq68/dnmh
GUSpsM7pOJYCG/TooAkOCXHMeFtJHrxjpKsXfwuRLDRUkbndheS9dSkQJYTb
KbDxGOf8XpC9SqWTCUJ7WrpiylAHmX9HvtCQoazReEKCOaDTPTf2iJTlKGQG
oF0LJUD6rXnOHjb84zKqllZq8mrE42zJjRn6sYxJKLnbKDU5XB0xXPzVfjKP
tpnrp6VHkx5yuo0m2sBku1O55Ae9acVZUn6cnqMUQCt4a513wlWGP46Gd6Q7
1s6t6L9EE8OMEu4/dGCp3ZZU7AwpKSn+hB/qeLEgm+ZlEFGLeC6q61cs69Cw
2p7HzrTFEcB3UaoJD0GyJO5De6Z5CxiwgjoxGbr91alnlJWi0kOKK7V6TQgh
Oy9yNjQtu7KE8apuF+Y3DBpUzLXkC7bCjGt0P9XS8NYOu2/GOx6YQoqnxGkl
74R+XxV23zorHw16i0nVpftxXbsRc2/JlmrMQNQzXEcB4UU+bSerKoj8X8ub
Tt96ZW3JEhVjvgo+sCUHX40a6fZ/xtjn/MBmslSK7Hy2d/hD5Dx+vYWh4a+d
FEDNsVodK9gS6yaoBdwkvXLe5EXuG1QoASyg6OD/wGyVPztfGQCqLC83vFE/
VAVIAN8bi195M8b8P8ZILHQ2ySEad/WcuWENlJ/hw6F3Ogn8WXWLqojc7VMt
LmtRd2G0xAcw9VGHncg0aESzfG26P34MCxgpAE0tpY5uipLm2pRenCM7Oi1Q
gYKBhGBYODZOcOhIdyuc553cWbbkVhu90oRw3YrBXf21oW7AkSBhwATJIVEl
WOtlr8s2pfETzfk5R6GoiG34MygLvwNmZNM91zecVtENYXST2GM+HKCusK8B
1ophLYbVQesf2Z9KNFdyOHq50HeScwYd/MYfecLqwgL82wskEXWagTwpAHyY
z2v97Tkvf4ui3KkeKxBHYxjZiJ7YZMYoqXXRnyfrObUHij6UyZDuvNU+DdfN
jvhStFXruscLfRVk4ZHSJ5ctn/4/OsCUae2CdNyUEMjfrhLOGRKNWWVixAKl
7kUXe1ymnR7KlYIfFXKKCW6HlXXy/cSigye6F0Up1HzzZYPvqmKGI0CSMJo1
47jd55oT1HPaMIRoPf+D0Ldit2YO8Epiqm2tSkRj8KRqc5kdcHIuNBdBXS/a
4+UqXl67XnYXKMW8MUOMRtDnJymr2qmmoW3o+Nx6X+K9Q4+M9rJ3zMMgzbWM
q3gMbperimov8IzeFpwd7SdBuQwnOrc3hzXvF6PZ5Wa8jf0b5h4QSwJWMhfA
B1Nr0PuQaxHRQH7661tq/u7/Ttczj3Dp1Wnl6f85/hEluLz97Tdgmqpz2+VV
5KmqiOwfBXxEY/Owja1COJYXA0YK9mtXXgR7vTcAYOPUAs5K7sH2kDzwhWCZ
xK+mHBba1LXFv2Z4R57I8jIojzABxeBQD+wZTngyaLdngzBr/qVAQiNm19bA
UgiGgiT3h3HUAY9C6QUHpwtXnAu0tRCKh9lzORzHUXVzqvaplMUreRyuajoZ
+dV4gR/wL23ZKsnNZNJuLrON5EUkvd07jy9xV/ZbN07HzkEd4qAJJT1QovpH
IeoTBOl0unx6CKqkF+WG9Rjn6pJslpQaREIGUAJf4YCiQihFMCeWw9/E3m6t
OHt7uYOzpQDrlEogXEn81m3NyNvUhUHV4OcQQuxs8l6ST+Wh/LwETX09iWvn
waiGbaYCduH9umkQZ2l+g0TKvB1BL0LY+kkSSU3C+XofV4d2hNWBylG+oDsT
J5YQ3Q+y9M73EJqEII5g2EF7hdKbP0LhjWpTgJS9KlgXL1td6GY569c0rHIe
ipQuNO78PXaGW0BULlmqF8dIhnDV2puJt02Vjf8fZ6MT1kvQuZuWC6+CXs35
EODUB31xIWKKQ1NHxepoTh/yLdD2dyuC330/o9/ifUkt8Kwoevqw3IV3kfRK
U3TJoWbn3Dew3DkBcDvFT9eEX2Cqb1BoCjSdcfT3iWANs1t3iRuCrfuio2s4
nEyQaQ34SOK2ZqnKt1N0XwDkzCLFlMqdAfP5hnWYzgAI3CLfTAQNAkchOuoB
GVAYyZ7HOPoTFDT1otL9dtPUVS9i2LL2zcFrrUdAjYXQ0PCt5zK0P/BzzEZD
XBXIbZ3bccsDsgjW9WaD4TBmZdkeqxqgswKMOk5XLvhHPRxnC0VDNy7Xb8mw
C9Fmxw4rr+SUp05nbO0ELoAywJi4SDZpuThzF5ZXoV4g+q36E0pdj2qTc52+
adLX5ixXwEK9PkmGXyZRHFEkDD4Qailbp0boDJKCFi+a16yLG+AhrROBZBqS
RESTmy6sN+PHN1A/z69DMz0yp/IK/wPhYwudKumqvRhIUE2PAlLbQwxGsHAr
VrjO8wAaFTGwjVXl6ik3+sU+MivxuoqSr/w0dXW8yjydVF6+1um2dtDGqfFN
xUSKofQo9AlmonzqtxAydGpz8wU806mj6kcQXavj46IN/MVBeOa67dVKVGSn
ECRUN4z0MvsRUa72M0HceDkwWdGGktU1Dh3uc/BJOmgZGrVBlL2hFHfB3DY3
pIBzVycR814CpooFWt7mAgiRBCz2oer++R6GGvrUhCeMmo4HfDji88bDaH38
ICVhjFrVtF3RX5m0ezTSkBn78WXpxacNt4JxPrg3aQh34VMWms7d9HCv+71W
bi8AeNA2gsw7Z9ghOz5/n4NRCcb+HRLs2foxo3ur/1rajvC8PV6JyfsnPxIb
u3cWTcVzpamhSbJIu7I14vbMyGgYC/akKh4zx6xYtkkVQF/kgyZjTxgpD40g
syD1ZKcXfDuoAYm366p3hVyqXQdhVHbU0sbnp8QJMh/EuAuXTMabrXLjXfOq
HyqfsoiisjFr6LC1fdpWNW1ilOID10r9zE23EjHfDVJl94jBYoDiJVs/OYdu
N65jAccBxDX1HKlI6N7s36ultIE/lRP8trSTW1rC0mfj4MnKF2IMA8Um49vG
YOU5sfRNjKB6TGg6ITl77xp5qjqoE1pZTNjiRFGt7itT9Y55KI+Wmc9gjPX2
nJwdl1zt5qwbq/BrO8MPyHGAQ6bNcbBRrdPPZK8Z9Aw2FFYj8/sDbwlUOwzn
rn96S/bp1EBd/K/PydZzPsupai4z0KqkIEAooMl71Z7NOErBxjMEIjtxIq1Q
srQwunET/ncYPUX4HwsnStX6OT7zHuk3YKdC8rnSIE3kwyxQ53V3kpUl5Y6n
C0DlSUnkd1ZtaCab+6sQOIGmsFtQRO6NuhwjABfPfKJAFx/YyIFOreoqQWif
U8m1bK5QecuDF5bpCbQpEaaRdCjf8OKzH122VFe0b6Rh5z8o7GOAjJrvmAgo
PnbCbP/havxQa9Aa9MVIljYlucSTlMv5W7fp+WQo/uUPMHeL5gnv/fqKl3BT
s/vSWCY3M7L+now9MgEIT/QFUHnTFNaNZMnyr+ezDDiknFrQpxWS+yQy2IRC
tKjk8m34Y4T1PP/vUG5DH1NuOUDkX/rlg2FpIMrZRz3oUkIDAxHkxk37aSHh
dffmKYVxHQTRP/Zn0SjcRhEe9fl/1o+OQ/LwxlA1qDumnMYeI+v4w1LFyyE4
8IvCX74w026zVWnd77ew6WkALwYwy2koeQQUt5dX9WrZ3ZuXijauA4bQNRLr
jqvDY/2OW2w9wnUuIIdkWGbZ+RmSs1udcjENSS0LLtJUDSnvzD3tUuzdXICw
HgSb26Fsx00Wrwojjxb7yThAdxXd+Zf1FriYRJ4Byr3nc9tkFAnT4Xjjp1Wi
idYneH0J+E6IgOQIda1wiC/tcRFOFV1/j2tmQVNcRdjgZNmGoyUtUGXcO/0L
IkfvEVR+6iChb9Ay9ZtIFSJdcZoeLbMnPQlXMOzHfCZQrTpiQrRy6saSvGCW
sRGwX1Vnq8f7aDJYXJg0oOuWrH0J1c57XibKRE/F+rd0tKCzRjQ+CdT7VMZk
NLCDmaPsGymzx3YIL/8NaRnSy/ixZlnOcDcMf212YGm727NUT9ua8rkvEVAp
+PTolN2/zgH0qMQLlsUar0BrQBKJIj5fXqT+Lkc9ceFw880ceD/0/OCvdcKq
rbOsigeWOZ7sr/5a3hvxFAYU6CHX+DS+1Vc9eF74nNPTOwLUbDKXGv/skzrX
7ZSE+oDIxoW0uw6RFMz42LSzuEteApnbdBv0xBXitRoFZTzZXCDD5geU7iYk
EfKngI25JG9bfK/SNreXyfjw7bTnZvqLfDIJAaK096s5323jFcBmZWCe7/Gy
VP3FRDtC3Orkf5YHQksAWDxBLwKf6r5o2qFM/rxNK2z+72w8zBSpmlqqkh+2
1LJnPs6sxq3+lGkFASBPqNJHGPcP0urmJ87tt6yxsaHYeRHZwIyopmUbwgph
MLZ/LdxakaZesu79Ak2Y09AqBehdvV8Pv4QkyNOoApVfX6Xl6Z8WguXpsZR2
15JSppaaHMYuxr2bmnn98ACM/W/rueo22yZ3eFTm8OpqpL9JPrdRDmrlKxZ+
wJ0z2F/IAdkX3ciOyUxk1b/tHA4UKZjMJi7/tAwD5Aq3gaz9wij1YOf9b2Ur
pEWtD4p4950cO+d3irZ2dxhXCWeHXU1CZdeYk7b8EImxzGBrZ0KnO5B2qmty
QKfbk0iv7kYP1ufOzGzWbdQd/uWQI9f5KlJ013n2DJoiXcDwkjIZJhzlisFZ
44O3cBsE7poA1dZNafWM9WRMCOU9dUK1v8B7KHwffLvofqcDvpr6nZCTbfxJ
sJ2HwlLUlXrRD9CuEoCv1s7KqfcI9S2TdwKzz6ZbFn4VgOYMdjDtjRquq4Yu
+GrEYtLazP5LH0hdW1bHuo+RcMWUJrU2gQurrRJ7+zbRbKugPY6g9V7jWBsq
l1ZyVNOWqZ0WptW13q60mgDKXC73z4oRPVc/rZU/Mmo+abaVQnbjQZm/qpZJ
qPPsyUn6LGqkszSNCVnP5bR7mGvkn+EjFGa8K/GTU3HD6j69AEVBEnNZNK3E
zqkvDgLoqjzEozcn3QYAFTo8y16fnlSd40wriHPHMd+HQD5iKbvUBXxcX17M
fhLuawQPAhRgRjjY0t5bbFAQKBw13JWV9oBLj3Earnn12S8kO3gw5dl8vwTx
mEBptPg5cgD1BNhuHZkdAr+9BmJqosi8dK6rQuO86eJZSrAK83Nnwv9ctg7o
4/Resb6a1ozrJ9LFHd4e8sIkjETgcKDHslpzJUOns8XiTKsckZI1CpGJx8ZR
RSUnOyTV8FUcOAPpAh+RiEyiCDgTPnSl00K/scOsN8cQskH59FUwoSY+m6RK
ItIysC3hJnHwV2bFB1eUH2QL9ZroIn25rkQTB2WERMlaslQ2vJoGtySMa+R4
xRBweYUxtFn5Ci9KbbjCSuEq4hY3ltehPfZIr90Boz++Mkm6jzleNeAQa6HE
nHrUhR37fAE9BPTZRvBwekbr3gkfnRJXBqET/MOTz8qojMM4HgpsX6cSpT3t
CQTeKdcsn1l08lopSPBAMs0GoiD1zMC+4Sxkb5uIJompGqiPKmBled7o1tVG
XWnreMCVhIhMa+vV9u9SsIgQOBhOV3gmgLM5KPDZup9xGbZvKBv4YPyUyOiQ
jJq6IsMeFils34j/vJiixuG/GyNiuz45SIIM4kcNf/Cqm3a5Qip95a9KVXp4
XpKmwrqumFiF7JBjbMb+lMrRNeYg3VOZiUdXlTHexq+sowWp2y3auhPEo0Lu
wsbQD+2mQ0mhnwBhpObS6e0j9l5XHSaXAHr2mNuCh6x+JkkgfZmx/cwiCzWm
Vc10vdV9eHbVfOyd/yBH0FjIwoXGZqVrOFaKOS4lTy+VTxnZn2iC9YuPVqEc
j5eCdd+TdEgYJKm+DDDmBAiMKNYWOQA+0Dm77LFiGh01xAO2vvIkIoaP+uXt
HHkumDEXfAvzFZ0uaNAIpVSifJ1NJSmgk761kwgj2wLnkL7+HoHYjUn+4D2F
J4vaHHUjrAtXmnp09gDcXn1+RhgkUjz8wDsNTE+9HUZC0t46ziL4jt9i7b72
iZZqEhkxvI8tEZSyjNq6eJHJbLSjFWjAl2Is05RgZpOiE+LGGDXMWiWIzm9r
6GZ36iQA47IhaQwB3ZtyTChCpg7Wb9I3tTTNSNYty+1MUekWG/AtuRTAuimg
IzropUI6V1ziIZXwwRmfOG0tzRSlzZ0W8ec4qe5/J8WBfrPsPeagE771ie+A
qJuZiBcJnhvg3A+w2TNW+vfhyL1PMQE435deskFbwdYBr+Mh8xf+T8zLsq5y
8pPPzEj/6IXVV8C2lh36hFZeSIMROFAY+YAlQnJOkVINuFZ5YplFrF0enWDc
DLRYdVMFWsWo/yDvBNO12mnh+2IFRMJHwTguXO58K+H4naeEWsrM5lvEjp/a
mylpLqGIOsxv1KVSIuxYKo5wb+XvluS7ks3Ko1+a5lCKq0P0dzJN0Q5kBK/U
GHDjys/FZ06azAGojKuNKDctexpT6860gv2KgIIDsrTd0zZSx6NXbwH+DX1y
ikLFzoT6tZq35KM108egnnY/88MRHzirlkbKB2pOlxtY6+w0LbMrbykGY/OA
lYw65fcHPlh3AIfzBgCBK15QXH57ITwfUuE2hqkn1Bl2NFpaqcX7eYpOVNTv
7DjNlJ3JyXOWiCYHEmQqLen89hSj8wO/l6hrG0iBgZg59DWDm2rbv02okCXQ
mnaMxVQTZjnbN7Ip5TaU1fspVs1L4er5jNEV+0dmwO6aUkJaMivXauFeOy7A
uxoaCrS+B/C6D03p8PmgXm4n4NetvKVAlnafRdIfv3w9pqcoRnBSYAfF18q9
AV1IGVr1NNJNvMaIopwmC2OuZHfv5dCCWLp2NidVUHY6L54Xa3MfPPlBleWI
8Wg5xZn98ukfUlZ9BYaf6v6+fvo1O7qD1K800TU4a/6cj8i8LGMbntgZ6+U7
GVOTqA+y/YnCmVOKXXHQFJ216mfHGP5jIuqYJm7e0QKVSoqNd0u1UAIejwiH
YJaubfQTDBSwhdT+BvWo0Z+rAwtRYz5LBdssMWaY9GSfgbC2FB9vyu0/C+JJ
DWGHHypH5mhPs1PA0eP3YUG2K04BLzpOe1v8c5Muxf3ID7neYyh5nGz2oXJ2
m3s+N1a+exWWfpaysOQIy4FEU6KerSYKMc0iDGVUzXvk2l9HtJ1RoskUP1vn
fgt62Q4KXcOWnP9hALXPC/nGpUqDYd/gVdt5glziSqDz5eeo+qyRFxbVSb0x
RTWrYSmp/H7k7fG9B9i8DSymbhSveaKm/Zw9iMo4lObhEbVApsofPoVlhCnG
oXfhP3y+lXiZ9yeuRxLZgVrSl2nkc8yE/9abFS5FlCOrX6JzoZraL5/+lUy0
816vO0dYxqXeunRMSehXZvKg1GoSsn3nuCByaUf1ZHd/v8MUV7UzEoWkuDHO
zbaaQ/+eG9Z6KsbzIpdimJOCZAhbE6NuhB8SF8lA0cLub+uFpsCX9DpXtbm8
EA1I/N5gF+XfqcROc468a4j83vq9VsqlVyUltCrFeqDqtI7u7inMMhbLRNcx
f9SZN5VYPGXW4Xv4x14G4myOWr+q32AfPAKQeEVJzDNjXNUvhITHVb+iwP4R
2FA3jdHEQO+F6C0wH8ycuPUg6HZqni1bdTffiNBRdzl3z17prQa8QBdraUi7
9VpstOU6ajhTwmWgMXdKtykylNkIUxIPKR6qw1gI0Rk9IaxVks7FEIYMe+8T
MFc2iK05YohcEhe+LEDGzHuami74KjESvUSsVWJPPAKqkNnnZ53duRl2D1ky
jHyDGzU/2CYf9xnSXctFxW4svRO8cP3o8Jii1U0Urj/FKlkEZ/rBjlKffmw5
28UAqhr/U8UxQW636nRuX7lniyWPSxvyjtcB8XbCgdT0yFzbFTMJ7+XUJJ1f
TU/tmpf54LvvdlvD4ZguHYRk7EDgOBx8IqZ3//dOoxhdjjC1gzkwi1cdscx5
TS1kT+IsQ3qXObQraudUs48dSNRjS2jg8LDAATxT34aBrTZYcU2AGQJdY8em
hwGuy1CpAnPngEOaJpoSSDSBL7iMqlafl6+gkmguNPpGIS05+0ueXPp/g0Hn
MGqulJ+Vbz3ya8dyhAYBTpgMuJq7UCNJq7FyyGeg4yOTv/C334k/wZV/phJh
XbE8DZxqEFR+9gkP+JMNiWdMrHk5GBpK3En5lGknUoqk/+IzIIgGDFNSY8Sa
5JExPIVJ1mcmLgT8FN1hOWB+rXv29lCu7ItCnrahxlWLglUaWth+k68q7c/E
VXacaGt7EVwgsb3B8bLEG2++xo7yDxpg9W73r+1loK8JhWH+zKT2dSWMgzAU
PBX6lQ9kUjGY68ZVgqA6Dd+x30JSaeW0ZgU8Qhj6VkoWYJueeiSm6vDhuTjg
vNc/nBMHN+yy74rK2xjT5vHP/k6G/3iTXDh+M4WTnUWzK/N80M8PxY8A2fPo
m//nYi3U7WsqzjdVPtbRpXwhPSvEll6QtXy47xyz/4fx9nQeaQ8jC2AqOyzi
esPMuNyrAmB5vw8s3W2SCbdAyj/6sZbYX6e6z179pnZW8Za205IAaDtP/mDc
CS2R5li5QEn7HOtQGnqeIrJNVMU166Zma7eYPIF1ewo3h7uu8V6+i6SqOnsN
UzmoeyU4xhMESPbA9wwJ+cHVvQIpsaAj8t9CV0xI9XMW6H9+/rH5g7SbKBR8
/m0o0gN5j8JoPiTM2QEzvcksNKup7kbWQBt6RkFxibyoY6agiYH8l4bYD1Dx
Uc43YZyOHmdfI3e2WMQstj4t8Hl4kAnfDD3LzcDammNY3yfK1Ke65wCKjOE5
3gbWI91Geb5rxh2JtBC+nCr7HwBMuq9caXnMpZug2m0z5CisPM+uUZornc7u
FIF52S06lGKTiInnxDM27N/m6eFV+8EvRYjngZxXESRb96DE9rOxexQxlR/i
MytN2265jUwVy4AixTBgbSVN6nZpCLb91ffSmkjkN/TSBWF8GotBVeylfkr4
EBgCW9Tj3MqOxXlTmygx9/kr6kcXV8aytsg6jMxuDcOcc+EL/FFnXAOgnqfL
wL4MxNcBt+rCxa5tDzj01b43dgaQzIB96qzL9gDfHcHQMWyBKsGRUBtTrI2b
iqs24RcInqCk/Kvx5vSBeqVn11MWc8TxchGOQo8L4MlE49EggLw4mmJ59MyT
qhcZwFEyM42n2jwnn/oDKHYrpiBNEzttTOsbYeRZW2Yvsc0Tx1cffJZOUFF+
7cdK1yS+4cRl6dgIDoJYjzvgQC76mwW/mqcusGqabqDisHA/iUse3T1RDA3I
snw9UZW0Q+nGpNOlYQeezM8RwH61j7Iyszsy+IaNSC/7RVwkl90A59UaNXO9
rh2QEaIjrIgPT9U/FaA+BBYQdIElxXo8nQqDKE8yk7dbnUMqizzlJbojZldc
mrJhVrZlIUTGlYncZB+U4FOt0MIiIjoHMOflgUIjjuGwptiuGPNcLShI0Hfz
B+Y1wbN9DSd4MoMyktahHnKyLAxeHuJ4XqZYDq3yZ17Jv3XaUOr07a38gBGr
J/WtyXHi15pPwGlcsLQTb0V6M4YBI/GvlrDiT2+XWxd+WmhGGg4fwHMjKjSy
ukYAykEZIlOq0mcBqNF3rUFe7GwQCyVwuhlG5wjkiodGZF6Y2d3WyZxUqAHV
dBakxL7AxX9jJEazL5+2lQzS1mSCTdx1G2T/Z7oQxiu9u0dj95U9ZUaJFf02
drvaATri+1gaZ3PLqoyuv4B2awb32AJgWR6kEnvZaoYEWKJJnOjObnBtYMSm
gKrMt/9PIOZqN2RYdRKgbUZuRnN+9nO3xuuJYiBgm8eZCdUo/CyM4mS6M8FM
xZYj8eBWlnQ3vCtdZr7rzLjaiFSx3xLXsaaDw6h2Nuy69Zn33D+CWmZLGHNN
ioTp4+79VATxTPwwv7Hl4u/O8E1duTPfTuDwJOudV/hSRn8vX2XwK4ExDZgY
pS9/nxT/XUPkTu//HNHCk74V3B4yG6dHejWKTzJ/GwlIMECr/V/Q2a1VNrBg
XTULe3U14O1DphqUfbRIP8qhp5rZlyDXqmupmjG1IQUqslMHMRzf7IBglkmh
H7mj/zxC8VENVFM4Pp3SSscOC92D5ha2CjSlVzVqqYOmQqWaDihb7qUygsHC
coW5Pko6MPZZ4PBaSjLEY/qdvqs0JB6VjbwmXcu8OOJQM34t3exwAn/H6M5N
gkgwTYNGxAGaCYdGD6tmnY5Uwvm3u0fcqA6bQNXCn/TzwpsqRFJ250Xy5plE
qxdYcvxuQJApeGPrUP9hkMsJjrAy2Zqa+oY/r+/ugtI1tTN0mqpc3PHSckPj
nBBrhdPQ6Nl7Uug9fC7Cg4eS6LWy+R2i9sqTE0gIVrSWsoj3WupdBIAqpjkC
m61tYlZYNsd2wWiMtAYcnsip+d5JXYFfzL6GjgtJpL+6kO6WhgCsGzPPBy9n
6IbCFB0BGpoUTvPbotfQA8YLfNwq2kAxZ9r3T+yOAil3DwxPLvnKsUIsfnY1
VZ/vnM38ope4OsVR4MYB99nZ1JGE6IJsb/tV0D05J4svkaI2gJ64Yka2VrP4
ASSk6WRcO4y9//WLf8E0gq3VJf2HyU9IylP8K4OLSchWKQ4fNvO0e5xn8mmE
PhBWyWym2vb+qCFrj6JYQ9xQqmSObqDdHC3mlyC7quK5uTuEoH9whmCijALz
+nnXzqqRYH7Y71gsd7619UvndZ8BtAxqnLBc2YmhU9nPmrp9k2u1KLimLxH6
YpsPcULGuKYbMTygLhpv4UfKxRUJydwRnSMoSRdexs04rvpYLZxGNeg2wvK0
aqaqjaP9lwVFKsWYIbe+LtBvLsGdAmsxXtpwof9CXiPPaUOHM7KKlMft7Ams
CdlqgAvOAdNY0r78NZ3nVfXQrjfyQqu3p4fSyTsQ7duYblip0w/kKz/CgDFO
qCLqrlNOhBm5lPsL3CTjbJjUfemhN1/2kQ/qAeZpt9weqaSqO5glpoqRO45+
Hy7uRhvBf7uSHBO5oWtAnkrYn637DxCHHGxBE0oXck+5duZyMdj2fApYfCS3
FOGphcztKDMP0gkHtMGPTUzAGZgN0u0Uga3xPQSDYBxvai/Z2AzcUdH3KfG3
+cq2GjftWtlqCMpTswTW+SFj8vL6hvbDU8u0ICQ8ZYxn2/2hYLEtc8ftgE77
dtEOabC5pChS773csUV0asWNFF3gIhOi+Pj9HnRhfnXWPHBpv7h9yH1Jdr/F
4+O0In5a+NGSEL5DpW7INvJFEr9jjltGZMO5q3/bmZBBdjpL+T4qjRLOtVpW
U4pw4YmksYkdb/fCuL+yz3uRIEcdIIHc25JJ5KWXCbdXlZjSsAyUKmmgQfRc
UMUy0kthk7Z+7qa3GUQjJn1z49p8sMnoc2Bpxuvk39jFblRiLACrVVMdp2dg
cdl/eQNhDegNYMP9gja9pUTvWiEeIXrfbvxrwj3eMZe+bNX5AiLNNyq8JeGe
nMRhvrr1DNR7UX1PT+B8iwVe4v/EzywngC842kif9eu1wpcpXXDCVnY4N0bY
mSP3lN19p+cM+3YcSzeV592VYwTg1tPyUW+C8jmgq7mnvujDBgCr1+BtXueN
nxvgbcUOam1H+FuO0qD3kyM/1lZQ6NJ6dpomaXfjvC11RiWKpW1gq+QhENxp
7GfxQueSWNEcMQP0wovda7HHSQtzYPsGFel7ZjbfAnRzfrQUxI6klqfuMum/
YE0G8IJ55qH4vnArir6+dG4iuxFrQXk01jPFAUJBqTuIMqy/HKPYzFJVwMoB
ETqlYzjzdTY4ipI8hPHDxu5zqLAAkaDpDvjXS+KptNA1CM1PPRmrGHD0znaY
NU01quGV8LrghoMlB9/nRGEYbq/tvjGp6lwiF8JfVpR/yn2ApG7dwD/B8aHZ
WPN2nxUSZlM/+Cn6PXErU9xxtIVRoF5vZjrDJe+K5r14oSEs1pyvI4SF2PlD
uHz0c6Tv6hsPNL/klHRAB0iaUsc0GXxgWq+uQq55KI1piiWHObbEXmKoQMZm
cOxGJVVQPBzFc+9ECMUQ6FJsS+KR86HZrPYDC2sKZ1rU2B3vMd+dOqzaZJhZ
Bzzws73zA+kR2zSATeAW+Ow8SzPcsfWU3W3kxO/XTOSJlFZZUqr8CD1N+hE2
WAlpCDCswYj/sy12xrO1/PDGW+XLFIrrwCJC3J3wJHoEfDgXj8GrMgIK6krK
Ec/zDqmsmWskeCxU20F2NZpIVkPL9ja+l14JgKMFV7rnY9pm3+z8shGgduZo
YM6ROFVtkvwOvF0LpWyd6VfU34W/nytJ4bWFHrTStfpELc8gDdGs1SJf9RqK
W9cxN/9bdop5Mg62JqEE1I6In2CmmKQxjEijDJxMHxt+C26vURK4jq1GdM2t
mn6X4ppJ2MtdsChHsqrN1n/isP3T8antvuueZXRhqyVSvO+EVtCUBWUF/cGi
cNXuFT3ZxNQj1yGCy3wHjvgRfEA+Ed5wD5qDph0tBzjpOVM+maO3k3qZbpN2
BTDU9RG8xAKFfUPDQgEsiFlrOMK/bKB2nidpk+YxsZV9OzRp43CLpORvLBhk
1A355dLmAJeMvTHcVQL3S4TsTe4E59g6dWTB0JyBCQJZCJugyv79KynA7jo5
AqzQLhKEwA8TliLcz8jO/LKkW/3obTCYymhu7K7lzIrjk1IQc3JKeHTC5cF+
SIcSWF8mBN5qHlXwg5zkdZkww13P39gce/CRI6ZxCYlNbHuwEAbocL2M7ta3
AVNnWNmlW8/f+VFr6jM+Q7gvmjciyVIzoXF9V/xPq3DjmQYOyfJ9pS0lFdsE
QVnfIcJ/a3VGp2M3afeUBTpWx+tyJYj1W7Boy96Mjj1prphQgDxRAc4q8eL5
CciKBQq7jhzDm25eSGMkk631pibDZhQGI8RJIjaLIZMOkWiw29+mc4XZAuFK
u23TyreITRBU6fnS3YaCPqTaINr5SEQo9K0SYEQCywgH1ig14DU8laoXacha
ycKc2NABo+DNlxGTZeSfL7jVOmU5lAxVehhi2niEEdmkrAanRtRioFoWCzOI
D9lD+rMLByxs17Q9MRI74InIjn2V9QEo+uxqrCJbBxFgJptan+tFwSxf9mp5
lzLQyPPNNvYlYy09UQeri1GC3dLkupHcUQ9ymUPfNPWq01udkeuCzX6wenbV
1cd6iVhuLbEeuKuTL0550Gj5aiPBbztvO5/gGv8jPTtTt9OwE7/DqMyaQLWF
ednvl3OvlO9nFvifddqXkdPCShL1RCYvBLoiJEtvIVErsk3Vl2qYMkBblTSa
uQ1GdIWNzcLSatiDuf7VUzWNi0x00qvjav2SfKiAoEIQF4FKtruYhyP/xYjh
i+l+ehHN8p/bgNrtaKTEv8GZ90s1K54W0XdkC8DsuZam8mR6XVCE9Sm2o7e/
B9a9vjVlUjasCZqP59c4AtvYvE6ZRHagFeR0dvROws9h89cpTWWy2XiZbHsU
u8Df3rRHdZ82Up84+0QK0c50c4O1ekp+xTLDBsnqHhyPJJ02+1PDvHjLoP6L
N1Q0+1qeFo6WXWjaBe7ZPKz6XBeVVAtC37d7basleX2T62hIjFIWCZQc52Dg
is6Ag3DVd6IEhhr56BIl1bSDF7JP4VoAxdsczPhNRe0pZB5dXd3UqoTWAVwq
iBm3DQ7di0LISd9XCcs73d68VwWak5MBfR4AL8RkdD/cfjw2IRwbWb04JDsR
waAMdE4f6TFdoXXkYy/VMMKZfVX9majSoK+R77i6N0VmAogH5olx0zT8AJJ3
lt2fO1vX3E/fEof4+4ljS+thhxOKtAhCHLorTV5BPaPFv/VuFJrNJf/VSY9m
MzElifFqeZ9Wr1jdMDSj8ph1fBzclWgodIa0I4E0hgbO4goOyPWsHoz0w6k7
W9QVoWBBWhRgBxgt6UoO9O4y1ktHCRh09uHe2uywrwEZ3vh0cdO0QxDtY4xR
zJO2GPD3UOpHTSvwdF0j2qJSFLCY1FkIPauh7RLz+ARBqqTTHHYGMK6Ug5xA
VpWOgm2mfh9XDINT8eDyfWHDewWWp8+38EmkwMRXbiY/5M0pgUC7zBW0xB9i
eHRyEZPi74s0Xci/WPbgA0G1sEBsZGJ5jtRit9GiNRO49yRtMRWjiKSWoZ26
v95dKols91PnJb6pcAEEKeXTzUDWBVAjgKT4j5Ceq3raduSKaV3C/hOfn5lN
qAWxzRVpxC750K8Z4lwn2zcAcTrYr3VRoYF/pxiOjIICn9p0/3sqYLng7XpH
E70MAA2IfaBcgz8CkzSEmMZeUXE/aSn+W9N5jk8NpEPEXYUkaoxbVkn+2tnB
RQq/h7ySTHGS5uXqufDwNY63nevB8fVyPGEv5A2AZNwEiYTryiwcuBbE91EQ
nI/yBNoldIHZAQOEOX71I3aOzifGP+qRYHAGAOcZMq+mA0Dbp1VtheBnUYd2
Xcwv5TdMaX3/WugWnbDT6P2lBlF7G57bhgsg/BZJpsSnn4ZAwF12Cr/ciAKv
qsfx7UMIwtsPzvf3lzNbkTruvFY49q1Phm/HPJ2Uy1qcqfs7pRSMHdxiO+3v
vhGfJJ/dQPfOyH2CM+GbragFK2ixZhLZivs7j0FIN2cJHi5Jk+8ytdQqpvBU
K/a8bcLwnWeP3dHi1cXxzkUGyDJX9N2epb7pWCMM1U0hJ+jd9ECh2k9YvZOb
U6q2PkGU0eTYc2jFL62pWYXYsG0iw3vrDVVH8/bbEnEDmJX1feMKLzNPYmtg
ma0t2gk+Ongte9Su9d07zetOWGAggvetpa1scrGEEMzZ74YPmaHA5yE6bteX
T0YP3V88j1fFn24pOEJtaEIKuqgDVAzuQcRJYK9ZssnDkLd0NpVM1q99/nxJ
w/l5w7RdFmpI1OENCJr1rDS3zAriNghqRu6wBDDmlneGvux59B3EConce9S3
IbJOabES+/FMaKavR7FcqVnAKU8dbVf6NmQJIn+kU4tEk3FMO1Vo+q5Y//2b
unF4TAPutz2XDRz5AUt9//cVezP2xABljKFErkHm4qF2jF7Mw5JWQHtm/eU8
51E4d79AeaMubyB5mUc8gZk6PRCohe8WLtxDZZVpfeem5Th45vDvK7M3pzWN
OAhCFQiuzceCgFzD5FrmXXoc/EFZTmPSlAo0CVr/fb+5Ut2pWzfAD5yxzqQ8
+EjCPkd9FrzUc5MFFPMPeC7GKZ8HrpIXUn03To3Y/+lcvI8Ec0OsAjyblw2V
KMrYK6ofL+mep8qbUR5cBfoIUFO9Tf+qukZQW0+8TIe0RFNcMnXJKrhZvvHN
ve2LMaG+3jvJSrPoMiROTQcmdX1WCYrubc0UxJEiNpoVxT4wfTMU/nr09WDK
JTzaVphO3nCG1j9ooqsGyE9FRdZM/yDQ0eNHJDTL4cYlCfu2QYKf35/vdZ1d
2/70Yu7SksNCK2hA6PFeAU312uGqZmvlioRolo14o7bxA1Q++8LgJaBGk6Xq
xEPr+bKhe7rf6z92628r5n8t6wOECvMDRr43ohszX6gzFPcYx0EsohjSctEw
N1C7c8WZ+1o4GnfFDolomK9tl40f6JLxYjJ2W/jBmfa+YCshhV2/CsjU4mwS
epXkpqkMZxf1jcozCKs8h0r4YA98dzzFIbGCQufEIF7mOJc291mpYK9V1wxj
6YvdXJU3VeIwv7QTKzDgWxSmxQaG5LiXD5h0NCy+YuEu6Yx9ruKPHOQqnYrI
Ue1iZWNGON3ueXgV1QvX1QFcBQAQRsJCK3EtQNy29uSxyJgMX7VV7Ho3kXFU
8Cgj7e66nwpEw1iNVX68I23tCoPSwsA1FNYiewbSj8+NO3m46mykoOJRuS8G
lBv2yWckHm9KNkgHJ8I8VAwuPdkNxacJXIbhil12eCJSiVQZMRv10Y2nYDbU
/XdP/kcc7sBpqSBYqVkK5Vwo1zpS6IMk7fYua6OR3YIHBNEmYKOlM+6KfNw5
zVqhDI8f60UXkS+en9x+XtwVcoaEEpHIqq3Q1zf4pzODJI7m9pJyoD+r+Kxw
SHBfBM/7xyPoMJPNH6pIln7tfNFVoYRKLQhCJhhBgKWvz3pSH1sgE1rBhGio
uiSvZP8Zg/OFeTf+W4RHuLKKlca+Qn98jcW7tc/jpLPMVPe+rzazhuAl2Zfa
HaIqIXdgCj/iNYA2SOJLSuG293+ttoKPMfnMyzz6/D6v9REcb1jtRIKNWHuf
dhe3cziubkreopIDvePp3Aj3YW+9RBt5GSvx7L9kr3L6XdbbftVNHItsXLlM
F4+swof1VKd1EVq/qx/R62mR+nnn4y6rzwTmzU5EskXQwPnCaOXcqKbLSYtS
0SzulFHjfKQ2wr7vCDHPHP0+ZG3JnKU6FiXOnOGfUBMXXtbF7M04iIbj1XXc
4xgWIE08koE8JgCGzkKnBTjK4Tqjr/baL0t/EPcWYtEQe+ckOnjcIV4ghE6C
EIw+Tg1G5KZjVLhzp5K969ZK+LNGkb783EIc0UZwTwj+4V98kkasg4dvVTFl
QKPuYMRYTaYVetV0UjpTgum0LTcBN9VsZQAya3gyNvWM49PivH/QB1FZAfEO
OmLdBFN3Oet4rq/VP8d3WQoiTBl7xOxnMsgYoSsflkbmiaJpR1q6oaFIuW7W
ZZjvl3KsdZsPf8nsR854ZiET0T/0q+RUX6qW9fICFRNK9ggdfZO83CeOnNdZ
lEF1W/qN4I1AnlXQryf0OJFMnoA4XgyCDbgfDxkPUG9KLXl1DroDTmZxeC7N
+Kx7iNmwFp4rJ/Z6asHc6WIcMK3DV0kcwqSzKoCuhF4Ma8b/yCVlmNwP+3I/
4uOEoPVnkIGWDXFQGNuXTScVc89Lxc2KdrokFNcpzgc/cKtSHqDG1dinEKhP
qV/USgVdbu36J1AAw8rUBhgHu6wiYtzmeBDOA5JneraOU5bRsK1tLBWTDsIS
XI7YsU177SLy5d1W9aO2AUoH1COlAlOCbpuN0HDcv4bPa6cDqxGwAZQn2AnN
q1TuQMkWVCo9veihtxV8KoX2acEHBrXBapaBomUrgLIhniMZ0Juw1TZk8bWH
ZrWBi755ME1byg0/wWzx077PylwJJu29zMomaKzVwPz629bxQEs8XcvH1nqT
1SWymSx3yW7V4R17QhaePjnjLhqRb17B1n2Vw7b46UQ+ajRYcXw0Tg2mt2Zs
jXTWSHp0+xMZFFtcWbnYazuiDtGEBfTNX3hQxMvDf3OCmjSL5p97ho9MI1Z6
s/zTbgKl24fUVOZg6wepvM5MSspUfNEZxkKwv71gMfT+t89WxUz0tguLDcuw
F3Jba+WBP8cVlBmdIws6GoRVon5WAGbvizakPnAmqoewXK7LnwFi7vYXthCa
nu4/RMJQwrRCWABFG7fX1kxJaWOKbO8WDBl7b7/E/043NW6vjO1bpADjR23l
DRBGbychviRsi4iRQYglpfuy2Drdg7KHq89ufd2GYUY7A253/l02589iWq9V
6JW0g9ZcHkmQhjHOaPs1yg2DyvSTUH6fXT5KnHeDZUKwqylm0LNrao7GhsVK
/VL99D6j3GmNp/Vm6vmJHY0b9tC2cKi1LX+R1SUbA6RpL+9P3yK8fp40EZEj
mjKgwOtURSnanVN84TaF7Jo6ozMZetl4JCuFTkpmmD4VYOoXxxLsKfYsSZNr
RNu6jt//RGaYBaGKfN3vViHj3TI+YpUtqbezax/QMI+/30lq7igA8jXK+eEs
8k6E2wJHb0KRvELKN3GC/ADgXdrIXVnC8tGiKGQhN5gnj4dnApbJlR+eoKBR
zYiWekEMI2RDZsEforXn1G/YWi5KQEVm8Gn4LUwRUSfueGyQJH35PBx3SOaI
4BDBvxU734aJ0xk7vWH8NMBrLSXqnmGJoQmle2OjRcMFvaWYK1KtAOmGmjaN
4Wm6oyo5Fhm6Rkx3jUmVWcnO0Pm/235KhmzpwxoIf7wCXHE4pt/abinYco2S
YawfVreovZL+V3Tk7CMvn+WYOQJQrnLciZow1sMbzVOZwLHqzk90DHbCH1U+
6y6zH1grr8SL63LNKgzar/cGozrMft/wT9CaAgFfB0mMlpMAKQpov99wAMRo
ogQhaxAYvpmFqQj+wFp/CIo/vRoJZMtutBhsN/Wx4hIxIRgBsSm7iM/qfZx8
8PmyP2xiMMbxjwDU4wbsDoFjvRpNtCajFXvDBfQ+g4aXBd2i/Y2gtz0wtfFn
RYZHvfBah5fYTjs8rdiqYqu7nrmCJuBNlbR/xzsdsw7Od0FRkgwF4V4RjY1f
GCyJFXtjopz8men9NyZY/UNFwMOdSqaFmtRaTErXywsrQC7RX3/nYfvddSEA
puz8YrzYUxg2M45qgWcx298v0hxATX1KtBL/C6/3U/CZvNRuvhBlj5fwmab8
PXjdGTiJF/pD9Rzd5asktcs+SQFvm8bmj5e5IigkHrf3xZMgMmy7rvyjO0Hd
6SXor16CqKmoN/WH4Ys3zOTHBce/IareIYXRwnAdOb5rCux5EECzlS4Ve8OW
c3JwDQ7UCQ2rcxAPQ+qYMRqAwNjlI7sdbYr2x9my4G59xsLAG5Vd7jtGbEj0
oqL+dM9LgJKW4/N5pOIZd9aHotb68ySSsq+8sZR7rCldEjVP7y0othAJgKiN
kUEojRSNeAoJSETOtzVWpISkdT6uN2LHoUO6GlE2+xOfg+zzqtBb3CVIkROu
d+/jr34qsQrLeSAx7qPlmvvZ/VlUjG5cPuGgPHmMAWzRCjpcPygMcfEuWzu0
O3yzhwOYOyyAI932Bd37zaVU/EbLEQL0BGLaJmRREtbi1oL5N8Y62nGnJaA+
pRZuT9NCHaf+5EFEkuUjn6vDCjeipk+0/4b3L65xkdOVNIG1o9pTfdE+SpEO
jSq/ccnoB/isjCiHAFfyo9kBUgqh0Ik+nBm4337CUbwZc+G1hKPH/XYuJLMf
o3rAXJD/wmPlACVChLj0TaiALkELV+rXiUd3CY1I+LH9yPv90EuJZnXKshMZ
95NWdp99Z2rxEESgoQlTxp4JBKlLvvTjLKIfMOyHF5TQQPG4SYe/3CLoVcMZ
YiPU3e2QjkvcUqg3eph1FIoPoyk00n0qXU02F/KGc9j65q+4T3rJQAS0sMnN
zejSoRjBBazd6abmQNw35OK4q5MzlYYGDkLr6B6jBplWIJTbsqnIN1pB9ZzZ
DXWQEJdUHAI7XOzwd0+LbgJTCE8RMiYwWGNB34d95C/ZB5VjcUXgPhAY9QrR
pkgEof3NBL5IIf9oHcCL8zpZVuOQ/zO/ai5J2dmkMD6qfBlnIfHtvnKO6gK0
OTLhvPabmnOqNISH2aTuyKLtSIvXFNT81jP7diwLzcTyYm7rIZVAw8ldOtyQ
8e7I8c4uedYRwet35c4zmXb3UgBevLNUIonux6aMgeDSGIiwkruWGWNiweUV
1/1p9TL0HRTfoeiB4toDDmuaXSlV4zlS53Xql+Cz0yIdXx28oArfeaWIbxCb
NK8H+JU/6YJUggEiWw+1dEji8gYZOW864w9pYnW97kjQFI961VnxPE3EffhG
kJXh44TCdn5FbxhcgH7SNpHl5NTiceOTCaYXh/3DNxfHnG8soqP3ZUM9QD0I
IJKgA+x/VOf8Em8P6EMZ5GqRF9AeFubcDiLYEoYx5ch1j6S1HXjXV+ZQVXu9
BKpOnqxH4TQ94kmzDZzKS6qaXJvOEE/0fk4jXwaalvYwK98tfsAPAe03xdAq
rLhzFrQUjNYMuaVo0oK+En0rFiYJTQD+emWAZxvYflbjareJi+hEL5Y0jQdg
xu4dkiNeeNlCxKM0yrLzF3f3zMv9fZkORS5wRqVF/Kv+L3FyeVgTfO5EhI4O
DVefA1A/+grjwnVF1PnBVpzAW9fqfQQ5FQ7v3TL9ZDbYNR1VAx3o3HU3dn8w
fxTOGZzKp8Xx5OVxfwAM7777nkAIis+LxkI6YtdVBs9FgBz0PxengOBLN43G
21+pj4fayzb9U0/ts2/ATsurrbBD48Zyn6FvBe38pf/eguUQ5ZYTBFTv0CLr
FrU55CmsoHLFZBevjeepPpbX/VrXGt5g0nLzVkrvBp82JgJahxor1T10C48m
ipkuQG/MKmc60cLsPwgussM12F2kkTXnzsm7rZPu8qv7oEJzEjoH+6W26+SQ
8s8YOIpKD5MyqLzOdqVBvYPGfPcJ/DqOyWu96s9CdJoyZsynpfODhddPAT6a
yGm9YjxiZreoyB19Bed1RLUY8V/frTaG2EFnXb5PnjewmwbjBryuGd/Q9PBG
Vba+Ne+J9iorCbOlMvjIjtQsw0EABkh0vasvvxcZ9qYA9gbkwYV2ZYjeYfrx
FuuQoPmyud0F1eTb7NDwoZ5CuzJAfo4EkGvE3HrerpKA7VR7Zp9y52bP6GC8
o3N9EVs2/nD2lFNy4PUHb7MCFJANYbUdNoJS3PxFr0aOHDH2uPruu8/3nJi5
GuvHcTrzoRydF3fhM7D946aQZxGZyW8IEGx9NXLlryNtvm3XyjgutwN8+DpD
gj1AVeg3IX8HZ1FBDEmfiuMVqgdwhWIjIcXQn4W89g027WpTvWz/t78ckNvV
B1HD5hOV3yNusqTh2VqTGsDl814fMDNlReM/Z+cH7lAutADg5k09iBISSUmz
UMrp5J9VFQsJpW92dTiyULt8BKSxjko7Doxei7D0qGAJ4GkwU64NaULUcwj9
SielxXkvvQr1Ni6rAJTQYo/4ukJWnFAedOwV9fdcbcxxTJbLIyX6HGvbKE+j
cFyy9xz18XPCH2EJvOeWBbq9vjzIiRqUbWzhOLoS8qeZwo142qKVKhY5S9tn
7O5t1kOWVw4eLbk0RymDmgmUJ5ZzNBIs2fpOfKb2/2S/Q+USFqwZhSGKtPjw
9i5N1zpRUCj4vJRVQi6D0BJ0BaJlLmjSlcjQTD3szQZFnDvh+Uy+pe+ikIv5
UWsaV0Jqz/43j8rGlCLzFJG1HxYnhFCiqCELYitR9hOGFddHJL+lg/ZaWG/0
DW0SZqIFdkOA5Pmsp93lTzZk9UEyHv751mStbFB/IvBvKWFKTMl94DZe9phl
TzBSVFhNmYYUvKRRW9thwtvNW3U7ghYR4L2hrSS0adAGMYZHdiub3Sdd2xiL
ltRrUM3RPvqBAoT06fh7gZ9p5TxFxGcdtQ7oA9YGMSlbkq+tIX81cyIZzZDq
aC2FNj2TD56BxLwBio4nS8bQqv9I/diHbGMwMLOvdvhccRnFWhCCqY4kJM4+
ELPfv5PNp6n4oMpfpk1tmYUBt5e8ZXv+n9fxeW2G3ohM1AfMOK297YV+4EGH
ffqz5C/+eVnUVJynLkRtDa01nMVgnWMM/u0PWWFTrWH9nAhdtbcW+K3lp9Xf
BbTxShgGUYD4Y83ZFub0SLYvTzf3qzGnQTtgeQ3r4KqG5eVbxSVlhwmy/BS1
nvJ+7jU5wBpfb5WYoyBpwhmmbSBGifYkNCPrKF9RGVD4wDdMcirWyHRQvGs7
OXEXK/fH2THv0YQMj4b9IMhfh4oT6P2Sq6CKDkSJAteBzansR6S78f/k8Cc5
2+n4dDqUsSk7GvPpD6f6PP8beUz/4fVLdSsbpX4T5E1mg579kVdJCZUJHoS2
wPoxiO3m1lzT6riVo0obncjCz/SoxdN24hQlS8y+hyT77guO8Srs2s62GvXx
EfYxUumzUqIm+TJvGy5o/TDHvqlZMEthOzbpkOdjO1QqcVgrVRXeWQlW0jfU
qV4jTUMINBjOvChpDLq6m71lBtSRoyT7qcioIV4GSbzFrnVZ6JfvVQR8M++v
R2U47XV1MHAP8QwBD6GzGpK9nw1JRlZGf5BzkU0k3HpAqncOMW6CiXcrsFQP
xUi2PeUV+4Ct9Kfi+Mv4xnnNJuE+/5AhcUpI6I4UfYtejL3iNV+E9gVsPycc
MM/vkFbLTiUpupinXINYBLTDGs8n5IyxVzznDVfFRxuS94X3s7V90gbMwS8o
I9nFWAqq9uTC5mRwSHcl4WQLJr403PC/N7KhRweFAoZXBeuSEr3628YtESlX
PcaTjD5eJ/mk5QeziQg8JXv2F/3wNZAMzajrXti3ROLwPrT4lx8XfEMdR2L4
SwSNsopSgRCuVqwfh0J6VNWlfq0JB28SWrspt5vp8Ls9Vv6nNoZBzNOJB5gP
8KfeqQJzYsIo7AxFq+VMfdIcMq9vCIv1aXO2nDpSZ00VurMy63yd/150O50W
3OYggyOQzA4DbP3OGeAP+gvE9n5YPeNoaoGF37ipPI+Ynbb2X4JBrrf5EHAR
yhhHSZeSVJ8UwdI+XTpWkpolXv6bQkrUo9CId+JVwzBk6dq4AOmxQUtj3L3c
iGD0W0ztyLxG9DjSJt4bAm6ciA1CqcZjzxsrvZoKOI9Fj2UT4IRlVA1iWXwA
iHosK+BsjcdHuz4ofGF01bLkCjzsbL08vXlxe6TPvDRQUajASobM077qD20A
zH+J8zdITnOLwNaci8U7kvgy50sbbMaezP5gI51SOKGPQe4SqW5hUnkQEKii
HOfL0ovYjNxjdJkvQVJDdVH6SxJOC4OsxCdF+wJiSRpcr4XQVKbA9VYzLint
TJJ7QGnF07Hav926B6X+S0x3/uikKeYhGS0MfaBDJPOwx/yQkbuxu/1TMb//
gO7bgbtXzFOgX8jI/5H99FVpSqN7bTAtfWnflV45kYn7fYL/UK3pIqMC3Kan
v+l7Y9dIqofC522r+W2OjewuRtN3CSE+Nmh6tsDEPF79rswL9ZKmTwH/kl33
d7dhtmnQ1JP32Z5UOZRC7I2CiZAGFIHWvcXE3lJnn5uOBeve16o6BOu5HJgO
V+cb7wgLZaFfQ3vOGtZCqgk7KkUpgktbH4hu0GhQDiYTt17MYuF52r8wjdKD
DNDKr0Y24WXBk0LeLOGm5wBlH5a1J8PZoLvWH5kBT0ElQhkwtgcaLRQI4zYR
VLsSCYLYfsd4iJdSWSJ1m9vH1CDvsEhC3bP5mCf1RnNYTT121HqZZy8xoGn4
PDckx5beD0b4e3Jy2AwtlLCLf9d+eBNHTXZ+mpSyFoQbi393OWY9Y+kPjlnv
6v4SfNyQ5yNdObIwO0jXMb+ry0VQE2mMf+OHiHR/7cjII9n2DXHyU9SZxCC+
v4b6qDs+4GwU4LR73Ua/M1/O4ZFWdj7461HupzM/hu432Pndw+fnVnRHyIVk
We1B2WWUE6HTqp70NrB/8frXrYvq2yhde78QRrIlOjAdA/hEBD9ifwhqXMxF
pJNI9C0N60ww4H7Ivh2//TJHTcFB9ccsEDCrcy/V+WKuoVMoOULI1rSD3SUK
k8Ul69z4+2C2CGawvqo5XhUy1x4trifjeywjAuOmXQBpvSMrz/HL0E2NxKBr
xW33+ZDVSHnRrOIJML8qhG2FOqPtq9wGm1lu4GRIOaIqiSHeFOVg+lwkqH7x
cxowFyBHl4RWHPhFqbkZMG9kXHplFTRvENkFZjAQjPhiFKjIxToHx9N6Me/5
hTn7C8u+lsdWxT0QdjrqCco9IXffHm9Darl8a8VkXaGtwDY7yWzCWaOlQD/U
5yeg80RVp/E5o5n7q7tzLTJ1i6ydNQMzJ4q0WRj2i7iIXSIEfPL7NzEjPSKS
JfoRfap+MoMrQ7MMNUZ+o1417cVyXTZ0ztb80Z84gZ7YLu3uDok2jZRkzSji
wWVX9dbdGKIITkaFy/9fIkHSFuRGtooXmA6lWihMNOz3SAkfFT1E7WWItI7L
TubmqeAd0GpXYs4ZMPM2kQtD6aTjxYoHC8/1VVzxrsoYWiHBY0L11J3AgBWX
WabQZ13npFNBhNmespC47+vyZLyqjHrmq99irScrj2cW4KBFAaavB28Yfa7a
q7X2Mzg3Xl4ERS2fvrohfK8TkYjaMAiMoyZv7mUKwkp1CIqwZh0ptJGqtXtk
SVrD/t3QeZWME7qWJqk+K3YWlrwPMjWWtz2OX/mywMC748ody2kh1dfSn1FX
5FFSUiEv3HHxx/8a/N4lIQAJjbcetZHhD4SGDTDBsUCA2N45uAK4jt3t+Je/
0Ql6VvCQwUzAiLWg+Unad1CtrbNwVeFUAXeglXbB8NEFVNCjvo+vVDyHHs3a
SemmSHF/jDIQUj7wx7JG90HlZmirwJR9qpUfNnHxmcy49yhhz2XTrB5GJUWm
Rzn2WJdHL7ZHpt+qkg+cUgOx9/Yo4D8UJEhQ9NMumw3bIDWG6L3qnz96u+9f
VE7STYj7Y8jdjFhl5WGhoddtDTLP10yd2LG+BSeHMoYcBwtEjDWQ0NAv4T+x
GIB7GMkvQx8vgpSMNZFtGRFXRvH8dHA7T06ZbNsvusbSl/3RYoUN/Y6Bc7Sc
YLrrS8E5fMr0t+XdrezBfkkswFXkIaZKoN9wz4AGk505Gi6cY7ZRfKuhmJYs
lqrCxlJcHJJVuZJEcA30C2m1pmYGaB1n6tsBgQvAyLMBA4pDhEE2vQUBFkzo
9zDpLGPPyYMwvTYu82nWw8e6Ctdg8YSBKiBvDWLOy1KGklVQHKIURJdL7Z21
qTK1YNNya28TuSvFM+GNg1vKEn4vghI6qIWuz8bS3ykV8QzKhNUi73oL4Ati
GSTG5mtDV0IHo/xFPBZOBSPQzGOZ0+3PKg3I96e7z/GHE5R/TuV61mNGAjXo
8vRHFpS6gVa4PipxXv7EAQr/1ReAALSS4WPRN+j+VmxCTlxnVqsXqdinlB6n
MUAfQJJcDnTqtl53VV6jJze3B13B40mEKJrK3WTp/ShjXEzbDTgKpUWPq9a3
bKDoXURYZzehGJirEIfvfcK7dwCCgMDfpipiuEOtlCh+TcgMqilGANMA8IRW
BBhvlPAKFg3FU45Z90ezhJZIePR9uWcvtIIlvehhpd0MB4guuSfajieUn+BI
EQrOzx/+PtDIqIWqP/rmZZJcgcioHVq0F68z5GZZsn3RgpUxp4aXK/RTVcCn
CzoHkza4O2VuDiILHbAkarj2F6T9MuCtDspsYD8J4MJl/QWxgtgx6Rx1wqzv
jLE6zDJjLpraMV+GWOWjF5WVl+e0gFSHzSV8KXvOgT4WShRG9maZmj3JGHHr
jTqzx6DjQDqhoH5+/dVjuDF8rrsdTlbgX8Zb2v5fDhUblfehVPMMHzsi/sCY
bQJS6vOkfEgYTG4NX7rQDDOqKkulmvKfSWPt3SWz8Gf/9iPmgnY5soUBRvI3
1Dq+wMLuXWcBFd4cnaJ/1g9Lc5y1VGVid9PqxD2COCYy1ixM4v4i0gAPBQCw
zghfg3JO8TaE7DVNs0s51i+gokrqWv+voF38VBYRQHXa5/37iEw/e4WwAaLz
EghBxF9D/HN9Svt+5G2Ufg4TZQVhbTO0OiUluYgL6nk9jOnTvPFXbEtIx/nw
94wk1d/6MjKCnbYqfTxObOTZpAGGcBnXwQ4IrPP9vXR8G2IKi+3e/kLbGYHF
HGQSv9IMIutD75xgp95xGAfM9CqFdN7iEn+pMnH782jWpewm7D5OzdVi/Xcr
spSVMgtTF9FEvAHOA3ScegSfafExWyYiQ+U0qrKqLwq4oS38qyqYZfyVHtSv
FZ//spFU8alBx5VtgFfcHfuX68r5TALWiUH0DjDEJVsTaabfhGiQlzV8rgc1
+JkCqQ+pAjEWs4iesy7gOxi+/b5H0vxQhLU59eWw6Ak+CyIauwygcGBDDyDI
JsvsKKFZwhjpBtWxxVb7t0KVRHFPVER9R0KXpJ+T5M2PmjxvX2H44adw0YtS
PlP2BGjeT0xyeDC0vFi990MeKfG6mtY0eM7iTDbSkC5duVkem+t15k+vx0mh
zEsz0xAkCi5k7gvyZO55vbOVssu1CU1dnZdexGm0IvDHoCcZoczmY5fkAbua
DUdNkmHXmH+VAsD963AAtk8JYu35hxuiY9Pcubc9i3YjnxcIJ1/euuLIkRA4
GXRlc5msRT95GRSADYLChUOoGp2ff8sMOu0Tx3ExQ+7v7xIvRLBaqII+fDm/
nhPcBQH/P3CJNCHBMMPBmxlHGaG+f5QvGkl2m4ptEcirF5QzMkPqF9mhHbMz
OQA6BWfVyky0TLu60crQv2WiYJ4QuzzDXS+CUWQKB8k4zMy49AJqVW8H82xq
FyO00nD81pwIFfmecG1OKgQbsINEblvQPpK5i9uRSw/KTneFdnWnH6YPFZQD
SRNZmhNTMVlTAzIcvzTEMJI2MR6NmKiT3HMy5yqrBJT29+9RJWzCQ+e4TP15
/mGoTij54tw27zM1ZlybGz43ozgbxFHR2buDEdp7skUdh9PLB38rSKa2zl5p
QCTkIvUvfvTYXnzALTbfGctd5bXK/QffuHE5rWtjiW9vKXeNUG44TzcDDBBW
ZpBSv1tDI1lyNYiLgxqJ+7SRj8dhkTSzkW+V8Vx7H3F5z/mb2SpChbFQlwAY
eVs9qMZ0/wzyfZJMM/OifK+Q9np5ulNFGfPz4nH+Y6czLlTyFA+NYtwU0532
EBw5MwCQSZhFvPCHTyePzKFmsJjeHLRuPGxaah9cHcFGRb+WHx599Bs6DFR3
6xLSUu0hJOgFwqwatwUnFfHo7i0dn7SPjqIkxsC9XXe1frkdLnLMBaX2FE13
O97RcRUlBAIwYCPxKGCG9+nFu0LrlUKwScwz+AQWtFqE7Bqu7W20mfXgxG6X
Y5MjsmzzVATsGEN2whcgSRuKNdFawdhv/86VGFyR3uWHS3yfuFGJq2DDFYX6
+Bn0RoOuh1EiDUHcCBrfU7Emu6/wFNh5i61DnDFDFwqzoybvn6JEUi3/FcV1
yplzp35tXOoYeKfjjEJzydlsGCmyywDLDyxJTjE/C4wp5SEKZC9W31qscHCk
nntKUixDs+NDdPkeQXf3jm8pwCHvn4HndOgWf2b5g78s3oaHkGIev/bPKATu
j9wCGELIdOUncMQbMbWhaGnw58nP0g6ZFhLou3MtIY71BRgmKs5TXW4mKMr3
/eUdxuYiCBtr7w4YR1DZiJgIjAEFMwBq3d8wii1wEWcbXlM/1590KD9pujPy
4SVRBxVBNC0MX41k/J/cpVu7z7m1saOl13VjF3vcVOle+fJFTNdGNfcBApQ5
DpkizYn8dSUeQNpPDL1Kf8HJs+ckwAlXV2v4F09N5WfnrOJ9+hOZgjo/3BNg
5vslrTRzd3Z9ggsbtZGniJqsqB7FEwCunNSCrVv6f65PUj5zK4g5ktaQQ7EU
U3S/tJQv0RwVzc+cp3jzTNk5UafPQDPs54EMlBrVxAo7MEJ8Zur5083pZ1h+
vY+ZZ94cYH9RP0ELp+9kMfkY5EcvROlMq0Z2BC8orKchIdTtwawNHifeh/fH
qDR5hXnOVHUjjWQhLw6Fdc9h6dYmM0jvsX3FYopocDkDzHwpWWo/ytTHwQDT
mrQJUgqx51WPyVcLHQVVA7vsd1IsjW7KAYHoGqcJhFBlr6VaTWjiX6dXJ3nK
fr+ZdXtULN9JHv1ge9c0gBBjrsgewRn7GRd5O156edRJygbAVQX/zWW2lHG4
FCm+1+1O4OsbAP+nu5CobH4YVMYxxKUobxtRWM0RhP2gfd/z99ZEsCYQ+nr/
W1SFdbP7CmaGo2vtC73fzr595ruy0+oQXV3iS6mBIFrOJvJ/ihhX/wY18KyH
4dTLKeM703YjWJbQUhptwcU+AkNBSHLJJtBdcqO5UgQyrFbl1xj4tE+y3ngG
PUQ8AyySaGTMBB0FzdnozA8O5J7IpwuNveEpQOfEEY/BuU6d5UAZ6x6JzyFL
1IZr8TegPxysylsyW2bojcE45zIYc0EjMw/MSDTJ1RB5u0EhUbkyML7yibKW
vg81eky9/k59fkyB+/1BDMRvL9aD2MV4+gMYZymglVvs2CGIl4a+Fbdr7aES
lj5iRcjHXOEBuJGUDMxyf/4ZDSt90zL1WkvA3zFEhY7uu3r2Je6dnkwmXKc2
kb50QaBoHfYRpsVaRWExqutO5+SJTY8TdGEbSDsoNOfSAjqUwv4HIzg36xh3
G9ax73YYF+Zhsa/3D3nxmYLs4Ir53JvyZG0R9TkY6NqODT7S8+5wVJNBmkY6
agHJPR2270IqgP27yiopi5zSHBx7vW86KEgqK3lRs+mKgt5bcK0oeQjkjPPz
+3NAneZRwXs4f8RhcAjKmwGNV3Dhk2QEag/snKjRVfDaIm6SSzOabZvjJDrO
DbvSRUSOL+0FPfajdL9pPQz2ogA0HhaCa0yCXqaEepwxs+vyfatZTqaZc9Ea
mejqI7KzqZpQ6sCOU4KBlnDqUf+vh29Opo7MPqN89NHX7+gozozndIK6mFjR
svS/I3toVsQ9hyYoFiW2uFScrL/uYxNVHyLy/QVfQgTIj054+j3xmiCRnsQe
IpNTO17Kg1VLQvGXYTmNlSPdTYBm1M6cgHqDJnc1777s1ORgeFBtdMq9aCqP
a1f+MIt17xsX20GOEIO04kX5lZRwbDIyBhUM52hftAF/c1ROSBTHZaynslIs
7zc6yAz+je1tobEnZRSL98JRzK7Ad89CpecTFm2FWWJvt1mIZlUFub3eBYqx
BBEYtRdPFiB4BjUSxHKaDPF1R4qSrh9AtyAPkcMApxQsRmm8DlqvSk2X1Qbx
/Iygzv1xtWeeEwuPwaPSnkEfqdbTUW73llWIU+r9joO2ra4NUKiokru/Vxkf
pfFPE7yJeRiRA5WumjigRzjonObspPvIDP66ZkX3aJXv5dmdjPSEpjBsCz2L
AE5uefXbLNDfG8ZdKK3oMEvYGDjVSHOS3Zf9aWcPKvzStht5odD8ZwmG0L6P
7scjUjKXTO2Y58Y6xRupFQbl7luADtHtDR8uLW2LshL2FM/exb3wbidmEnmW
Sio+xg0ETSCzu+vCZeNdAkP2Q8qqaOW1SHtWOjAT1y6++v1S/4W5gp4v0FQC
ApyLUUzkffHxUXsImGxXMBW5SaBYd3FqFGr6kBeWpiwObCfzsuwTaLMcNOJO
MzaWqKLefvbiyJoayzjvQJ3ow+LTlyAdbP7xNeQjPKZrp0YiN+FnaLXL+XY4
S1zUNvgVky/sOhdjdbpKpi1OYa0ZjMVFIKNxK1y39gms/4PAExKuz1ZFHkAd
2roJ6v7z8kRBeJRoC5H1LlPNWS3xyzmRPSZTSrnUBhN0Ylelazf8TwSeIKRJ
3a14BLAV/PArTajYIzOK8S1C2ISXSRZdjgTlmTv5cTek7auAlwd1d5dkjhjD
feMMJqBa8iSOjft9wypyRhHhMGTPASyHDYACUXgtJUREEKWbHG5V8FphRTZ9
BhbMTxJ9GfbmXl5fMxZvKqX0CF8ltBCjB9qsUhoAsNw1zeLCKEgqWiy6NJCk
/eI8kFDDAko0I6K8KYnPGf2z2eruGzQ+MbeZCaTHO9bZrDwvInxztZeIGUeE
4yQBRlMfHxKul4SFHoVYCpABrHaINpvjWHI89BDXeSEfp3FuNud4YMA4SZeu
pZoEpauHh51r6ukRZg+VoY8U4pgyHw5Ua62NhG+RSI2bHaf8RvsLRBTKi4Fl
3/Drj4936Jv5Q8aRXcP1l4zEL6m9B2IWPmTpvjRWOx/ItH7UOldP4sekyppP
dz8+5w2gYjiWi+EVOVFP2SApMwH4Ms/2iHjHWRk0vanj7Ur4VitIQzq2K9yx
eySgUWp7bEd97z49eGCobIfied9HX7ntoKuxgchmLgIT/BhUu2KWAxA6r5dx
MtzBvMtApk7nt4/qOQYi8PDf80sL1KBLV3dJegSk5b2ZC/cyNyMeykXJOsd9
tST7Qqbj3T/I5SZC3mlMLY3hOvOyBlyZPa/W5P54rL2WwulefsCMc/uI/CoI
ZkdfvrEZTgB/sMlFajfeIhOCaxBbU+Q2PQjYPAHTgXV1DZwXquSx+HQaLRCT
meGkcfckvFInXo0f+evMvmF9sET8gTlg4G9tnBFkoORdSFo4NeHxpmpjdQ+Z
gYlt803oB7pj6eM373/UfB4MmemBi0yPMIszgWbOzh2DaoVz7I7923S7xZSb
GayF9TgnKkvCyAIAICJXPBL+AGBp1Kpa+72n5jJIQZFSCqQwNDLh4DmEo1Dh
C4K9+SvXK11umlQKGyp2gPMRHqHZ4utwZQg8r2OhHMxXFbRPk9ZbgdNkOqXv
LpNm6OE+TJy4IDhQcfK4tD1MZya+1qKgAnUIN5o5Yh3d4bYKETmWNRpnMyp6
UpPHRSDr5dOcrgiZ1Yx0PJ7czr3VQrUDWWQG5lKyGn294eVEwsvMtyaQrway
XANxq3ioukUapJLFweWFZzWCfKjHTtSBmReHHOnlkhyEb5ZoYK6j5xkrtnJZ
2nWygCq6t+dy9+TYui31HTRf4bl7I01iv8QnOwSSU9Efb25VdmrkRKaIyhSD
MrZr332V3A4tI9y1BdOsXHXE37+n9U4euPSZeMiXhA4miknIH0To+XpezBzx
Di9JFQMEurmuXM+e9UlXc2lKGY9nnobkcmbjte+Ra7ihY8LBGvJhWP89YwPA
RH4CrjM+mRJdl8rzDy8EyBOppl38VLxVpD1HvC+XQswmTcfN+YFyDTv3tl9c
sztaRbnVRsmbcKO4s1fjR0SMLmwXlT2CWZ49fOl+aPveHUjN2BDh69M74PVT
saoLYmWRUWulxe9jvd+C1YzwvfvFpjpRf/LrPcTC/ZmmcX6q+xyV/Gb8bFL1
EM1jB8qv5WJMxcgt/9sbR/bdJNCVZTeQhzaq/XiqSq2O/+EAjGhLVcJG3q13
v4+XqTRpl6odHrI7acIcXF9pwahTysu4jIv49x/92vP33MSDk6y8cngjATkJ
od2jVMW3IC/l6g7o+rrfhQ44ga5tGMrA6wsgupCvvzZwGBcpgLWZIyScPSgy
QdtjoZoJU+84ptZKf/RrLqCbh9L2bGbEKopnyVPzcnd/M2MefcfWBs3M6H6m
H8d4e+39Ekvmb47jTJJjWPBEjcHay1J1tSnI9xDeh+Oywsyi+cQvJ28OxZn3
J8wQBjggQonBGF7m6rIINDLx2HxpkmlAtTNN36X4e4GO594BvW9PZ25EN+VM
5GQlGcWQWe1RxhCyZ26qWr3pw/0J1z9Vwt37WZnJEn2z6wv2EKL6GE/nXFA8
yOWp5tzbQaUERivjLhWFQZ/hE8pL3mOdjLy8nAe8GeJYWKzvPDDUEdPwKylT
WtBWnIuRoSFhKrrlA4rJG5Bqjoaqtfte+RwH44/+6CieiENkQnNKfOTBg9aU
rAkvS/pMdJgPKbuvba5j1sVGCSoy6Ggidx7GfbGWLRyja8hbf5zpOf+DUPaX
04yW+b2TgjWV0UvOq11rZK1vEeVCyCqH88GAfJ0FaEKgCRBEdcl+M7gx/Ye5
0cs3HGd0bfRPAVLULmWsKoqXn7Urf48Fz3jA6FpXIGhGMcr80lGqM+g/Loj3
Tr2hbXTJOzq6sJezM0nFLEYHVLarUYrFGtcgejEeNXSDGuS8fy6PQCgfevGw
QaLzqpULtFIF5uTct6I31vIol/7+g/1Pba3tIkExl1KqMJwB1LM/qvxqTDHi
qA7Du53pyXm349y6GHVeAbErZiAGW4kudNY7vO0ONVS3C8sYGVn9JbGZHdNq
7ctQx8hzbpT4euh2ppypVNnT+TjdtxI7vzAH2rvSChmGwRIpzY/mkkChMo38
v8RLLe0sqE+ReJxb+uQ3QTJBBewsQCzz5enNRGYKF0h6/fZF7QbWJ+z6MQBp
IFMFO+a9mMkAuuB8c3aJ/Ou2sCWImjNJ3AyyBQms/JBf9ZPk4PgTN52P0AoB
m85MRVh3m22wRjyHXOECV3BWl14ftllHwdPQNXvSpmSGO3ds0emcyJshnarH
FBuvD8CcyiLeP8+Dy75mjydfq4m85kQasjAWrcBt76V0WewHl05v20QabR1X
73dNYsBff7TaFoH4/npkGIpNGj6pAy8Qh7vlnovQ8IshDfxnxI0aJf4k5C2i
WX9ATUSETyqtZ/F8Ld/6XoWugVoN+bSUSI0/pdosFb5EZC8y/lVeaUuUaror
W622bnCYEMUtKOpjuayQFCznRuF8QUU/s2Wvuy/m6/uFiTvMknfe/LLP8TaA
Fph9eYQO7aSyBkibiLFwMT3XxZQrbw3jVTt42wq/nIhTxXBxObnNku7Z5oo1
WMuMONPDDRKUTlmWqQbFpuMWKk6QyGhG+MhDfZt5nka0GLQtRdPfS4ZBRnxb
ncWuvbBJ2gyfUitxb69V0ZGMQla6mWRCfdcyhXWlAc+REoiF+OZGBY/efcKD
Csy6R+8BxKhTPI4GEaRiIcnrmapfryEg3t3PAnFj1E9iNoexLwyAm5QLyoCT
MK/pAlKiHk1qmC81VpC6sxtX/QfleMFzhoTY3a4ESkwn6Zwv5p9tSnV611YV
+5q8tcXWRfG6dyOTQhszI5UnZgdJfDinL/R2gNPPIwHOuy0xg8jpwPOGCYmi
ZdxBsA3huglEQtTJHrCuTnFjkJPlDNfPlFLyAI0W068o8WDsJzODchyGFU1S
pYh1gligNylDiQozxnPNQLbHompwvLlh6e6A+bYbqqSqV29mVUPTeeuHq/Wf
MYzNflqKaSZKBrYO1EYpA+cpEGiIiWuIRiGs8PQJ0bLuNFmaYcmst3rAPq4k
hYlrN/ug9xD9m7uvc9ukJaHMW17+pIyWjJFaMlmcqhk1vChqJdOMzh6ds/ZA
M6NnefFqPgTBXkbgGVfbh8LS+iQHFP4eW8LXmRE6KYYEEca7FWvSqJkpjHeH
qJDoZ9aT9byHJTrQuMKKmDgucXMrHxmHMzxbwy0U64va7Dq1xfB/3JN+6XFQ
dLtr1gBUQHDK8fzeN7HhkUrQLJ2KgUx4fnQzlVXPKksqPv92uihVAxE2cxEt
JAzohKyvyjBSpfd2i3rFS1fj5xK7T8hDsOSZeLdBBVgd3E+ZrkwM5OQMDVp3
ZEhHpmZnIBK4SEeY9vD58sNIaMwbo89PR+9e7siiSuvoQD+VuhX7tzEDcI42
JbgHglEKyirIDsczL6WTvkEB/mvYb5ZDCaeacdm+WEKLF9v576DLzlEcaRFW
kRhxvMY2dZMKUkueuBSZyAhjiY22R8M6dBXxBsz79ME4DOM7GPgUrMVtOpcr
ig4KYFODC2a3AJJly+SkugNk98VFtnYPHxApphwBxKFW0Ora1QOwbU9/Co1R
f6L/jOVOdTJte3UrxmIQv0KbYOxuPaHhCfzl+F8ufIhR1Gig3U1BWbT+k126
4CT7QV/twiR+vbAOaQDYOfvVoFdGrOGkr1FyhMkd2P8/GiBU4UX30vg0AFRD
sP49r7H9+tv03h6rTc82xJe0rOwryYsRCq8nBKKRlsM+MqW2YDUDu+llXLwY
DUIbHSXl89ts1M1GFMr8tI/9zQ+M7SthLTW20PJfOfLCSeFKQfaOptN3bsMu
Nhr1//pQ532+zShlNOoEbcScXq571Fk8nBx4YKgzNWRTdpLvnMo96eTcClmE
ACE60I+bUGBCf+cCfSxDAn/B752WWcUNRDOiX7GEt+bEgabMDBZyJIi+yT++
OB6G5dARXqIl4cOLAc8ngxY/41GQDMSrvMHBL6SRaniZzqYunq1YqJ8QMPkw
cav2rFOpLs8y9Ia3mYzGa9fzAGYXjL90hoCUGhVlPgf+1bi/HfXtYy9poHii
W/5Y3rftRhoz9BE8ILXBnaVnQlnZEfwztJRE6YjOa7hPeBwNuApozSqiPpG+
hl1cip9W/0sZ3e+oCjbIW0+3LE8IvkdWhuLLrZ/oEHVxmqM7vX1vXMppLdiI
ZOae1j2Q+4zsgyoup3E9Xgvx9wn2Aa3wp7OSURSv9mzhulLel9VgHt8XHpC/
TqNam/T/IduxAJBA0fk9xaafw0h3ILmR+lX7wTRQLI+cZwg2Cr13pFL/fiM6
epjgTt/jeFvuRddrFLxSlrEq1f4dMPQYz6wd+TfjVnRcbF8+k9g+WFvY0Njv
LQlFXNwkSgrfmSc0N4gqv3IQ0TonPxaINT/vvAgzeZBovAlWUDo5Bc+kHyWW
MJN4eQiLOPFajIVr0VUzJXKEB6HCW+Q5vftxdGMwgPhzfwME++P7oqj5dmqc
g64ogp+c1uS9QqEQL7hgN80EADF5W/yxcJI0gwvlHuZtIcA6sW541C96oPMf
ZDtngQOKawIMFkJLP//2n6zUVMTbNuB2gYByBtENbZ6eSXDT1tji4ZKvndtG
FAvuoUE10oE12CgiT3NQOGLzxd38Qhn8pnX+9P1aeQvrBwtA9suqKn1WNtTk
fVoBMgM79ob+JtpVj/zf7wVKXyTGsdeYj0fOWtK+hWtpMoF6jmgEqZBYirWJ
UuUA4Vk4yEFsCL2nI4ucF9IiVu3kCr0w9T9KfpVkjULEgN0pHiLdkWYfpna7
1bGRhVRyn+Hl/sZbMnOeoaV7w0hCrKwFgcJFxVO7JbJfPzgW4czl+ckjYzJx
swqQ1XMFYGhX3CAhp6ShzvO/yKk4C8+9V0sBU4Ki4kCLobbEJarUU0BImc2x
hu+Rj4ZiSx713po0fiYt9zzey1marBZLqx+yb0sAucj2YXkmRci4DiSNKPS/
DgvOdo1dsO+6JKAvFvDiThMmVt1xiC1rvTkXCrBEzKtuCSU9Zocf6E2N/8k1
lcJPelsiSio6z+gMvGPCCs4e+v9GOH4EJ9rgE1NjC4TDi3Z/0mf+aND8o8wu
bnyfFW4k2YgtQi3eEE9rYfk0k9qhhtN7eSQVrouagBuYrB9o8j79TVFkmlgo
6gA8wJGxxByJ9o5ecnj0qZGC1UruxNgzMlRcV173sSpXPNmZT5zC8XfTd3GD
k0EHJhZqDHtUx6gwIMg+1m/UyD4TigzfYhmPyIdprdxnhrzxhJMFP9WcLRt9
6OYRYAOJdvn8+gVe3gHnpCCMtmwX2o+Rd3vGO7/SfEbtH7v/8lQVYhccLJmX
SOkU64kxWbcPd+p5wFqJoF4wYL+StbB/4XWW0TLey+YoFVs0G/NvDTyisCYj
vLZ4hMQvDriQuHFeUpwaZeveHjyqM1TBpA7r2R05hc9wrqVIPKwFVEertN59
SIGTx8ygh3M/5JAtKOqUu94m3Si+cZ8W/Ty5rxu23zAoaPGwNwMVoTyAKM3W
rRynXkQx9Q8CMUhwrb93aD9oa4oYbiIngaS0RXREqfTxl4ZYsX1jL/Doo/n/
YhUK6EDBmguUMKsO1MopcnYLiFEeeCxFse9HyCExf9US6XRbg69v41w7p3aw
qqnRvC3TvWq+a+qmSO0IF0AVFxxNXsi12SxlBbUrAkmf1AzhBiM3sdAiCWJo
dzfcGLgseJ4MQuzi+Qqp96Od6mM5u/jwsxHMqwTXzsOv3AsFAPXGo5h2kfbx
kEWm6Mcx+NouKa7Nuu6Tpe9nyC4jCCK7Llj7j5VtMQEb3jaficdtpD800Vqh
m0tnToROmkf8y0JWqew9RdFl87Q6Db8JW/JflaaHlhVeB6l+y+MRnxgyxdSl
6CeoYvdR9HUWMwCh5HiATUbvX5s8tFm2CM/kAB9WDz5EiuafqmrrJRxlCMyt
8p4SNgQKPT95xth6oJ8Qqb7yDV3xNb/hevMNrzAzRgmnXBw1SAH4O99Qa21B
ZvwYHQ0n8SkSboBKGsAcxEzAynteud9cIcKT/WX6JmdVLMTxH34LaWr1iAD5
hfH1tkQwFQc+P2bYgCLSo9O/siZRJi2jGX8aWgNDDwbF47Lhs+z7lGnhVcFp
ZpMnMhHub6Na3kcZh5LdA27TctGYwgdzQjNV3SZzwAlJpG51VTOfjB6NounA
KH6bsms1TY6x0heiI2hhz7IfLp6H8J6mK6YEAFGCOcrWwcWHNm0U1/LZCx7n
RDmA4DBULMa8rSjghDTYcDcS03Z2V4xublTn14LkolUY5xUMeYzow/qlsG7i
YsqYCJDjo4mhHB6LDzWNpJEHxhFqloWjcIMo1ZQNTSBlk/kg10PT/7buDZFR
jSrMjpGiwQozYYE7PJm4NNKdYJfRc86sWKcGE3GD6bBGjnlVEKbu/Z88nsOv
fEyB3twrWzX/IfLa3sWZ3vpzIKTd8ftSjLcCDnkHbCXwbIEcpc+ZbjwMC2ny
txhJMZUtvaNJTUtspnzt2i78Z4kXro8bXvVePdm5HsrxZ/5cX1RCAardZE8Z
U8kkNR++/8wXhil6Wtj6KgeyQJmv7fh1R50MvnwkQDccbPIwoEIaLzX7nyrL
SfFL3yz1P8HHhIo3aR84KLHEwuZhTX5bDCGAIgq37MgexpSlL9tKPyRLUSqW
MGiS4qUZL1epSagDuixCyjWPaO4tfn2Suja8n24RL2VuvUy2cGiDwVxbWEh3
MGJpPAk9Q3VsHgNaI2XMfHJqaQuVkVmEDD/gRhDse4YcKazBMeYM5R4omawC
xgYtPWRHI8Dim20a9JR7a+awyVQ4t1QD+9C5nU+aCheQqkOQJFGFU5d5irzA
e/XdxmlFIHFkoxfSxmTMLD+YBweI33KdC72S1/AMhHch72W2YEvZlSL/Ochc
I/tx9Jrimwda+wrY9y9lfp/+gDBULaVZhen+lhYwMLKwBRqKi1IdMstiDJBa
Xeay1WAmNHNOPkj9asTlglUzGE28NXq516WC3ne8XBPwT2u77s5f7t0t8aRt
KrOh0p8rUj3/ALal+KXMq+j94AboBCVAPZ8+UO9p2VFBcZklwfIg2CldYiQa
fdKfR/PJ+OUcplUoa/mYScp88sywl4WbY11/JpTExX+iSnXDd/3E2k9NAhv4
QcGgb6F3Z7e6L9Up2yHfZdVLO4aVBqUX+LUAw14XYqi1N134/3uUTfud6zQB
29JpvWkOal+cV7Ix3Jm6j1p9xTszqj38N9tuqNkbqSwApaXEAs2SAQViXbrE
J/7WbSRrj4EeZby3LUZ5vMq+0O8HLCUqKhQ3eYxnGPS/rSClNeWRuVfpZTqf
3GHG3R8nMMoKnhvnD0NH7MNF1yGdE6ejTeS3VEdhjiyDPs75jaJFo6sy94X2
qVfwYJSKT5I04uuvg9p7WOCO1syuogDWGulUGzPJ6Vwsd4w5ZQDd4ADML0dl
+4kdBACj1x0SA/WP4PELcKeX5t7Hv4ibxkXhkNPI7Unpe93NDhgKrqj5GGUo
uL+GpcZH2XZML5EYmZymwm01sLyPI7PJ+M9OH6uj9BVYP3ZyZH0+7hWO0Af6
zk8P4lJkLAMOy9sauGTi4tovGBTIEA+Vc5pDk/jABbZrw/t44EDPr7NvfLgN
XtfAgj22ujgZ61MUdlFZyqok5i6wFcnBmQOFRtshbPgluyK5MJyksqvMp1QP
909O2/XlpVA9mEry4PXNUAu1qrIS4Hdpb2DctPbTRumoTSmB5FTpOyKyJOTc
BI3ikUiuSrk8JvwDc07JK0zgSqYzTmghryOfuU6Wpetb7emkDqYRSN/fO5RK
9fcY3cKwRKcQPP3v0k+BFaI/VR1LKDtOzCzrrYInypl3fZpOzY0yNHk0n5a+
FSclODPkW0NQhN1hOzXDbWaoYxMSmxKcwzuGiyKmbyLtWfm6TJyJh9X5ZbUo
MLjtjEiElAji5kXJo72oHv+XJlspgdREm5d5xWDEdPWoghO3ISL3cuIQ+Ety
9u1LHHwpv9WLes5RcyaqJMfjlW9OAb6ALex7L3OCrsiFUhjA2u7Jfo4iRU1/
qf4zvSEETmC4hf6h/sNh/Xt0GZQMJe1QyFQYdtlIvajFkpGXYfw9T5VYyRpC
J2gqE2oc/Hy/oCdvTYt8Pa7SxVj/GCsR9EyFExX53ym1SIV3Vjhx39fbVF1M
F7yDLVkGEjC5E5HdTgLBrQWmn+1TOk89ezk9rATxczRjAVwo4clXyjktJeQh
RLoR/ewBoHbY9QizPwhUASioBaEisMIfAQwcRs5Kr08lt7PFB6/nxkSP9s+q
SEqLBJcRwFN8wRtUSDnKj4Vry+/n6lCB9tCx8yhSclGE7LyHS2zVVoKBPxSo
efh+RnKkEYLYsqofDtaw6+l9mMCEMbQGFc1xXaOL82Eutp37Toj9A0P4hyl+
b6Q/v29s5bHEjYocRv2FeJRdttBf0c9ifO+Fxym6BLN+H/rYUyWmqR1Ea3pK
/dxUMo1/+cuWTb3f9Hz8SY8iiZYsGbGfEz50cEnK7wP5wB+SbXcPVFz8xEru
yPBqVvwtQSfzH2xJ2ycMR2DCXbjISiv97y9fS53Rlasfg0KS6i3k3ObVbubp
Vh/7cmpiOahR3XMDePClwn1dBZbLVrwpqBorC31VEXSbITv6RAnlp6JJxzLc
GUzGRmDpUmJS19Q+Ol6NycyUzHMJvFJa9vH/+QQRunTSdG/GjBeCCBX975An
f64wiaT3WFabmnF1PfAiZm6fbROH5EsrNUOdiZi3rcak0vXAPbkorHCFirpE
X01e1K8AO1UbYOOo+xgs1ecArkbnRTQ7v3g+WgNapajFYUnaWi2+J5JQdecQ
StUIerjg3MrAR7TN5cJy6Kkdp7qkda2xz3UlsZfjd0TeL0AIrnApnUmShAyq
CBkPrKTXXanF+BWtMbadXbG4HKkN3I510lAFgcjmqQBhFQnUfpmYwA9FwcUT
fmJSVu1//irx7B9G+fUMdResu266E26+GUVY5Qojgd+ILbf7Xj68hrDWI1M9
I6Ect3wVn3b0zTGbfO17IHi+zW4L6DFFJLlj0Tzfjwx5+llYwWGjr+OdwQH3
zkTen6KZZpCKUE/al913Qdc2gUratvHNfbfmqEfiDzG+E184wctfVV+cS+Rn
N1ZiDQz0AasNaMwnVShCBOe5ugrWF8+a3cA+mqs0ZJkutP0yeUF5my64KJwv
uJvT3JHgX/d4bE+/EZV0tpLBBjJRHxeAxYPeCMbnUqNTyEIaFCYqjI5Y0C84
y0djTOa1YMHfn0L6OUfxFM22MZckKJHmaYLR76DY36naA+XlpACBiSOpHsru
3NbkhP9M3elQiQOUvKex1eMwrfcR7LcZJVYhrIbqGIu9YRllWNBeFL9qVhQD
gVwJDOT8aLBrBBu1XF27w/qvzSjxC7Zox50XPdp7aKC6RdTTcdEALQtbZj8k
A9HvhUv6n9TbSG7o04dshBFcRUjuQ4GTsxUYN3q/ZEELDzI91sIhw2cQWXPi
bVhlqoNUUWwvyxQaUDHFf4zZESEwa9Bmp7Mf1kh5kQ3aMo0GNIn9yqtLflaN
t4nP56FA2GzEcNpQEmhjW5/2jmMcCGR/DEC7iwGNPkWARKCNwgIn1gWg7ES4
RZeH/mns6XBfz9/tJseZH7G/HXd7rw8wgProBjHNfqYmhtfdRt9BCL9/0ksS
SOS3PSgP/nAfGavWtNW4vXR+TyqWupf6nBPgqLByF7GCvk7z8JOKMDW/pKXm
em5/3xel7BTh8ICGTEnPmumEJBqsRBvUhr0NsOrYFF8CinKuhe+KZ5wO5449
Wu/q0Yk3mEUMZNg1K8NYOvkQKvedG1f3idJEEGujtMDWA/qyQQvAM/MmApWw
AACv4SPkpvAEMI/56gROPd6klaRwFTJs5CEeysPoUKveyJQ+3may5fmbKNh0
gvfDsAPe6ewaVpQubZ65bPl+1J3z1/uoVv6KQuPZqopJ53U/h/oOQYd2qS6Z
f72d2DfalgdCuGjzul4PALwJdGXQxtUnWkfPApQPhKRR3g3B2d8Pc1v6NTPN
EJB1Jp1G4h0sjAauYTlwZw57MwHIrM+AB9ljYKgQ7nWEwrcAG8IMrLhrhrsp
6kQ1vzyXX0ohhP1Ivd918b6n7AUmJmaEHW7geQASUs6DsqfVDaQgisVqAp4B
p6AAP/78Ih7rIMrUks5s4qb/J+28EFjchEu8ouCr0zPGzy8XISqDHgNqzhY0
wgFHrl9vQUUG69qElDbBwn5XKjSuQt+9Xd1R7CyLwL8dLylAo7iMbZI02JJL
vxSyWwqKHNRJpc6BbDqDc6GzUq7rJ0gdzv49IJvNIkoUjpZOjFDyT4qxmsds
sa3a8fOEeDIgW88jvN2R+zqR6zXAO2anVswfe8f7cT3ahXl9tIJqAJBAWk5f
5TZKkJ/7zdxNIHK1Xc3Jx57ADP6pUSrmPEhVlKOBMORKtmJWP+hqtOFGlQQk
4niseZD+lmXGxD34jd+WVTnmAGLEHVCVfq+j4v00XV/cd3xL3tk0km5roLYp
uhsl/c/8nsDS0AMcpTgX3ClY3U5FmmlSS7iFeYLRcKjLG7f/48v09OfVFQ1U
VcObLnlvNz+3XH6zlruJdiIiC6oHM+ykUcCg16UFHPEC7NeLGaG85qzAzSj1
0jKhwAqu1smHs2NjRYDF17AcydcUc0SJzLcjZPWmuq7ww2YDBCVXSP7xRwnv
bkB86ID1HCLzgn42DbJnP8EpZS7b9/vwOlL1O4Fbx7yFIwQ12I70mkV64YtH
dOIFic7/jzBIoX52dSkrqdH9GzydeitsyF38OHtyUdnxhd9ls04r480F/oYz
eb7RdIfD9dE9n6M1yJc1UQjpt6rrsMQzhXvXVxWGtXx9Chi6au1rONQ2ZRU2
7synjnoZiJAPfTcY6i1WYiYHXzZ4nHeXleGslilv7bMuGds4JlUuBXsYatDQ
uWp3HYv2baGfbJC1saDoOpZ6wZgT/DL6s612kxqVD5gAlV5MW5yMOPTVtgIm
wCDnjVZf4dnuNnUObsW5Uk6BV5GqDQfEbA5z/Jqq4nLmzXGX2R5EL1YwggHg
1l7+TeoBbA5HYrOCZ1tYnMuK3rWW7h6iqfxfyL3a68IeUpjXW73CJT6CsYUn
2ECvf7o/5aoF4Mmp0zGsL3em9eSX+PNWFZ/MOWs/CmcSwrYi/cux2y1VNg4f
QsvIa9CPh9gf9nghti9qOW9mT2k6gQfN3vP0KuT6QxdHAZzKGc6y7qcCX5Lc
2Qdt4kqm8fr/HJ7HA2HoMU+g1clNbE+l+c/QrWTkneumFWAYRu+GIOPazbsj
yGwtX96yjBCKwiZdPKCry3IW3Hm6O+a5p8QnW62uThn9Onp12N+eJfbZbvzC
SNX9RXgCQ2Tbdw+ZHq5PCk0HG3BbQohHDjlIVLhsoR54v/3lMMzJkxrNGLVj
NUrgeKwvZyyFEjGkfn6rul2Kr+lFv3lusGZo50R+0P8ch8YSV+UX04SkWvhG
IUrOLiwBE7gFM2qth2M+Yt5M+yHRVwkGKsxjkFU5NsTRgTxn0ite6gXEW8Ou
bVVwubGxz4i4sSCsNbIluPPTjFSdiaKhyzBW3SqB5VIv5DoMURJeqPM4/WyY
RhtOi/HfYdle1p2c0E3YPvfg2r13EaW4uHj2ueuAzJXEy0I4+X/oLQ3NO9B7
Fyvb0gK/kg==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG0FODxuvZIAoPhrfRpQNXxh6azi6SD6xJNICgRf+3S7XLEb37UcCz0C0RZieri5YSmxJrZis3/5mknmyX8+owI+kSluQoy8d3pGfvue7NP2hNrYjvDgp6pclzIRgxxZicgkqVBajvWiyWgg/xxAiUyPBgiwfgRAB7tSCUPxpqT1mpPY0iyQkGrUrf5ybzt8D+HxiJtEfgXQ5aDvKL3FOsyBIpRQXQxcTkOAA5l1ZCUBPe1BIPuOUjQ/1I3zULZLDIEVTzBmO/FS0i9V4TAEMigTtNkbPYAdBCmi3bN/Vm9krfPj/1/ha4CJZYJoTGmwLZR/7bUb2LUZMnu/1j0ANJI6+twsOk0YDeuEWC8iC+pck+QgI3B5aN4dvU6GCZHo3srgWrkutqpiKOh8Af0Uo5L1GLxqWeCxD14bY7pa4xCDNwFNxwncKNjHxim4UVfVoIHlXP/dil0mKJAuHLGeeH/Q14GxESpu1yPQ2fKZwiwQK6pxCPrhlEV8gZNpdtoCrVE7Re+IDIQCGBbDTLBrTiVOq9JsJVJbt37EpuB1D1aQAXKrqu9pMvqrcy+B4qml5ccjHEuNHP+mN1fF9KTSPigOeXV5HfdtFYDYx8hJlTxn0pJj/s0NP2mH9CIF/GhtMuVlknfTOoGK+1+jWUHiKKqyZs8b3OTyJyLLCrTlOxXd+OvCWC5j+qU7MpVcs1U8qxZyAqbkQN7rNkrQTw+UZnFgL6xxBOFJW8pClVkSi7kvf+Yj7uq6qzZ8JCW/lsuuJqFFZ6Xbwc18vU+GDInU3ZgJ"
`endif