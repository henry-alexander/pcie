// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fs7f5WoUROuNOAdRPGtVY+0ahrbFhLYYFWVXU1PYyCWhk0TxGuV46IxNq/dS
ffl6yspI3Gq+SKFlAAkzbgvoVjJW7TCdtNOrtQizTnMwdpLdWhtfCn5DsJmJ
KgUgtHkewwXOl20RwWG3uHavI5cuqGR2Wfz5icaLtg4zgBAfDbIYphHjJtfX
hpdQmYKHvkqz7Jf0QtD6qsrrQryBEYqb1GnjhvCvNZ3WCp2XN+9KXVdz6qXT
OENp12eKA570QKZ+DSdQKV82zwtQD9Q9ze193kantHcTAqK6hP/biVyYYhHU
CQkCWRzeSDmtlQ0DXuukzONYcJLnzBL0zKu3YTej/g==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EiVQpzYE/hFYpZsoj7hVyFkNcuakBtg7XJXRCxrHf0COkUdAE6/LjjmAdYlo
/e7qEEAH/PG6EK3ljzPrAMVrrw4l94GC05cvS5mzzm4iV7qyjPG8TzcU/iwK
yy0kBBB2JYX1ocnBleUMTJSM8kF39ho7vWRdkPRhTplpS25nMVRg9cncdCkm
G+4a1/ZoluLPtMhNOqzwHT91MWL4rMixCNXXC8YTx3EPgANzwD5BLYIOUV4z
z1HBfv2muIPz5qVGtK481LQAHQTdKpLTcHSinEIVBmhue6CSxWypMr3Je+ms
G5csfmJQe1tv/6QilALqubCi+gFZablxmUaGSuHxjg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
pfhHz1uFXQQYzgclfK0tloeN7wjEHfk9U3TkRxAyYStxu8uBP5uN3f4Whx0n
fXSuxR6WjznReciiS8v+4xbDEFqzj+KE30N3GGQJeqcrq1z9LZQW2yQ/9CKc
LuI3xfueaideWtX+f1QOpVoN5sarsghBAY+KlgQBG7yVGHMEDppO2eKJlM4j
RRIYdBXfOGuzRltjqv7ZFVKimRv0xABzn6FaSVH/vjwMldZasn4nUiL/CdqQ
9ppeFNpz3O0559g64STFZ814L8WMyTqfGZnsKkatIxcOWF8e9+mDvrFdH1ht
KNTwx50GCwDSz6jNqsAPCdnSq5OTdMdRbW7t0MQUiA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
FM2XZQJxa/unFNaeC24Er3T6XXiJ0eqwCjMgkOfFzLTCRhAAr0Bk2yI4spNv
oyfbXxVf+U0cE0XMh7n/583i3U4U8AmOvXpcNPw24fGWTvXaLeY3pWaLJkhl
KyT7TweUrvzGwBeQtSBjCl6mAuMclzrbjXx8vrd/Cb/1WxUzM1I=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
SZKq1+yd8Q67reJuWuDrUyZHfMlQujg2rFaYkU4VwfaqE20q50jAfiinTjWi
efKxgqfAJCzpVxDDSb9ZJOL5TqYIlJKO0Fgwh5UhZkpBiz71jGIJsoHnZoKG
xfe/GFEJSjYMhFV0TBtW3DOweagv4XKhuVC2fQrpL0v0PCbNR/2wJvKie/Rq
vNPFMBJg9Lqe+jB97JNm0ckmyLtoFjwhQU4V5EufADf86f2C5BXMsHbd91CD
9CpypDHXoGZJ6+OiVUhWhlwysgHduNE3KNmhAf1NJeRgY/cYZlAkchr6xFKV
3OrQamXvd8Drae6NJmODV1VX32wy6DJseJyOWLgsDOog2ukUWNY/2yFvkErC
+OE5NC2LcXrkPwBruFL0jBy0O7Un9NUToFttWiRklftPIPVdibUvRGHpNiwL
67ySucTvSqD79cL/QXarZddLPrp6K8Hzv4sho6v6OXXoK84ELh7K/D5WvEe6
8s9ZN0SUOfP46uTGlH9FKh4OSUh/GuLe


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JoofyIzqcIMY2j4ZkxtdPVfUNOHZcCZTMDGTwwclhcklCfISg735RcpuMGwz
j93qaAgOATii8n9NNjUCGYXN5Qkgcaz3iEP1r8uGV6Gti1Vco6vuoz1JFRUs
eWhU/9kn8iJwt6pztuBqFUMC3BqssaavLPyQRE8N6ybWZNSDhoA=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
q67r12ugWaJqe2aklCFmnOLbV6dWmCfw7U4XS5VrQaTf+tt5rtBABNkmxOTC
DT95MPfgH/ta38oo5M/2g+mCyC5NZNhkFwjUhyChEbeENbGTC8n6pxbWLGGm
pExyE9iM3jz5nMaZueKhjhLI9TAkS22P11LUjs/oksdLEIcbLE4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 12992)
`pragma protect data_block
h3StGglZuVUl3Ts/fnwirQRkXBzJX1LPQILAkcL9m3BR0fKleia0/dKtaFcC
LXJ5r91gi87TEKWkhZfPs/iaUOJH0x0kXKZ9g4os5ULdgF66+2vf5uuqwuiL
SRl/hyguDsQw6oPRuyHP7OpIP4QBWveYXYAR0rN63GpzDQxPNGoZSSaPyAPq
FXYmtKj25yCI3eT8B1tQ7OQDNerss9UGpU+FObSkLvrKbbT6x4xhZ2OHj4ru
vuJ3d7tVwEvXP/U61d2rXqLO8pH6FxyfgLZrh55ZK0aFrKXZJWHIltG+AQcX
jqogpWMgfEH80vg4+P1cj7Jnwiupnfl+n11cANt9bwFD+hYLSTlHJ/pbxilg
hk8nvQtZdpYO9AshVRAPF6v/qv3slUzRSE8jypUsVvNo7paqSiDoASTzGM0V
ImA3NasOq1h2trO7HYwezF3ihZiBem00EnkohP3Uij6+di59Qyhy7LKLm0v4
zCC2XQ3yB9CxUWQoCiPz9j4K8G27F5aYfzGx+J6uHd2cpqloTD6NuJHF0VZM
1HMolw7QVwG5jJz07wgOL49NoYApHlP1ZGVYcjMpofmrBYHMmDVvLNxBB/A8
6/70Rj1M4zLmHX+NX89PkQotYaoUkTiqB1VWLFfc95rP9WaO0XHXgKuVxlD5
mhDfwHzZxQU4WQYS14C09qfs1wR4/Dni1EnekFBm4fNoYon4UGSQ5EWfJqg7
alhZtw5Yp0ZTC4yBylxKP4cuw1tHjIswV9XILnp7w7RmjqNjUA3yYG8LSHeV
aziDE4vtbi9kpIDdoAIHTbm4ocg4CMhSgdh0yaSOLBjsv2w0yigh+vg80AzM
7+qULArI3t5xCZCNppYIM9xFfItLdSJ5by8HjlSlUXFalat4E2IzHB46BBt7
J0iJDyFr9BK/Ndud3lHKCIWJKfhz6wxy7cHGCeZQpUQk6KvmCy4YH3R+lMyq
cdZ1AHzGxhCw4nmxNKOkhxQijyvnEuEEqu8pFmkXu1EFYQQO4XlNPYdRYfuZ
A3MIHxm+8W8h5cl8b5irPxkRJO7uWzcUMMnERJmcgFcmKdhRb1JM1davLi9Y
Id73vr2WK0IsLwjO+i+8GitAcfDmlAa/0/DZU+zhlR279r+HMVXxP6Ahlv0o
KV4iLkXnFfgKfqJAEMyh49VvfJCN0jeZB2aYje00ql8Pt017A/O32ujzxG27
qEPPjRVSqcePzguKtWpN/MUAZsQBpus2VME6LwnZ9s7P4N07O2oaU9PrbvYa
BsIU/NaRgRVpvY0q3ZgbN3CRmF/J0kp7ufvJWrq3jVtxYWfELrmi4kgBmvwh
e87wpo8WOuIeigDAn3A/+ihNFVlDSF2aJ1DFAoA8ZAKW0slqzLw90hyLm+by
deuk1AKPxxWhRudQnHzvecYqSN1x7skPzyZC0jFnqjMG23AjCSsU8MAxCtNY
tRV+deF7fgx9vkZciaNsdY8WjtExloKwZhgatdGREkdZOOKkb4+yQRY4XiUX
cfWiI9FR5BaWg77ww1P+xBeSsSp9/atlT4NrgCt5mHklj7mx0ygU09yeDVuw
FA7tu6ni5Fc94mmtbaV9DQlzk2NDESXAGVAihhCkYxUzHUUymmGDK/s6kjvq
a0HySjqdNTG/kU476DpnwzTMAUPF+TLNWO2+XkGQniU3MDzBYUEQUMz8hkkM
eZgjs7WcTLpMqk3yraP6fhPS0fjj2JmtSt4KjEz+Ygl7JT25u9G8aYeWXLl9
GILycySa2aGuZNvtb1B11E4brqulODaAq4heZGB4EaTQg6w+alwH4kCJkzUV
vkG6AD4pPKuCkVPaaHG9Vv0vl/JrqRFF1sY9am3WTPyZHXk3tAWYd6PLtUgY
Yz8bnLlZ8HZrbXNFy7ZIqYtmZWESM96ylYHqnoOH+5mmenUcF5E4ye0g+ozC
9Z4ppP9VnRCAETVNtkalIs2COmYjAT9lEoVarkK2Jlyh/ixWBqFA1w2xTMwJ
VeUo1Vsjq1z17LlKHPghvjM7SQbE8qLfkf+ijY0lGCZRZvBvN+c6P0H72QQN
2upHYlVqkjckKHbBybyVhGUrRvI8EddF5RipYLc9VQHWXo2b27ZO2U4dheU0
DhKVl66EMazU8FDaKdKmou1876VRCN2s7yLM70fo8xbqrqE8j/qoRKFLs6NE
HDugPxgP2aOJCdO5nWfXcwCOW7UvkLFefvWNdbzOnsh+RoKCrOPUyRw/gFuu
IruBA7LdC6COW0PodDr/KIynkgpm/YZEgWT/t8ygyX9fjrqePsOIi2BtwGg3
/vWCJ8HQ7v+SnwJmINaajyTB7mD/54Fs7JRmjgnpR/lD+bFIL4BRrshphlmF
eY4MbsLmLy4AldYDCZH1HrSWSim2fPakcYw+d6/n5XO/EapwNrU6SCB5AQS0
78tmRNuwTFrHanD8htUw8mpk5Td5aCRdG6Qe7cKL/ld4UOKgSF6iG53ESQFT
ZhGSJcuMAxMuuKv6cMy0brmF7Zq6OgiLSM2YXtMSWFsi6OuF4EAKAnFME8bE
Yuwvu3DfLO2nFZdWYzKIbvFrFkZgjM9Nd/FGEZ8WPn0Qj4uyJo8T2cO77KKB
+8I6GeD4s1vhXJsR87gFP0kCuaSAzK1DPGmrkZvxMQ/wAwqoK6ULQWJbj2M/
8RHqSCq8x65QTchsgxUFWn7gEALYQDcr1hDdPbgXhz/bL4etEizlh5eIBon0
ySd23Uf1LNQFLlPfuZg9C76hBiJezTBbKdcnk3PBHEysFhx03C4XDFUkVx/t
H3VT6xWRzMB8HxH3MGm+7iocdlAQLjOTMN9xEHMkkAwZJx0IBwPl7qUmhcbw
gD5JVkqqy/OjCmdEB91hTA/IL05YtGlV3C8hWtsITTgwhTCEnhn78OQM0N3u
HVDPbakxS+GU/FsxpzY6+jwwKFYKpqwCHP3d+iU2DyQ1qlC44pQBDr8P17DE
zHfonDq8E4uJGpG5xgsogZWS/AZHlOrj1Ke5em011/RH72YmmoHCeQuvKLbr
vNjDGSA94I8NwKzpwTgXqb16+4bWL+Wxosgbp9uDKvjmWmElypxXHYwOAQeI
VFejQ72Z+Fqe5Gv/ANKmlDYBCNp/745TQAHmt6YJ/wPvKEIoL0CaJY5klQwj
VBxt6K2yKN+rDu8ofp2FL5ZsYsuzRsNh18rhpmv1wbX4ISEj2bT0HdT6ADDv
5nZkvRDtkPz385s1HbcjEFcPwWRSYIKOU8mMZKy8DsfKYSUNd7Kk/tU9xDQu
k9F842RAl9k1HBIJ/nPj1NWxDtL5Yggsm0UPA6WHmYJF4MSh9/vlLTRuo3/D
1sgKT0WWxZFgFo7LoDdaKiYoFn0/P2dUpykWDmW4i7m5BBJDqryF6WdpJ8JI
RFdoS7lk5IavZrKg3kQBYRdwqrvJHjVCkts+vvIOVfASiGwA1ox9Btf7M+xE
9c1ANtUlcikNv3CZmRF5PjQqzBrJMvj+AwpRCZlAJyM3fvO4kPuNCD/73N1+
ShShqbiqc+C75cLorXTrbVCY+zSY1J8LieUU7HM2odWbjmAd71cuC/ocWJ6c
o9jplogALUbmHd5MpEH9V4o9IFI8AiFVYI3/Mok32NevQop9utAYejaokK9w
oBHglvjDL07pTwy5j3jp98fnzLCdST709b9itTUfcFnnpV3LILFgT7uyXHZc
VTReiKukHPc14WrRPh+geMyBa51dmEUM33zooTNMxhi2CprKo58e7hMySDBc
JQSh0eRORSJB3YSPPN65dOEZaAPYbA3WBA10+wb0R8IYtf5pC2wvgHSdd6n/
YSap5IeEAVrpmica90b6AYQcpQDXSFzzdbExwiCwbXCKi8lIkMpmC4HtNQmH
XpvlKMWjojZxot511SdG2zT5qvkCi2urzTXqpToHOtUXgA0k86Mx1yVtIH2U
wfQdsrkjQ6pdMRMi5aP/U4M0F1Tl0Ub9KP8P+XgE2NizFOp9ktO+pXfY8wQx
NXgEKODNXctpfgfHNJUoRHMVCqTUrRTNd63uxA+54XYqLKXmNJaM75lNHIt7
9DcBPJwgGk243EQ88Mz9jajm+cyTbjp9bNW8+xUHNLwm4clNlzjeMPT8frgK
AufIPLp7jqcARgr+YBFKrr6g+te23Z8NtTwS5OGpxCouWPhFs2NUzNTfSWjp
xFLVswLnCI1A4tvLY1UHaochGeiEjCT6EmC8p3TvBe5fmz7X4fwihMpG0hW5
Trw+Ikp42nmA9pKNt7zcjRgRv2WE4x5JAUmZrEYe4aluy5zoFDf2Un00qMHP
dZ7jza4kSysr0KhTWRqoca2/hXr1p+SL86oYFfvCjS/BK0reJQmBpEi7oz5H
ylk+5KNS7hpLSI/bY/mWuGPhZ/EtdROwVIXvNgyb/fxD/I3QgrpC5pWW7EjD
Z8XpWjZldCH92Um2hfQO3Mm2PTZkqi21MHqbI+R58VxYmiPZ+JBtEOO0OkHo
WMTasxjNHx/okZrke+FR46ne2xgjk6tS7ktc8AayD3eyZ6Zdc4hYH91E+l0c
OO6h2MiVJpqzII2buYDiXYuD+C3l0iFz3iffuGhXuo9nyk1SAM0qK5epPixe
WxzBc7L/WvoO7u+8tV/a7ej3jgzOEFNR/02NiaFK2MInSefQFwDZ0fuCR9b3
E7+Aica6qbfbXzV4HnTVOVzgRUiuVZmN64ZE9oGGe0Ciy32/C3SNl4/m6STs
i8cWJYuwAurOH3L041fPe/vaWWYQAyufX1y3Il5WsJQELwOM5hoO/pc+umFU
9C8NWgEm6amgGTDIHJqe3G442aXAKwLNc84x9xagQj496IoSFWUu8YdBJFAh
4yEbj28A55WSLOCjamhgxd+FpHpEyukIlO2zWdvpPbn2Ttq+6hGCMK4a87J2
kQfmojjjrkTtu76O+FJ5MdpnzBhKGDLNeWbRG24fWt5h4Pv0ceGY0ITLU0+9
4DoSDKBDLvBkHP8QC00fONL6OTAiH3XMe0j18or4MfhhJ2VisdPdVOzKowDZ
DkrodT8VKesDpe9ZlMNbzDJM7gCvhogAI3+CIvQWvZIcUdlvSooUbspF4MOJ
Lvo9VR6sXbMZNzQIWOEAv5Dd83MaMWp0sQVoz8xwSUZrFraIgihayktXHQWw
y8TBql0gsV9TfUx3nHg3yeN9ItsnTh1Vja/7HRQZ34wAj8seCwcJPkA5cwKY
6MqCPfBOmwcguCEKkucwJI2lZv258GAMB6t201abF9xNj4YV4og0FDYkQeTV
CGiA5yNA2jxFwzBrihGWI444xAy3V7Pem+xKfuQZovDnyTPfGoxnWnqksCZe
DK3M2YmnaF8x5QR9bmy7H29TjTESVPh0MW3g9M0fQMebXOcr2fMHOdjXUHcu
2jIkjvNGqiWG93OSd0jobkXxAvhwLzItbE3QvDhojLrkAUR61miJnF/9p+D1
2y7RRHZjlpTBHunSDFlZleAfG4aFi+80vdXZY+UIw940gSWSa46i1ycTxDGk
D0oyS6oR6wwo8kZ8SV8WP3emIjLo+QjO1HcEHOSoqoEMh4OP8BIGOFG4FXkp
Vn723fZwmyHszL33n9DBGiJGemhSVB7kyQ3ZAtaTezAcCyXQOHBJ71wDQv7n
LrE6kx8Tpm0zdQToI+Ftsu1+E8jydHYAtAbDbAEiDydob2c5mhf2N8nFNOOK
ksDvwFuPmqCHlhw1iWYIhP9eFGiicaY0qgyMLY4W/CJWSYcTRhvi/+X9gLdJ
wuQYpNXyf0102cOaSyg0VIweRuv5HfRDl1I3+tIgodTkC7gxoqfXI9OV/4T9
XXSgS9Wp9q/TS7hUAuVRoSyDVZnvq/PgBx1oDXbuDwuB/GrJfR4BU4z9ckbZ
hiTwz38InEkWYDQCo2PyrlrgvvKDx+W6YYICbVlFa0X1dB2XB8Xb71AXkqjw
S5gziHkYPCEWrCDY+5Y9gJSePxI3ETvkp+KbSK3U/2YaeKWW2tIFmd1Sffdz
LTGLEaHN62EY57cEJTIIH1jgToqQswR35g3uFemKoITaJWuMqxdcM+ilXpHU
05GHryizzkQ+DoCpO996eOzcxb77HLGwHGGsdIsJTkTrzo6CgkW2fi2W0Ypo
PNE+ioKZTGug4Zh8noJV6zLovk7tDurPu1cmbgWD1XQqBlDKREcBylH8yLAE
ZD3weouQvIZ9pUxsYPbCU0GwJAY+U98OZvf2ZCXrbM2tIvGSXMjqaFeA4VUr
UFwwuKoo5yKknI9gwZzYtUBpnJ/XC9Bzg8N+IY1/6tLvZAM73BVbWncPNgB4
TXU5tcNgvY95yIYS5ajWyDZ0IVUkM6cIRUM28GLtOQ4PP/ES1dC//9jZ6aIj
YgSHQllE95mXqkGyjxqcFYH5lVaRrYIKpZ0O49WaLmHUWG9CHe/Sqy7XDdSL
rd831+OTmTfptIcgKZAd8r9jb7BuaYnBLR2q+mVbWJcAjqj+jgxk8hR1jEjw
z9/RuFANxj9oGdwujJUVYSDVsU0qbl2+Dlq/EI/vwKdfch8keJhhnK0udUNA
rmPQcCEa7Xz8jRbHUjud3tGBLnz2a9xJ+ZnmXNVI+yFdmo0XCOyFp6+t3lUg
oUYRyak3WCEvVbzjVhssw9gx7aIuurVjGpYM+8eLkuw6foqBA0BkoChu/1DU
L10ArfYtlfiihr5eGjjCkN2fQsWAF6XixfF4SLcg1eYXWOGhsNPRk/pPG2bt
O4NSctOA23u8bky55isbX6RJmfnzgLy9WJNByshxoo/uw6PoNKgIRitmrZS+
C4bp5ZKmjo/SoQv++NyOSaF67r7vI1m7F5kRjthQ0Oqw9C5DeipIkIo0Jczc
ge4ZWuygKcCOcRI/yVQjh0GEvwOM8ldQp9w7BbmMU/OdP+OsCwJ4cpiPgoXq
AIJR3s6HxazM24whhizjVFJY20cZlgxB+S7liPzmlF9oSzfSCYX5olLxG7LV
FuJbhN+FuX0PDZ+JmXm5P4mGhUcGCqBTPjBk1PjIZbJPkncxfhYMNqc04F+R
UnD3aeb4/JrZJC6DdHd+WtU4Ep+aLiNv2F1o8etSltFVafaN4Gcd0J/ZYURx
IPJ9i0X3WoyjPZugthlYwOx1j+RRp7Ouz/ciPSRgzUTt6XWvE8OBjTl6JlUm
9ndfpnV5OFGY9nBAQ/tuc3YiUhqDIxrQNb9rIarkd+4B3/xpyrlhS2tu5SI4
bx7y7aaGzGeDun3iKqP3Td4WiHbwDEQC/FvMGkKQyD9wFNwYQKEUhRRcVIRS
S/Zh3tAwiuR+x1CDez3ULXlZYcIR/WFMcNEVDB5YBnUf/DInFTQyFu8khgW5
MSi7YyvziiW4uI0or4i2HyJe2RPQM35+JkghVL1Fb9Ma8lDuU06LzmoAqzr+
efgjGu09fzgSqbJ/9cAsJre6+kwhJG0iFqPi8AmkWHbsdj5a7QUx9gHS2vYA
gHveizqLiO+b0ZnLngvVRFTyoZCchtG+qa/4TtbdQjyt6HtoFyDh8g+SHu8x
pebYoJFu80qjL9kYdIeu1EDTmBUvBll4gn1g6a90XSYlJrpDpkEkzmBpOLdE
OAAk/otquy7w/DIh8Ver6BgirRfaS8v7FBUe1rPPqsA4ApacBjuxQlJIuwIi
G8syEZJUdY9OK2W1If6hmsUxM4hHtZ/q5gqzxTJadokVI6vUFKxoHwIqghzk
phCkBeXF6+tCg3R1bAcUu0qwPEl7DwDQZf+T8Jw3oQTfpi5fr9Ed6EbpW4mn
0ii7Nn16TUt1q23j7Va/XCTdjD2eEpeRxMd5yquPFBKhl4MTymR0rmAdplpW
f12hrKBPHSTstqi87YbjFsVfsFL2qQ9sof6IjtX5tqvRnbIrOhzCj+2Wtkz8
UF16YURbh8ebfsvUfJLVCWUA+DHYCJroTlRb4mo2xMOAoe337s5lm/+y9rr1
V3bFSwT1nd1PwJmtjbjTVwzurwNc2bT3ed3lJXOHl84pYbqjZtaiboumyttd
TpPJwfR3ChdWdeaFxen11cPl3ga4duXUHogqohDVD5hUeBmXwKAFwVSe2QzH
BwssPKZi5x9LWvMFfPg5p4ymqQE2UxAceDFqii6IWkCN7up2YZcKRqlnzUjP
Iwt24Z4JhbNVUeiX7QpH5TTC8pvqOLNv0APq/2rrvyG+6TUrvaYY96xCLKpB
aIxpCXUNvbPbSxAcNfoyW3RsYAbrJxbgEVA5672PUMA+RBAbCeErXmkJ1QIB
JCtkUYsI5kX0LFeASWAIFefV5UKjs5KJ6RWkjhQAKrOtMgma8+eCqLjoEUw/
VqMNA9JBZvEjfpKDA++LLATWlAGjFV7QtFqS9QFMEnJnGtJgAE24ZNWXOOLB
TaclmuRlW/DU3o7hrxc5FrEAyrJm98ixkqgixEPS5mt9BSQSN57qJ+jwleC5
pB/4ylaZQJV7oM0WpCpsHZ3CiKFCu6ck+JwCojrYTrVSCYcEvZFs2W4c4A59
kjly+8ktCC1cRwqgjNAljNyFoxGmpo3HjDb20FTPTURgXOk0Zvc5DdlyLj2y
LA3GDFPNKfS0f1WnWBq8kMZz0Gj1YvihDWoZpHIxM/KMJay9bfpXvMde8spv
RNa7WEyI8C0ONb+lmGmfz3FZi564E1K7e4aBmUeADqltSb71+m/QWcqZiUAi
+13relSXOco98Bw94po/Z4QlfKmNzZ+6IhyvtAQLAsX5PmiR0QIsgCJDB5PH
ClSnekltDitFq2ked9aYdUrRytUC/bBPJm4oC+Epg9dCvVCUea8kNcbvlYqk
JEvMMUWIJM18II0vAvme9mwN1NVwL+q2Co+MeqSHJBmdSjuzC/zBCCLs3SYN
a7Pvqk0cOYOTzARUAg8VWvvUvE2iVdGLkAtbphms2NS8AxLMMNG4pH7ITmee
UtvllfSs7w0rPGc0AI90VWyJg9Ivi549WjOAbSRqvsiez8Dt4qJhBRStG4vg
aSavsw3njyRrlgPWP/KcBxCc5vyhTy7bj1gljNDjFedH+UY/6Wn8h/kQMovQ
TxHkOvmQ1zY8ZxZesN3l7zI+ZiBeo1V9KImWVFu6mHDqH5bEsGZTwv9LfF2p
1mE9TzDe/PP3Ncm2ZxWrEJjU42k6/QNfC2+/gb5dnTL8aUZsiyumhZ+lU9VQ
fv8aJUunB/JAWwdszt7IsKGLk9q+XiuT6fDfLtxjCn3ihukII8bE24O8WwI8
1RKrrg+SeQvOI7VFiR4cpCFHikepoNTAPAqaWFGeS31R5aEEtbi1qVDLPSK1
Kuz+hme4z1v2z1UChWz4VmV46MSDtFA9rpZDX58Oxl/q7dK24gx2l3EnhfSo
8+qBtybZa6S68rtlNkBGEQU/nLmYIedXJw1DltcDbLV3+LyuLEvQgdtlLa9w
oBTuls8AMkYNV1+sdEYGx2ofMEZ4vgFqs4XF4F1dXef0PvLzyOi6LXUlsf1q
UCDaVksh2HXxx1Vxr5mqir4A9VfFQ7e84M73o7jz83q8xA7qhf9x0B2FiGm3
wrB4ojRXhUQcUYM19DUWILU/bHu67kkpXSVVnyOpSkGgpTD9mAXdc8MvhsiY
kpA2wrWJ2IpGa+uPEIqmiOtyYpJkEfnkgB2yjTIWbdBHhm9i7rQTcpuQL7u7
kOccStTkrbJGn2JiEb3rXYiYnqZ+HWiXo7rk1qJF1LQ77gExl4zAcbpDDX2J
R9wSMuwB+BvaILFqL/hRj9UwvBLYvIUMYLyL8B3qrKagknoubG9f5XiZ994r
v0qCS160W/ZssucoBZ5ikqpv4Pim8PV/9rJos92rMy8SCmS0mdLxO/nhwqrT
s6YxBVXilmUXQbKnDJMOizBCg8rlI4AlTQoNuOvHltmv85LsT7W0IVRzIz3R
LTuSUL/D64ZHwjN8qZ8OlMFRGVKQxKJ+EYWnKpwUfAojpjtVYlEgJjAN58/p
Wbm+FQUD6E8qksOcA0aHWc8hlI/xOxHC8k1hUCCBk4t8WJ2FuepcCOTWDTVU
ARVugdvqHhNhl/Xr8M8eYqbNWP9GYUTRdjGtgGeHCuqqsx68EN4oduDrHL/C
/0tFCDV520aqJ/4ex6cSoBxlE28VxXxMDqBE5qvlZXWgPQHRPbY3ZXOAs/qu
lRx8dKeF4jJQKMmnkm2pbXcWn8nRKlsPxoHHZ7k2/Hfj8ANJD+FckJEYIqc5
PID+hjVK7e8B/hWcYsdz8X1vIRtyZ3Xr/c6XyM36MmqV/j0M9E/LhrRQCZFd
VjaaaHwZZdbFo5b8SVV+eFPmK8p79zXZKM6jh1pKXOAmHYlTD2D9p3ETFGLS
SkHOtQEyDO/bA75S5KyX6GVWxyxna7dg/T4Wu2y6mXeYweCRkakahunG4QmI
1l0FGTsIwxHMxUjIuMIQr0IDYL9tP8pcYOEM9XbhfIxQKlVYFN2qlOlXBRay
RYe2N2UJwMaIjqRX7oL+7zEgBm0NuZrh/55rgPORfwhtLomyQubTCJd8Xcu3
x1Za1NK7CBDr5QrVPMpjFUxz8GbKxlei/3BBTw2QgAFotqtGlQhvQd+bjSUM
hmLIcE0iXzYAPiv9u/nxTwoWxIN1FPj5QzSBwVZ+YtmfDmAZl2YHcw26zGF/
nAnnjAm9kXjMPzTe9yjuYskXzLwe+TLr4jzh1GBY3yxA7pJ3RbE238HUtvql
9aOARnYBUH2aBs+qryghqETI43vjeZwO8VMVv5OXGKSClPvIVKC20RRv7vL5
CUMo1CoYLvRoxJMepfrGFoKnvQ0xqP2sOPcUc3HglbvsT5gjZQsNfhtXQM5V
Z93pkiVwvQLiK/icglbdhrJAEOsC6G7Ked6IoRLzqVrGbfIDv6n18MQthOyf
5gyGP+2RmWdLb1bjWTfwmB9HG2DsNEhTMQEOSFTXrnv/zAA1dK0vZvb6kSJL
5doyJtzst6f7Cv/HIXxlQdZQtLuo9iJ/N7Sof58f0Va57IhO9gWLRUThAcXF
kpjkH0VzpfznY1WEX1P0Mjb5cPVGqG712iVeaCzyEn0npmSVmtiZjDeq2/Xq
kPDybVnMwn2gC/lghkzd1BonIV5Ck7eQo7snWC+smFF4aBVXkLvhLdsV98/o
QejuIo8BeRHIWY3aMRvxR8udFrtJvyo/Qg0bOpy/mQDyOvn43wNLltsXrGby
8o/qCQ9QPbRGskyGlqMn7rM6YNrTcc8ORSZHUwCjoDJBYsQE5wkfHva9NQKb
JgN2H5KbKcKiYtyuIsdvdaVOx8le5zx5DjK4aHsDA53ExBWBaUQli0TLoxhc
2M7aV+TjPf9G69x7ojNDAGWRKCXogdef3LeSWqUhEL/Yj5gC1PgEgiKAqL3b
rFVjFy67lA5AyB39lj7EgN1/3uZTli47epLQsZcmDU3uJni+rHwYAA10fbIO
MsmeZHbPMNmU+P/JLyRutZeFoGcaMvpKD+41WX005lSe/B/yM/xaHUk2cmGo
FXPjYWb0HAZYjk+AzS0i0yq0jLZfAj9eIRCY30eA+QVg1hmQR41An/6tlfpG
JidvfXTfX2ihDMHLHGZh+0tMjZ4Zx0mnlQ3671sZCNdQXmH+sCl6LmM5NycZ
CxHqLBw/MIUVzhQZAGCSkUIwv0UgonDkprM80iCUklya8FZM+UV0oCCeO11n
zsE7dxIqghLIwil7ZZAqA2wTX/iRTJBWdsnnIOVzBptEmcH0AnnjFShXpE6N
QlvdxR+eXnTtH41nfTRyXvvlqjfQCcgsCxcYncAaFLD+xNjCK3vRx4R7rHuc
3nfAZRHyCqWjkQv9qSLPH48J3+PxudMaUbhLrdSw+0CVt8IjDG/BsK8BakL/
inP5EZB5KAcnzGInIU23sNpjRAhxjeGjOYHZC6RY8hTb4tTc3X4fZhN3Wcci
MZV/tyV5+Nwsod8A9x+ZYl0bWVZjYprk8S7ap4vauHjXNnRG2JDW6z0Ji2r1
BhH7VIj7iC79ttSoBWoAguAHS6F+/4939tnYO+UBzajtiCzRWNHKZLuYsLKK
jwsbl/BmsTLlEpgZQWmRN3xKcTdxdtV2nml0atg+ISSG2XnGJzmfvuM8JJM1
chMUhhlfHFL+kzd3SnsZ88pZLVrZ3RpYW4rNB42/GTz0MB+Wldx17KOhS+1c
lwpl6Qrg+ihNXwMuUkXZSlJnyX3GQJAKGPmNlfvx1Lw8SZM9GhOqhGn4e9sq
fwNmzpGppnVYpAu/Hm4n05lh6ZXU0J2zcywVaoEX1TcUgJwPN822ciDWFBnN
63prZ2UfllTZkXgAhUAoVvmxpbLX5NX3hsFj3hEdDEXlOp1ckf9u1sqKv7Mj
r6dZmrJW0NIXO+HBUaKI5TPo8yACPUly3uLQUM1jECd1wVXoRALlFhEx4ySc
5ftrj8NeyKqyzHQupZ6ZKwwjqBgMlcI/v2HR6ghO0EqvY3mxu3k5TVZqKT8a
upKt1GCNFob/XNGVPR5PdcJxpav3eN1Bk7qe33GG6KrfXsdb70N9SQB3G4AD
jLYMeQvmJ3FjJSatoLNT3zYVMFKOXy99QTUsPMyTJ/kR678FUuL/i1cUgui6
pOD0kErW1L7BvUaPp9FSqPvm3ksIyd8xCkR8dUH/718r6PKZNSpFHJqf9SqJ
a3/q2lXOfA7qTeISjGXL2BgknpNqLuV2jmA+rb0F1CzDldIBE6G6OSq4Twlx
eTrg5dV9cF7FLfRpCwQUJdcaUa5XBeysZVoF/VyFu/5RgumaZk3HFmvvVenC
7euaFb+lfYmF+UiMBbivMMSRdNqZpCcFLfWwOS+TqcWD174F/OC5Bblq3vZD
V9aYXFjTervedNWTm/6eRwMqMf29258dxLucT/AYk53f3i6UPHE++2hITxmu
AbqYtk+388Ls8lckdjo5O6tmFU3ZYc7SfDCV2AJ8sYh5wZdrp8JkoRSm0PIF
Q8TLhvzkGNChn7YvpZd5pbqgcgiNhzWlhjX3eqFaiVBkJ0Qflz2YAXmxBDr/
2jSQ+biMixZWRqc2BKZZZyGFZswDJZ+Gaop7XbHBJezSjGkYIlfOPi1ql7w+
a1KFoomX1/GamiKTWuT2+JF9OIYj5leTI97upMaFRdD4MlQynLkzHcA16wYg
uePYpezmeM0TUA5H/K8il+Oe14GrygLISsAPQ/+pltKUMwW8KvVvDo+P8uJ5
nT1n56+vEtgmHKLdcIYkquBPr4CF/KIcOVtHoC2n/9xtEw2fRPFaT5FNvw0u
Ep8FLt1yNGEfaqVrEo/wdNDwGDP04ndZUXIrvXpGBVLVN8tmW/LaqbXkXyA1
wkkz1lYgyJFd38CljNNhme0TbHIMnGDKOO0RPBUFpVpcHzPA9REd5cwcHRm/
1+PIF3syjHEFTBDdT28tX2umViKF/mgbVc+l6y0HAfH9B2f1xCttaqOguLat
2RNY0h/vSTLpfs21h2ONCDAqJuoK7iBKGv7vD+hnnv1sCfaT+1s6AdhADLMx
exVKuqb06VS+jSniKtcWjN73p9TMFpTerjIUCE352rtk0h3oo2lIDfXf609M
AfmBE4g/vM9y5IpF5hOanuqpe2sp43xllczOdAHrXUXavFP4prvEZ6eNvYrT
/3lmtBfpUcdQ5QQhlHFhtpDkr4viw/yn7yeF/uliZWenmLkzU0kqnD9Zacxq
1bD/rgTmk38bR9aozesujRKh0VW+BWDtRCX0OuqqIpsyv2NMW/7JepM+Yjnn
/j9M0p7KO/c0GbQg8KIjLbLcfpJa2YsIFI4n+1mJOAzK4XelP0mtGWm5XJ0r
9QbwmnR6hm0IqNS+0IAFAmm6PYrnQY3d/1EC2w8+D319EyGfRGVEy23+QTkM
8GaGWPgvcW+Cj660zwD31FqLvB0lY2SAJuQu9AxE0dFdhc63HdQNx2mrwKMD
hnA/iT6BVPHbSeDQaJMCfCIoP+POZuFhi5SYh+1UPBIDqwwJt82AAGE+jdt0
A3m5b9+Ftot/Pa4VUCyNBGK+6c+ZR2IS0xR3NuYdmcw9M0g76e+fzLYZYPtS
05+t5Gk5PhPoGPKPa0aWUx9RxLT+JYuKLa39BkU17IuA8XfMCGCSuDRVOukG
4Od8Zox+pRwx9TUvPZNy1X5Vjxu94T9Jttk83c8wrSHOcM+F6KWd8q5u/OVg
7GI+Zi6EbnXzJQOPnj6Y+hoI1IHr5V+Mq8I3wY5Jhao2YwdCmyg5Y/H1GdTG
Huw7wrgRQbQCRB+Xu6RB9W/GHM0UNmrY+dJO7Q7n++Ho9nvmZt71qyYfzwpS
fdctoso1zxfbFCos8dqoUPD2Ozfp7OY5zQnqVl7jXFkSc2jVaR9CbdPSaJhV
9n+e2ogkbPFz8Ro8az0v3mp7LYtITJb3KcdEp+PDZ+qi0LxEAXfrKkE+5GVA
wX+suT4+cSulwPDjF8nOJzrK7xjuN5lPu+6Ph16H5Wr6Jvp7RLRBAzEUqYpJ
r6bYHU98fxeKoXs0U5KKDGGpZIInFaa4iswz/tdyniyWOs+mnXQzbXLdrMTd
RN8B2PlC2BSW81Z4zClUPAmr/0fm/ULjXKhrA1uC3GE6im3kSAtdPXIZPy7l
gx/mtkfNxJODOI+cEtozyEdxYTGx7cLciFXj+e4XOHFdmpX+8xT3JlaCUimE
X+bbvJjhycf7RpmNqb0utSnnedZZ4AP2SPK1KQLT4FWU+lyqdoFA8TyYq42Z
HkD30xsFjWNGnrBHPD3V4nYudmt0UiGmZufIEKsfq2hGYb16YFDAWnSn3De9
rsiOmyFB6yPxX19xUzTn2ame+X4kobiav/wsMHGDdzGjH3Ie55a4dDto29Aq
aIFRGJG8WSsFIUYyACKeIUPJLIWuz7fa191P6e4wxVef97gvjADkHnURb18f
9Usfkr2tgcMk69EYNF2aIgSDuU/XgQqzHLC4+Tep79TJSlDJYURwKbOsbByy
FVETgs9YIJri0Gg7kYk7eZ0pLyPL3TZhzC59PRF7iw1SUnCUQhkpcEloWt7T
ZAeS9HDUXs83Y+R1nlhHjdydpY4IEU7oFQQvvPIdeFMaLH+kcSXoT57zJSn9
mUmZZ6W6OSlCaIDh0E8OZN5o3bm5Ja76qxOpf1tB2GAF5em9+4E4BVs/z2c2
/CHvz40m0QhQhAQjcIxLd/Iuzle8DKGZv/q8QtPnTLuVc+7Ki07+I7C4Ox2n
WN+vTO2Wj8kNb3C/XPll8+8ZHq3x0IAbIaMrznMRquWA5/DlEcsXRHUcJsWR
GAZ2Dd1lJRNikYtmbOfU0tOzGILBDg+E3K5x5IyU/gXIsg2SJ1TL74WYDVqM
0VsXDoJfHXJx7IBSlAhKlG4rqYBI+3Tb7ggqfj3urooGRHXh5DL1UPL1W0Ug
GryG7i/K2Fhm1k0hRNo9OVW1XADej1PCA8GXKo3SIWYsPHAL9LZDm6/snBsA
jbbCFqfbNFmozrXHuaEOqTFPyapzNZX4VK5s+sOf8VVX97SfhSm0JCM5V/Sj
5S2fQAGctHWGrLu/76nXUqvSNlXeV2ZPRf6j4L+phNXN/aF0L/KT+f1izcpg
tEOxsiMaaCwe1ZLoE3DC5es2pYJLkhkCShTGNceQdxrLHBbr3bfbd7jJ1LSF
CY4Q/BUbEzTuuJ/l4SP64fKW/2bkwq7NQm+8HrfWJaoWKV6qOtz9JBs6Samd
Rne0dHZWz06ZNTjWuO4wR4DWiDjQb6bQr94hVPptu/F2PtSgWQrc9UVysnYi
lTQk/x3XDfYLQLJNwsBRyLRn/7d+gBfAKdQsuRhnnZxgWuSuqfmQqvlEUliN
tsMU3sjeW09KAqjfWeQWaND/hwp/eRQsfTVEV5eWIw9jsiibqQtTapcQhkxe
gbxCWplp5Ws51c89WmUVzpsJOea/INvZOyBqrRzTBVJUUC4gaxV+M8+7+GZO
STW6OioTYxvJJnr08irdmGVWB3lR7xg2a1BI38o79tedK4eWykTUKySN2goj
c+wbXeW2ggO4G/aGC+UgEvb25l3cTLc5I3/u8N7JmBm2A1hBnTvPirEX1Zmy
BhdZDIovIbqV1Fy4G4LAf6vxYxD1qjnB33oRWu0PcETHho5F1C1wuou5IjlU
/TsYY09JezMb5xRatkriBL2LEaWxRSkQE5N6UZr6HpXt9uWUnfyEpnTIYqNx
V3XV+pBLzgEpKfIQNtcQv+PJXw6o0dw/jqovMUMuUMdcXyE6JjGBXEdfaKNL
yw3PBi/LbfhpIfWy0Axrj7DGPju4E0orOc8EL7IoJktNOBPAxp5IpjzmGSvA
fEHK/0+wJ2Ltyy34hG4KWicUXtE7Ul/KHIMBhid0ifPsiY5zICCd89tTicCS
ZB/9JIZ2wNrelERgahkR+akXeE9wXihf69xKy+UwAoRNiRaiZSTBdiJIXyPS
OJG7OwM7yBXgG+TpTmhlX8jEkQLeBtw/B3uZJ4tP4vILysyATbE9Ema62X/+
hYF/JrM3dHbIypBatNkshJ+lDReH+UcZcpwWiHZBnXDo6L9l6GHLsxVVJY6o
Yv0gGx4eDAN2sUTpMxYykexVWPkW2wUlo1gjmGI1Wct8lfFH4AG/noo1alhR
dyJLPexIboT17vTjcShzO8DScqtX18PIC0Z7UXEW31zM47OzaJoKbJaeBFVR
osncdICGymdbOrPdIY3aphiJLwDl+hc2nDjEPCgB4s5wnwzb4udd3mRlYdwl
qrLNOvhb+CijUA9v5XXA1tRQGNU1fQ++JcFMv8LCgJZ/z5FSxCDwO4NMmPsk
OSGWawyn5js+jRIqxGN80JndPWFC89rtQduyWkEeKDlkzvQMqMItIxcO593A
Hmb+kfMei93rdrd2BUCrBCkQSrNYuM4HYJzaVmwMBAZXXv9UfisLu92XUIVq
93O4dsVlcMMT0LfBWBzV3B85UgZ1Q0/V8rKllhP/s02VPTc0Xr/XcI+RPHYx
uuR/GLHBQ4RN0va8DdjOCa2HZkcdd+isTP3qQPxcs0ozrGirF9zP1Bmc/mhj
xwJokWtZqiTypkK+C6Oh7bCbWCRw2RM8eBlLt1J2ByC0yXR7f7OGYbnMRcjn
I0BJh+IoEs5OU5H2sd1BobD4svPSZIIWOzWTYmHx/fsNuvXUOaJmXY3WWusH
zRAh1GEC+dCtxadxov8lET1SjG9Xmx1SpxhbVbwQHlCLe9CRSxpYFJcVRBO8
MjIdk+wZVEaWmFsNt/Nj3MpLHZs+FLwD+OAv10hh0aoC+uKOmntu5CjOZevL
jUX/vG1pO62ssSDY7ce/plGzkmH/kFNujcDMlvHUOm40G4+JNNwcvuoMWPk0
Tmj+Z/U0n5zjUQXYQKD5nLB8F9WMf5kwUskAO0QZ1oHpgdlFxKipWIqpNpa5
S98fqLTbHHli05+lMA3qRMYkMJ3mD/XxZ+x+bbPBFi6EONfl81AD3kvZQiqT
DB2SXmLG6mkY9hcbG6oyG9lUw36QyPtPb43QbWMXfgwBBjJn1FD7Wii2CKnE
AR+Z4kHSC5VOQ1QaRkiKfc6YZnp5NEDT5GQOBYGnSBs=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfRsdy5bvRZxXQLE/7AlWIZox70YFJUeMm0kSNOuqZR5joy8vUN+GTDfPU8Mzmixksn3DqodNO8WUl/4VJLdjU1Xc4D56VL6l3GcA3eJC7uQoh28ZWEBdZN3iuWeWun5drsp1MAaxaAZskG6yd2oRQ/XF3PrURdtSTGNpFYBYIr8CniErX+CQE89VIB6V+1txqm0ayuSo4QTnHomLcRt1zCd8tpm+UfN68szEPSZcUi5JraSSY+rKnWXs6Y4JGoLfe1Fd5rrMqo1XK7UrDl14Fav+hCvQRsgk0OaWIjDGhFWGxT4YrE8/2vxQ3Jrg0im+7wTDIbB73DTpmup1UCjeQB5wlB8nn+Umycfwakw8NkL8MSkQVgq/fnDkiYNkUWN5j8imRuCJ4oganZESRu/iO3BGP1lnz/p5cL1BaisAdcJKhxmF/LbJQEYxZOHeSNDtbLYc30J09SIRo4+vxDb5Pf2Z621SFX4poDeTubBoeG7HrJ+G6+hb4aDMMjVeRFy6Ea5uDcRNnX9v3ZGae/ET6Q7yYP5A1cPVi65T2apLX4Ee3NO6QPNnR6zpjGvTdtnuaHRbEuAuD5751CMhuETgPdsw8S3kweCmWgElkpqff5foynN6QyH5oaOh1I4j4go1+mSt/0YQ3KV/B0C2CbysQpty848wQvw0zsz5b/omzswSSG4ltEjZWUgbwzq1i+yXZOueWdFEn9joSmlzvVhubvq/sPyU/SaUnmb0L4Epq6j/J2coycJax1xtyBB+48T9T+g9On8K1EdnMWWpEGJEueu"
`endif