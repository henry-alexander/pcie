module system_intel_systemclk_gts_0 (
		output wire  o_pll_lock,  //  o_pll_lock.o_pll_lock, Lock signal of PLL
		output wire  o_syspll_c0, // o_syspll_c0.clk,        Clock output C0
		input  wire  i_refclk     // refclk_xcvr.clk,        Input refclock port
	);
endmodule

