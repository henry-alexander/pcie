//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
nP8jf7cnr22cOsZ2Wfrm3YjzCPv3Rrih51OMR8YJ8LLSjnLa64Ca6BxLGegN
9OweA9z43B0h8DKz2D2R6D2b2Sa1U4ct2cAp2XlObp45hwrnizlL2yx4iowf
I2u1mYeXhlsvmL77QMWvRApZYB4H1XLPqQBSH2Jf/RMM/q+Ndq8NvoO5LPC4
iTQTKk6zuxtM1abo9TNxAS/+Mt3b8STt8PqnVl463DAK3PQdm2EJm5GhNYc4
7grNm/Hh/+k9nAD9aCUiDgbMzOD+6xkPUBfUrgP5CDNALyQL6cAnWY1t9uhZ
n6IffIY54PjgUnIqWL9E6tAcN0KBKsi8wZScNIRv1A==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WDjYMeogmjTruENslDBmAqUqPK9mT7YFXntyN3tlVQOwY36lEfK4WH4LxS5z
n9HXyAJHnHIVkZEhObuelj/ug+JzwfVsSq4XoT3b/FxWV3X/eHIkm1bWVPcj
LeUxBFFAiZaDmSuAYFVYYzGh4e69/9AjPOSsjNFAE/tACpEf7Ho47hTfTLPs
x4of2mzVD1BjUspwxvr7dbASfzSVvV79HIyG0ck7oCfMse5VWQpGcd7v+A3F
EqIeKPCiT/zcvEHZnCZ4A7oQ9Cvc2MhDcyAysuismpsxRXVDPTVlsHfNzYJz
/UP4i0eopzqRtiRa35jsYf761HgN74MS/ukmAxeotA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Oj0++7jnnQ0ZL77s17i1/kPqv8GCp3Ye54bMVOnOQXSEOfx9n7Fy7CrXhQ9k
JJjxiwPBjvft1tiCg2VzjyWoHl5gv32BC3Sm1rRhGjJj5Jyc728dqbz2XiGf
0Rwr539EZjWB861dPjUftC1fRPxzMrgC2XGRhkdZiVxSuBPtzPzmHUSc2ibJ
DmVJHkPPfa+YNvOmVHDUG7P2GQdDmAnhJdIeICSs2KnZLvZaGIYDYbNAFZu9
lzBdfWgPIoWtb3cObR8g9bVtdftRU2StzLlcO8xhcvsR/wha8rUXINz9KZSF
iKguJ0CTFazco7tyU3+BXFvEneK2XhqL0DP6DblYrQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
XJut8tUWFkCdwd4T30fxnpetrnX62JBH2Wr9M51fDhCXJQj6mlogN6U4iAil
WI2BjIvUdrmzkNczn8Kgmrz7g6B4swCWI7oAws8+1Ajt7zqTkEtsm3sg6SES
SIplFtvxHV8ASPcOZbIsQ/M3XBhMetsIaSh99xqRoD7x5C+TBaM=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
h5haF3VN/h6Qy2Idwvb+0lU33Vb8jJ2t0/6jaMCtaZpTTKTIdbhmqOTD7pdP
mUJ+u1MwNUSeyedkIRfyMbt155io/OoDAXnm9zv5Q+PWyJEfLX1vYZehJSq0
w5+gxfCaJdkBjalV/irwy0GOjn4Uju7oQlZuvkfmy3wpEPl+1j370vmFEQP1
16WY8mVtDEsOFR8FpNHM1gviVfSGDv34fS8gcQD+FGKsPY5wammc1Hc4hNvl
Lv16fvxGjdm23NwTpLZVIcLUdtfadTJLg/HBPN9sjr+2d0NC3+LLsTKZxty8
DSEcbv+EhZXurMjMVlIgPdAAZW0sRetBtH4cgQ+oLrFo3XFPcHOaQBe4da4S
iQPbxOy+skdGn+Xprw54qOzOVACmzo+GHLZcLm/6FaNL9bSEQ9OgZj9JGuxa
bphza2C194aEfrqP42FEr79qkQT+gHsXD6sPXTLY2Xw+dXEJ2TDyAu51L1f8
D3dYIeab5QDV2Q2ugReLCzlAwUQHXHkC


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dxYoI2pfGN/EqWvBjkJ1mbX76kiJzNwklU8Aw7/jGDWDTNmG22RsBpC0ij7c
357YKk1cJYtraQucq9QBCOLJE+QB027b43kKfbSVKsW45gA0qa/1RNing0Kg
Ohfs19H/QhrdNd9VkRONlW9xTx8XhAFhGaEffyyIHAuKbhYB7QM=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
X9/+IpZjDecGafTG7O0/BOtOPc9rmDbHPqdfiv9z6isEft2XMtCCHmjRyGco
nxwCqbeEsXrdbV5/Emag7T6Hpdcd0vSoUvpfHMtAVDpZwOTrHIVlaLhIVAQi
Nx19TFmWBMm4J4QDmiGeKoabfJlTqQ8krvaaosuBaxn5qrVJOCI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 7792)
`pragma protect data_block
rsKvd6mcbN4ab5n91dO3imhNFwkYo1Xgyk/4RYL4Ab8DyXiGA/ecd3iy3rtU
/mhSG5zOf6Lqx7D1u4Y0CsOJno7VUFx3eLW0QXBj9xMEVXa7n5WD+0uSPfix
82aV8b2wPpyEQOhyAaF8t/yKqlKASEZDz0dUU65EU4PFiGstLGR7NGxc/aJs
elGRelyXMq8NII/AR7cFWrb0lAnT8tzEHBXajguA+/dXXyXGV7VLbduff/RE
4MncKBE6PkTf6sUtDNf6QZUSBmaikSVL/OWagO7vDizU7+shhheapcBe7bhD
sTlhiDiko1isZ/MWRzsUNjfX5vEql47YkhApUY90xdZKf9i0QGTTiwIg4ItD
Kksz6mG+8eUcdE+kEy3L30fOs0MqOvmPhrrhYylS56B1qOORop69Q46VZ4Cx
iMLaTGtIu882+P+uDyVac84n9xEBXrVtQ2RLokGPyaLenZe7+rQrDsSByFE5
5mZsf/MV3EmoLql5qapMThjBiHPT+HVlcbd38khC/ixOzPBf4PWQZ0lZI6tF
ZzmLG+QmM9wPNRberPle4Of33L34QzI5ww7mr5atUBAOsHvB4FNkRiDdUjca
z7QLe4v2n2hOSuJoNXio9W4WmDFU9p3i8Huwt97Zz8JIpvdHOqZS2sVfFhhl
9tpQ1iikIDoN20/Iz/ghcsaRFV/CahAUZ5syGH4pO2xOKM+I4zNrKbgW5Iur
LGXy6fjk9q2wWFWeYrXqWHA4Mc/CpozWig8p0i+28ukuxc+o5HpJ05/EI2LG
8GsWwJE5F3NF/SjlCN9i7lHerNbUFhD9oOjQ3d0cTu/BoHUvCfepLaSEpNpm
C3Hsx5+C8R8HTsIejru0R+k4NBpPTSV6Sw340e9PuZzg6OHNtS/LqqTPIy5m
Odmk1dGrNUVBsaEjo8KaaCM1zzY/h8w9Gzhj3ue2it/UY416cwWjapj19x3m
GCCUpvXer+GvtXchxtOjjvJmBcSzlbE6rVN386CD++TmCnWKw/b8+hi8nGXW
VFx+YPCo5WLk9M8qe5PfpRh9gjAp/JuZxii9jkwe3n4HtB2wo9zJrEDs/cN/
q+cYxFP5OxjVAtxrPMJBqtsBtPLBpLvS210AwJ/UXFSxBh28nKE9FmHyUb6c
0xbr/1+vzDxGvbMBD0y/2HorCLtB5Qzk/AJ7TLL5M7KkpBgqQgLjuC+mkVCD
r56Mb1ND7Rem0QAEh37fMREsSpgLHGjpG7UuFD3+m8ySxrCz4ZCBEq/BC20L
siThtKpFuHMZam+gxx2XHkznJ7YvV4uBDZ18eObpbdVfYQ4gDXHO/9Nn02Hg
d6XAZfE89YkPQjZDcSntWmyFb6E7w7BdJsDPp8ppTskhqcyLIXoi/3GmN0uQ
xXEbM55vrU/CwpRbK+REKexCAtptbo9QCrlHOZ+/BQ74AQSYe5zwnace17Dj
QN9o2d1CcPQM/QGlxxo1RLO6qa1+dITiOVpRO5HbtJPck9LS0ox3ZAGMqiYX
YzulDp04S7T4VMcneRAOQ/CRG4+7WNd9LUsTVcJlO2/oVSg41V6xjAjXwPhv
Lkat/mY66YpmxgS0V9mlV9AlaZnwhtyJ/Qdd7B8jrsqQ3PhSuld1wO+prIjt
09CVdzY0l1P2Wymk9bFNO928KSu38LsO5j3PliDZqnwf0+ke+EY2EIPUZJZL
nhkZwK3rHo1WqeX1Qzsz0Umah71qTqx9L20PCVeh2YFd0GO0uHXCWw3xLEGn
jmyegsNJ0hfPpq4P+zoQk97+k3kHugF087qZIjTO7yQcvnaMdFTdMr96dzNY
8W/vpp4fcnQK40hDW4m3btaB1UkL6d4pBWjENrsi4jtxIZigTSF7O16ePDSg
9uw/CapA+HoJsHVHo/qAOBnSuU4cGWHtDzOAUiX+TZLhuBjB4zA9WPg9Gtsh
8EbRtedll4pj6tDttYRBjsBi6giQVTy+1TImXTlHA/bts3hNCEWKYwlu7pIV
nXu5v/iFsTq5WA+TXYigEG4kswzFehE1mAjESxi/oxNn/oh+vBVFF0o7dcIL
V/6gbvg5kNzQ3+FM3ypGy8svGTaKQ4dbMs7SYLSv9GMym6WhjNsEZHjkrYem
1e5frUilexxgrwPOcUJcOiJpnX/dIE9xq05xo7GJxZ7UTJJwCex0vusz0C7y
4sqqrMjBEzVXkmLgfZfpyBWQllWZjYSy575gIEsS2/ZKcnMXmllWKKFfbtvC
mym974Nwk9sIA5CkIk5hnNvfwCHQNzS2laTAoYdV1e4h8uD3gK2Xo7m1cKv0
xNU12wRjfLotDsDVzOVtOUU/K0ICesTqAxrm2XaNrPKp54EyLKQQywvNsW5Q
CY43oURPbZDFQYJPYCmQu+DrzY97IgIV+l/QYve1/WofQCT0uwXAOtmDmgbN
F5+Wvh6bSvf0FKuOiUdCucfnmm39ophf3hE1mMho08re9VoJct1ZIw0fmAbF
51OaB44vhr0qAaRuI6pgjJNPGjcuVsdYTLLCIUdYoPorlcqnAAsu3AuKJAfL
BycD+JrXQvf71ongZcJjM/3Hzoll/3YuvxUCPj9TqZSlHIINRjJQYI8O/h3a
m68WYnVCU1wZ+owXzdIF82gjg2rAl/oWooEmsQADGMs1vQKfXDNTuC27irtr
U+QTs/53Xme9IEkEt77NbwNEstr+gB5QyBcYSaWQMMjIY5lVzimvGAdSBq3o
E0IB9A1M0QjHFK99IDMsdQBwK+sD4PzJAy6WxbXvr1ZdpRk1xoAta+M1z4MN
FINiHnmiVzmsCQe35DP9VqSZnqf6ZXFPQfe1E04gMeHsOrzlJEteWCD5nKJt
U5LSNSVGL8/vNguC/VWh80PhiNamFayRYhsVB7VQfNZQvR9ZShjgT2RdKk5f
G1NIltOmtxMnP5rsDa9dkfNP88l3WAf3bk+V8UjIwk5unBMhFCpECT/datt7
yKKczFt6gBeWpGCdj0BzTbMat0XndcX0gRjlFKK0ZcOhtSBS5Ivsv3s64GJM
63cMEwkMnLbsuep3jIrgCRenUAEs9CWF9UrJNWtzvGZafCicZ5JSq8+tS96n
mZWDThXFn85voqvERvIu0/AijyrFSh4K5zVGtlYu8ykQWbda7koduSAVmVLY
A35rNSFXdcy0PcyrzT+4zMaaiPY9Qj3i/oyJeoKxQ9c5gCEi4Yt2tkZ6kndb
SEs/TZvTo9bXtEloej0WCS+VquXhMcrQ3vcCUJpkiKEt2TQnpUO/ULtCMR0n
BwHMIen2BVooZbw8+LD5m67FARTHn7K49o8fCtfuu0vbLo6+Ne6/tvGPOH/h
YAwAPWF5ArK14m7/v8q8/PpdIjszBq6zwx/Gpe9xAzCq+FIoU/7ybYVKEaMF
9HQxjqOTcvJpZ0FJvMruY5rykI2dXVDKf8mhlPc3cLV2X1ULGuKt0ZtTJuCs
dO9+9K2j1ebRkikPddd067KRBJ9oOoOpxDFTPn/g7loiFJCHnTYpN1E1vIzU
1oRsbWCI6J1mk/fU5l/SJ4sRb6jVj/CoJm161e96HYjWWX1b7IhM99wJgFIF
NvVhR7BYuG80V+p+WG2m2tWuObvoKPpd4vb0rLNZd+fgETRY8mbuY/tozyQL
AUgg8/gFFiHP+dPL/L4f6S0I0gCT7ZHHBcuL/PzzeUAmmi9WWIthBLk4x8oF
ADOQu4XwwwnmwJf5zRgwkYXnaXcVC1iMgRWm6DthQYwbPWRdTRFSzjWGWLE9
nm6Smz5c+AmDXaviqirtlnqjmlqrPXYXLA8PicZtdg7eoPDgRuI9U8VFtiDU
Xy3xLPwo9jHlupiu5a+T8rwsaX22mPVPvZXAieUx/ShLQza6c78ZRlUgHCz0
JcxSVBil49fwMYMLdRxzv/aUvg3WTcnJRD5a7FRElL4KQw7J8G5CES/Y2Kqu
VIb+t1AWh9mOCFg7yPx8OnxbEQj486T6XCZ2eC/H1sjVJOvS9tRex2BQOLLo
xJ+vRT+CUNhrl00t9DLVaPysb1oY9yPw1ZBGqG3fzw+HKoCeSf+lUfscv1pI
vRc/aEsX3LUZDnyreDkg+mspo3kFPpDvv+RBd7RSOjtisoYOsmy1qYmu63bj
KX65hDDWiGpq/5r89Ko35nPgTvPGBXrZwsErW72Y8PSMjC1PhHCUZeHXUcyg
0E7dHdvAO6+jb3jRQhsY0jdGJs3fcmppOnjGbMgxKtejkD7p2WjrRzpYzwH/
PAGKMLdpsjx8xn58Vfomw7cvBs3dGe/6g/u7qx/eS5qpMKNyvlmUFEiCCeNz
wS3bM56yrItNyhnDOlsQiHMQyTcngATZUG8BlqSSsDDwpGfygzmMDoE07ua/
UsE3xSl+ST4V2Rfyh0/krcEnyP6fM00Olsc/WBFivixrYX7XD8JpdsX57LJ/
3RMSoNSQH7dfIZctcumwjAPDZCAECKtr8FDPNWMJvnRSS9sUtDxCj3ZZVl1i
+Fmy+mcMrmkLw7da2y76wXHlDBbYtKRnsDUNtPjXogH6XSRysK+hK5BKMzYu
hO/9VlcEzltA9wYN2fXy/p06cKnuVZgHLjJn/+F0g2VvTDbpG065qj2Z4CkK
+43x5sQEoSGmIBmTngiVKQVpB+Vd7aNHMGQMFGjNkAw0BqzxZ5OEbux3p8Hs
DDdWvDFAO2UfmXiQEyLKe7AQrIJIgfmibMD/Tq0lYFg2oYrOoJi4Em8qZ/i3
/IbbDhE0iOBtxlacOw+bJ13c4iJ8tIbwUH02Obb9PzmFyQr+JHli6fJFjxQ/
FINUBFS98oGdwfiBfMcL5QIm/Eo7hDlrM5s4CQ1JrQqxD6CS2hSbC0UXji+l
q9BCNP/xIf22tUta920xLTpJmd7eu5mEpQAXHgwT4lcFvVq3f/q/0zoHTPkw
Qqs+F9H+SgVOgdUPZnd8aQNSEHW3C2UnpGm0PCse9Bolgv6Y90Km23samGQm
P3+SjP99Y7zHiw+w9M++/pzLkW1pD3o7KzcFmeGDAZsGQPqoQ+BZbAx9sL89
aXgbqPSsqtgclIUT17fBVRx208+YYKnK3MlWLKnmgt5mG3i80dJvQ/3o5iVL
cXh37Bgl45hgF9tCemBxzj1vOaNgWH8nRsbfrUZGOKNTusdwgjGbQrnyG0Sz
z9WZccrUAjlKGk5bH9L/vjxdxrGhY6TLyS2qsALFdD2ft3AkPn+g8aR1g21y
TuSHz5365ZKjYxnwYfzdGeLXNIHGEn3a3ay6sJGfJiTgOOqnb+12++BPwQmd
D/w2Z8V0gC9Ghh2E0oIpTW9I6Psv4rRPYjJDVeNkgt9fCtN8yDBORpLySMdf
K8DeKpRVrOrrOgWoYtHoWAUCt1WOnopOUkcvEKARPG/o41KxrOG93+AlvpUf
GE51ZrVgGAF9XGWR3tjdZ32GDXd2D1Q0nqBGc32GQDKscTrmgICYqA997bN6
MeRtOmEhM5JxNptMBd11OI8pKG98m2iej/UWn9ODTje7vqmdLr4fLawk8zoi
CbVwumuT2vdJ6tqhzJ7yMZDLTEB+1RGH7UW5diFVoooN+XwqUo5FQx3NIOAn
r0hH2OdkvCqqPEQdpFC7RufYwOjr24YxCGdjtjn9r3be9Kh6eewRj72USGVH
HUGkliaFWl0KUjpk+rLDxmhC1rY9IayHmFwquOglDbzoelSkdZWBaGphzeHk
QOJ3uzvYiG8OBDs7j1t7whvdciGUDNjsaLud8KW/H16v7CfbFXZbO3cFAOyL
SyvL1p0UVDR32+SRAXB9Ox17x43k5sGFfsc2AxrmBXl4Kz+TyJ3+sE674zh+
8WbMBDQLeOHQj1MSJ+RRwdWW72q0Gn/ycrAc2Ylz2jn7h2hwKxFkMdNHqOLJ
0jRhTAZ6iTiGOwCQ6FlWSVfVWEW6xMyhaNaADHoz27vIrG+XUYRmCtfBB/0D
EEvDonXDz9MUrvX58dwc1Dg/khankhA+hSmEY79g+CoVIZuSS+OM1A7tvkL1
Z66uobEBWB4iJmu2SnNur/JtQGIb0z9bWoe/ko1hC4Z8z4EbWiqqKIS1PYqD
PFbCZ1kWmHIv04Oy/SUFVVn4Pb9wda4AufdhEnzPRPIGaPwaPdqgfLHX0USE
d74Qlx/wQFBsxfXOOkMrvF9LncU5hAoeBH0al1UX0t6JzMwPI8UQPG8SQqPb
aX/YjUmTH3VLhvurD9UYAegYqZuHFYXo5lCj4MM9D0KFLecz3zSe/wq67LYn
3Jcxo4buXyhRMjhcDwTfx9LMAqJ9y+u9IbDxxmmagSa/3pa/GKlyzGyVSfg8
yMvrNsGv3RaVZPMrXfwcvlkmywHM7J46KrvioExKUHU7we1myCgSnoyZDWrH
8uhBn1LRJkMWMWqxJ+XlyP/zCks7WXA5NjwvpQUaeCaWuqT2Fz0U+S5k6r3n
G7rRKCdmNwFHupMi3COaOOEXWKF0DrxtBuax7aoSpw8x2+LLEA5mJQV3QWb+
AQkV+R0BhfcFrq7rK8INb8QrBJw/rg54UP39Yhvw+DeE9Stu+lzS01KB36kp
Z49O3qsO7G3ZBgVKVcFBnhl9RiWOSNWT/0z1uqxmVGaZgVux9LyQhzmlB5/b
ygWbUwg5XW9gKs2EJ+JG2ejR768FAkCuwFqSKVBXk1rX4COjzoY0xnLb/L7N
JZtWMSAv28KMWh9uS9qcYzNGAAZz/QPR2W/oEwod2T/4kFq2lyoY9MIpevEX
QfWKystIJilpPQvoOkCjksJZkc890wNjWszWy1ncbxgn1dw1p+FYtxBHPkmQ
X26IvMm79lL+TjoAGSjYucRHRsCZHkKqEyxuuE0Zkrsi66E7xHvECH9HyaNn
mpM23GfLwtpJ+xMJVLDhFR3vnfYWjUYkUAiIA+dEdTFnBfYUFxJmaskAlnf0
fqTO0Pne1flcN/mxSNEFcWcSVkaPQCHonk1UR121oAcg8rFa4bax1aH/ShtT
dPLFGobBVRv2KNkMXWKqsAEU4DcdabBVtOipMDbI0h/8p/jTd8pbrziew95K
OD2h62toJNP6Tr9SmFVH5Z7k15povSwhiS894mGyt99plM2kIOK2aYPnCdoz
zE4X6f9hGFrqXHub6EPysXqHdNW3f4Lfp4KLWFYbh0AHx/fjscS/8J2cPV2T
wm9acy1jNUzA34Ph/zfTV/9ZNYTv5a8j9yfxRemH45nsAoEIxP7xgCM8bk3q
DlN8chz69gwy9yLScijxfEUCCGpbuwYnxqMCCbL5CMUNHYc12G/rl9RP5+bh
B6J5QKL8iUxt5Z4RceWRlL8Lu7GyluYepqyWCrDg99bRK4QV7YiNscW0bohW
6N1c4ZpRNPQZu8HlH1KixuhlRf8/cfNxMJb+GE/NmyZ/5XaS5xqVZKcGoyo0
ZB9l155N9j5Kzs6pb3ZWwBEvKGqxcKo+mvtRG0efrLBRsEvDcS3UcqUN72FP
mMUfuSmQ60fxjGoYryF6FR6UK57/ohXd3JmqH8yUfCy6uMLy4ChYxebqiLQx
FX6MY62uHRkES/UbsO1tui0q8CgXG/9NNJoZDunVLYLADiZNPGBtFj2Sh7e4
Aju1tcmwH1qd367+EO5C7nlWAP3NkQ/cYzcSSWh9B3+W2g2AKyaG9b0AuiZ1
rVK9KGGHe4jT8wMfTidTgkhJV4cAcl5EEqvgBNtiJKbkbQ8MdFCcGSjYIPe0
YeX5cUhpEqjFNXA9NkvYDIYfSXa4ISoBYDQWYWEZHEKfz1zaMgeR5gP5stFG
3KudNapnu6jOZ9EEksuy0iVHZKWj/5ASYNqHrldySUyeTZuotmQig2J5X9ZK
V+rnkrPRG/F1irK9VRDYEWglw+YbMT/rNdOgWs2ExCKD1k61g2pOtfvvlC28
ORNIGb29QxpO4KhCl1Y6smczRw99aWqhS7chQaj67AVqEhIfEaIkys1bY7qf
20AfaQcNGrCCiJ660SFh5C6nhwDvzlnaq6I6byYZhzSRpQz5vXL9yWXWxSyQ
M+TPD44JmMtK5swx05gL5TlQ5IHyJstuGWtOcM1dv44zxo05yismR3eCpEFU
yJFj8nSktAzeYnvy99sDXSBlpFB1mpNncxRZ39CRaNY4ctQEImVRZdpb3Kin
4+unzueS8e9PfEx6W+zZWLJyi2/BxL9d/0bcye8GJ/8pIAEwE4hkojOCs9UM
hBj+YHR7O6DwXpLxbxzzxkqwpNXHF7mU+/nzZ4ynRFRv1z3HLG2fWNbmPFgB
KhUS0DjmX2izhtPU5KXxTKPgBjT1R6LducHs1LtiBbocfyIwnuU7QqO3sXBY
+3VK1rYcgZ2e3+HcF32uukkjUoeI50n3v7FlZOk/QOfq74M6yZGxWjeywLxp
SiQq0sCzYhl/OTG2HWtz2W/fUGH3IR+66AKxgzKRChc0tFgQJk4nEMsmIGkJ
IlnhnJ+AkZkpYUfvLuXNT8AlK+I54UjCVUVFaB2FpbgRMFQuMvFZOpvDXsXa
N426EZC0WuxxkAs7mgQN8d9tN2DI8ZhlYB6MjKipfJyRF2iOFLC+9ONlqgrA
jfnUp8iwsADRxYZ6N3+fMRcnhGDN77hTAkMb0o7t04ShV96fQfHUkUzTLLs7
kpshkHmay491fRWIdZtm+kZplqddQpG+HPnWygDvbYD6A/6oyLyuSE2gLWUx
nMtZdoJtMR5XOBhFOxBru5w7Z0Q6T3Af5tLHXn2aXrHpPrVSLSmcuP+pCSlj
36LKwAtttpf2xAbanEdYBqF3cENwHAuJxWLFYuLxEoaKxLM3LY4WCm251LTU
NGaa3vZS66MmXiPjsvOE0ASTNUEm2l8+JfL2uZGdODQqZIZox+xGFJOhHQQP
bsBS0Aik9hSrzkY1n8jG5tzR21F8o60BG4nqo8AM3TJWyl6Yiogekb7u+MF8
vdU1YQ8nUTPICBSFhvQsgVR4N2O3Vd1g8p9zMqFcMVCYxOzJeZb7rYvEqrYE
DGqBIfMCcE8Vbf9zpsedHAa3yuw7q/lobqlIwkZINK9vkbFGJoNQTompK4vk
5Si97tgSrZnAAJdVzZlcnxN30m9wIXz9S0XXvJSeSxAwbnl61HmOtdsPE43F
j9hntgI6hXneddh7oDqSAB5+96gxsTwKFv9E28ddf/fksOrBnh8YXveSTxYQ
VIUQxqzKIkAe5SxtttiYNnHSjfj+WyNOSKcrnOdU8B2a7BjYZx9RfhjNBc90
pWz277tA9qSEyY3Zi8zkkQAAby30sCvZVBQAPdfAXFipn/RqyZ+FwuGgP+z0
SL2nd/03iOlkf07e+Wz0m0aSwmTO97AA7gb0EPGePPPNlY/NfZaEoYsoQN0K
YHc4+8yLDUn1AkNiLNwaFlCa8xKl0PamDC02Vyhws8o7kZyOns6To2K3tiZM
jRpjpL+EDm9zVKYUmtb4fUn++taKrFPsKqacg4o9ZZxd/G8onh+L6XO46iI5
qmyavpjUA1M2Y+R0PXRfRj1VrfXt8N3HV1OVG74V3QA9r9douGcBlukh+uZA
xn4dx48cuQv45DSzZNSgqkZBORwfeBBwOnOPWEHwEFudINNXvJl0eKT4J329
/AhmERDPcjwu3Kwso6NlgPhh3RydBp+ge5Q7ZGXP4MhpxskmhXMvHb/6HoH0
BdUxexIsBKnUc6yTswICSo1OIKL46upTCpxhZpfTy4SneYU0OsZwj50yoeby
48B0LcX4bLlRyoTNLQmq6nx9isoTNSULrW8SlTU+te5cisUlP+ZjhNxIEbEV
UaT8Q7XkO+n1r4pN0MHZ53JWMZICW5km6uV2xKUUwRv/1Fm2kgytTg6ND+Gq
E2GfKCuAY3/alxgwkedjtZaF76KYu653v/fUC+zZ7ucWeKCtCVqb4Kldlu9k
jaYsr2ZXTWnm71fB623VUx1p9VcMrLlSghaYCHsRUkc+RR8psQFqtDgkIoy/
EzKjM+aheeYdwmBJKMy2wpDC/O6b+jm78woYw2KkMCknagJQGmWqPLqOXU45
VJg7gcVT1q0w+tQB9/dtA0iZtRkc9GEQz2UFTWHiyFu4vmi79fFC5t+tOZUC
JnCgobYy+cQJr6gUTYp36WyKG9AABRQEDeTZP4H5zb8Gz5ioV6OtBzPM4PPa
AXZ/wk+KJbspPhpT3X8QWeiCdJo3IuAdaXzAzSnDyNJE9upzpQUjXTN8UnVA
m6Mg+rif2MnJIZOZxI9kWY44sw5F6m2Z7oAUUUZ98r3int8/3hu+J/MFaJTy
Ofks0ttY6VtCdudy5B0uj/rH+g6usUnazKPNgCncUEreAHB906HeHxwnfwhY
Qc50raqR58uYgvO2eaB+QEIEY6q6jw4SmKo0bx/tnCBO05NF551zeO29o7Mw
55ssaB8xZ+DLWn7o+d3zxAMn7dbifRXD+0cg6cua4LFqSz76CW+ZueHc6muD
6PJzXcoWyamsFaJj2N1K4fvwau7Tz/2OEZL+fYDJHHiVVnqj6xUCkOc2zgCt
8NdGvkb8Ag==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG2/dMrjIwvwcH4ORMYpRR5mGUAQyQMiDHj9Mso78y2mZuUq7rX6milMW6FpeIczunWVZivZ15icxvcCESSWfw3U9NNhaConZv+Vyqpd1PT1xjTnr2Ir+Myk46Bwu4LnSOyAJ2TIUV3ceCI2PPzM4cPpIQHqwJk756k6ZrT9hcYg8s41bne4/GH0bNhRfPo5LWDCAwx+d3eE/rIDPgq8TeeV0++bPnTFOb9SiWSUNmuS/uBSSCSqSecy+Mtp9lEKAXhtLsyEG7YmfBf7hveBtLHe6c2JJ49Fp9FJ5p+9v01gY3UAxCoBuZ7YlicZLq5OWp7lSVMiRz6tMLlOh6OqCY63fdhdUwfDgaxNTRJHfLK1uomtDcAu8z520AC+Fie50xnczUNhQoCwagK0DiFfX5WUy6k/uYKzrtacGKsaLA51n9FicewbHi95e6/AyMuxlB/8fXVlSTv+MzwnGgxlVMbPmgScDSKiG/WR9Nhyp8R1cBy8YvdwqSl8hqxN0bIGtkn/zgR/DjTJ2poFwNJS+DXYMGskQblcaJ9zMzhatPjSxs5KHs8WXOAJHxmD+frHv8boCtjgvAlLnDMlEZfnFtRMQHCot0+1KYfgTOg651Sm0D8E+ztjGpXOf/VfRaWh+jPqhTt6gREnPb9FiTy03rFw29xpiH2I3tljr48x/31WeFQhw59o09cH7FD3HcDQ/tMf8nuljXKflDlL2qZRzIH/lhUhSBq3egSlWtJZvpxtwIg5/yHY7dE30KVPHElug8E/AehZUAlLPX7ECYOfcjNv"
`endif