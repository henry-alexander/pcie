// (C) 2001-2024 Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions and other 
// software and tools, and its AMPP partner logic functions, and any output 
// files from any of the foregoing (including device programming or simulation 
// files), and any associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License Subscription 
// Agreement, Intel FPGA IP License Agreement, or other applicable 
// license agreement, including, without limitation, that your use is for the 
// sole purpose of programming logic devices manufactured by Intel and sold by 
// Intel or its authorized distributors.  Please refer to the applicable 
// agreement for further details.


//------------------------------------------------------------------------------
 
  module system_intel_pcie_gts_0_phy_hal_2100_ebn43xi
  #(
        parameter ch_l_xcvr_tx_preloaded_hardware_configs_atom     = "TX_PRELOADED_HARDWARE_CONFIGS_NONE"       ,
        parameter ch_l_xcvr_tx_protocol_hint_atom                  = "TX_PROTOCOL_HINT_DISABLED"                ,
        parameter ch_l_xcvr_tx_datarate_bps_atom                   = 37'b0000000000000000000000000000000000000  ,
        parameter ch_l_xcvr_tx_prbs_gen_en_atom                    = "TX_PRBS_GEN_EN_DISABLE"                   ,
        parameter ch_l_xcvr_tx_prbs_pattern_atom                   = 4'b1001                                    ,
        parameter ch_l_xcvr_tx_bond_size_atom                      = "TX_BOND_SIZE_UNUSED"                      ,
        parameter ch_l_xcvr_tx_user_clk_only_mode_atom             = "TX_USER_CLK_ONLY_MODE_DISABLE"            ,
        parameter ch_l_xcvr_tx_width_atom                          = "TX_WIDTH_DISABLED"                        ,
        parameter ch_l_xcvr_tx_word_clk_hz_atom                    = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_xcvr_tx_dl_enable_atom                      = "TX_DL_ENABLE_DISABLE"                     ,
        parameter ch_l_xcvr_rx_preloaded_hardware_configs_atom     = "RX_PRELOADED_HARDWARE_CONFIGS_NONE"       ,
        parameter ch_l_xcvr_rx_protocol_hint_atom                  = "RX_PROTOCOL_HINT_DISABLED"                ,
        parameter ch_l_xcvr_rx_datarate_bps_atom                   = 37'b0000000000000000000000000000000000000  ,
        parameter ch_l_xcvr_rx_prbs_monitor_en_atom                = "RX_PRBS_MONITOR_EN_DISABLE"               ,
        parameter ch_l_xcvr_rx_prbs_pattern_atom                   = 4'b1001                                    ,   
        parameter ch_l_xcvr_rx_width_atom                          = "RX_WIDTH_DISABLED"                        ,   
        parameter ch_l_xcvr_rx_force_cdr_ltr_atom                  = "FALSE"                                    ,
        parameter ch_l_xcvr_rx_adaptation_mode_atom                = "RX_ADAPTATION_MODE_DISABLED"              ,   
        parameter ch_l_xcvr_rx_word_clk_hz_atom                    = 36'b000000000000000000000000000000000000   ,   
        parameter ch_l_xcvr_rx_dl_enable_atom                      = "RX_DL_ENABLE_DISABLE"                     ,
        parameter ch_l_rx_postdiv_clk_en_atom                      = "RX_POSTDIV_CLK_EN_DISABLE"                ,
        parameter ch_l_rx_postdiv_clk_divider_atom                 = 8'b00000001                                ,
        parameter ch_l_tx_postdiv_clk_divider_atom                 = 8'b00000001                                ,
        parameter ch_l_tx_pll_refclk_select_atom                   = "TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0"      ,
        parameter ch_l_loopback_mode_atom                          = "LOOPBACK_MODE_DISABLED"                   ,
        parameter ch_flux_l_flux_mode_atom                         = "FLUX_MODE_DISABLED"                       ,
        parameter ch_flux_l_rx_protocol_hint_atom                  = "RX_PROTOCOL_HINT_DISABLED"                ,
        parameter ch_flux_l_tx_dl_enable_atom                      = "TX_DL_ENABLE_ENABLE"                      ,   
        parameter ch_flux_l_rx_dl_enable_atom                      = "RX_DL_ENABLE_ENABLE"                      ,
        parameter ch_xcvrif_l_tx_dl_enable_atom                    = "TX_DL_ENABLE_ENABLE"                      ,
        parameter ch_xcvrif_l_rx_dl_enable_atom                    = "RX_DL_ENABLE_ENABLE"                      ,
        parameter ch_xcvrif_l_loopback_mode_atom                   = "LOOPBACK_MODE_DISABLE"                    ,
        parameter ch_xcvrif_l_tx_fifo_mode_atom                    = "TX_FIFO_MODE_DISABLED"                    ,
        parameter ch_xcvrif_l_rx_fifo_mode_atom                    = "RX_FIFO_MODE_DISABLED"                    ,
        parameter ch_flux_l_tx_bond_size_atom                      = "TX_BOND_SIZE_UNUSED"                      ,
        parameter ch_xcvrif_l_tx_bond_size_atom                    = "TX_BOND_SIZE_UNUSED"                      ,
        parameter ch_xcvrif_l_rx_bond_size_atom                    = "RX_BOND_SIZE_UNUSED"                      ,
        parameter ch_l_xcvr_tx_en_atom                             = "FALSE"                                    ,           
        parameter ch_l_xcvr_rx_en_atom                             = "FALSE"                                    ,
        parameter ch_l_duplex_mode_atom                            = "DUPLEX_MODE_DUPLEX"                       ,
        parameter ch_xcvrif_l_tx_en_atom                           = "FALSE"                                    ,
        parameter ch_xcvrif_l_rx_en_atom                           = "FALSE"                                    ,
        parameter ch_xcvrif_l_duplex_mode_atom                     = "DUPLEX_MODE_DUPLEX"                       ,
        parameter ch_flux_l_rx_fec_type_used_atom                  = "RX_FEC_TYPE_USED_NONE"                    ,
        parameter ch_l_sim_mode_atom                               = "SIM_MODE_ENABLE"                          ,
        parameter ch_flux_l_rx_sim_mode_atom                       = "RX_SIM_MODE_ENABLE"                       ,
        parameter ch_flux_l_tx_sim_mode_atom                       = "TX_SIM_MODE_ENABLE"                       ,
        parameter ch_flux_l_dr_enabled_atom                        = "DR_ENABLED_DR_ENABLED"                    ,
        parameter ch_xcvrif_l_sup_mode_atom                        = "SUP_MODE_USER_MODE"                       ,
        parameter ch_xcvrif_l_sim_mode_atom                        = "SIM_MODE_DISABLE"                         ,
        parameter ch_xcvrif_l_dr_enabled_atom                      = "DR_ENABLED_DR_ENABLED"                    ,
        parameter ch_l_xcvr_tx_spread_spectrum_en_atom             = "TX_SPREAD_SPECTRUM_EN_ENABLE"             ,
        parameter ch_l_xcvr_cdr_f_ref_hz_atom                      = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_xcvr_cdr_f_vco_hz_atom                      = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_xcvr_cdr_f_out_hz_atom                      = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_xcvr_cdr_f_pfd_hz_atom                      = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_cdr_l_counter_atom                          = 6'b000001                                  ,
        parameter ch_l_cdr_m_counter_atom                          = 9'b000000001                               ,
        parameter ch_l_cdr_n_counter_atom                          = 6'b000001                                  ,
        parameter ch_l_tx_pll_f_ref_hz_atom                        = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_pll_f_out_hz_atom                        = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_pll_f_pfd_hz_atom                        = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_pll_f_vco_hz_atom                        = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_pll_k_counter_atom                       = 22'b0000000000000000000000                 ,
        parameter ch_l_tx_pll_l_counter_atom                       = 6'b000001                                  ,
        parameter ch_l_tx_pll_m_counter_atom                       = 9'b000000001                               ,
        parameter ch_l_tx_pll_n_counter_atom                       = 6'b000001                                  ,
        parameter ch_l_tx_pll_fb_counter_atom                      = 2'b10                                      ,
        parameter ch_l_tx_pll_postdiv_sel_atom                     = "TX_PLL_POSTDIV_SEL_SYNTH_FAST"            ,
        parameter ch_l_tx_synthdiv_out_hz_atom                     = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_synthdiv_out_divider_atom                = 8'b00000001                                ,
        parameter ch_l_tx_postdiv_cdr_refclk_hz_atom               = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_postdiv_cdr_refclk_divider_atom          = 8'b00000001                                ,
        parameter ch_l_rx_postdiv_clk_hz_atom                      = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_rx_postdiv_clk_fractional_en_atom           = "RX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE"     ,
        parameter ch_l_cdr_refclk_select_atom                      = "CDR_REFCLK_SELECT_GLOBAL_REFCLK0"         ,
        parameter ch_l_tx_postdiv_clk_hz_atom                      = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_tx_postdiv_clk_fractional_en_atom           = "TX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE"     ,
        parameter ch_flux_l_lc_postdiv_sel_atom                    = "LC_POSTDIV_SEL_SYNTH_FAST"                ,
        parameter ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom      = "TX_USER1_CLK_MUX_DYNAMIC_SEL_UNUSED"      ,
        parameter ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom      = "TX_USER2_CLK_MUX_DYNAMIC_SEL_UNUSED"      ,
        parameter ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom      = "RX_USER1_CLK_MUX_DYNAMIC_SEL_UNUSED"      ,
        parameter ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom      = "RX_USER2_CLK_MUX_DYNAMIC_SEL_UNUSED"      ,
        parameter ch_xcvrif_l_tx_gb_width_atom                     = "TX_GB_WIDTH_DISABLED"                     ,
        parameter ch_xcvrif_l_rx_gb_width_atom                     = "RX_GB_WIDTH_DISABLED"                     ,
        parameter ch_xcvrif_l_tx_dynamic_mux_atom                  = "TX_DYNAMIC_MUX_UNUSED"                    ,
        parameter ch_xcvrif_l_tx_word_clk_dynamic_mux_atom         = "TX_WORD_CLK_DYNAMIC_MUX_UNUSED"           ,
        parameter ch_xcvrif_l_rx_word_clk_dynamic_mux_atom         = "RX_WORD_CLK_DYNAMIC_MUX_RXWORD_CLK"       ,
        parameter ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom       = "TX_FIFO_RD_EN_DYNAMIC_MUX_UNUSED"         ,
        parameter ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom       = "RX_FIFO_RD_EN_DYNAMIC_MUX_UNUSED"         ,
        parameter ch_xcvrif_l_tx_rst_dynamic_mux_atom              = "TX_RST_DYNAMIC_MUX_UNUSED"                ,
        parameter ch_l_clk_debug_select_0_enable_atom              = "CLK_DEBUG_SELECT_0_ENABLE_DISABLE"        ,
        parameter ch_l_clk_debug_select_0_setting_atom             = "CLK_DEBUG_SELECT_0_SETTING_DISABLED"      ,
        parameter ch_l_clk_debug_select_1_enable_atom              = "CLK_DEBUG_SELECT_1_ENABLE_DISABLE"        ,
        parameter ch_l_clk_debug_select_1_setting_atom             = "CLK_DEBUG_SELECT_1_SETTING_DISABLED"      ,
        parameter ch_l_xcvr_tx_eq_main_tap_atom                    = 6'b000000                                  ,
        parameter ch_l_xcvr_tx_eq_post_tap_1_atom                  = 5'b00000                                   ,
        parameter ch_l_xcvr_tx_eq_pre_tap_1_atom                   = 5'b00000                                   ,
        parameter ch_l_xcvr_tx_eq_pre_tap_2_atom                   = 3'b000                                     ,
        parameter ch_l_tx_pll_feed_forward_gain_atom               = 8'b00000001                                ,
        parameter ch_l_xcvr_rx_termination_mode_atom               = "RX_TERMINATION_MODE_HIGH_Z"               ,
        parameter ch_l_xcvr_rx_onchip_termination_setting_atom     = "RX_ONCHIP_TERMINATION_SETTING_R_1"        ,
        parameter ch_l_xcvr_rx_eq_vga_gain_atom                    = 7'b0000000                                 ,
        parameter ch_l_xcvr_x_eq_hf_boost_atom                     = 6'b000000                                  ,
        parameter ch_l_xcvr_rx_eq_dfe_tap_1_atom                   = 6'b000000                                  ,
        parameter ch_l_xcvr_rx_external_couple_type_atom           = "RX_EXTERNAL_COUPLE_TYPE_AC"               ,
        parameter ch_l_tx_pll_bw_sel_atom                          = "TX_PLL_BW_SEL_LOW"                        ,
        parameter ch_l_xcvr_tx_bonding_category_atom               = "TX_BONDING_CATEGORY_UNUSED"               ,
        parameter ch_l_xcvr_tx_master_pll_mode_atom                = "TX_MASTER_PLL_MODE_DISABLED"              ,
        parameter ch_l_xcvr_rx_cdrdivout_en_atom                   = "RX_CDRDIVOUT_EN_DISABLE"                  ,
        parameter ch_xcvrif_l_tx_bonding_mode_atom                 = "TX_BONDING_MODE_UNUSED"                   ,
        parameter ch_xcvrif_l_rx_bonding_mode_atom                 = "RX_BONDING_MODE_UNUSED"                   ,
        parameter ch_l_speed_grade_atom                            = "SPEED_GRADE_DASH_1"                       ,
        parameter ch_flux_l_sequencer_reg_en_atom                  = "SEQUENCER_REG_EN_DISABLE"                 ,
        parameter ch_usb_mode_atom                                 = "USB_MODE_DISABLED"                        ,
        parameter ch_pcie_mode_atom                                = "PCIE_MODE_DISABLED"                       ,
        parameter ch_l_ick_tx_word_clk_hz_atom                     = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_pcs_ref_clk_hz_atom                         = 36'b000000000000000000000000000000000000   ,
        parameter ch_l_lane_common_ref_clk_hz_atom                 = 36'b000000000000000000000000000000000000   ,
        parameter ch_rx_invert_pin_atom                            = "RX_INVERT_PIN_DISABLE"                    ,
        parameter ch_tx_invert_pin_atom                            = "TX_INVERT_PIN_DISABLE"                    ,
        parameter ch_rx_dl_rx_lat_bit_for_async_atom               = 18'b000000000000000000                     ,
        parameter ch_rx_dl_rxbit_cntr_pma_atom                     = "RX_DL_RXBIT_CNTR_PMA_ENABLE"              ,
        parameter ch_rx_dl_rxbit_rollover_atom                     = 18'b000000000000000000                     ,
        parameter ch_eth_rx_clk_hz_atom                            = 36'b000000000000000000000000000000000000   ,
        parameter ch_eth_tx_clk_hz_atom                            = 36'b000000000000000000000000000000000000   ,
        parameter ch_clkrx_refclk_cssm_fw_control_atom                = "CLKRX_REFCLK_CSSM_FW_CONTROL_ENABLE"               ,
        parameter ch_clkrx_refclk_sector_specifies_refclk_ready_atom  = "CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_ENABLE" ,
        parameter ch_local_refclk_cssm_fw_control_atom                = "LOCAL_REFCLK_CSSM_FW_CONTROL_ENABLE"               ,
        parameter ch_local_refclk_sector_specifies_refclk_ready_atom  = "LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_ENABLE" ,
        parameter ch_flux_l_stmux_rx_demux_sel                     = "SEL_XCVRIF"                               ,
        parameter ch_flux_l_stmux_rx_rxword_clk_demux_sel          = "SEL_ETH_RXWORD_CLK"                       ,
        parameter ch_flux_l_stmux_tx_txword_clk_demux_sel          = "SEL_ETH_TXWORD_CLK"                       ,
        parameter ch_flux_l_stmux_tx_mux_sel                       = "SEL_XCVRIF"                               ,
        parameter ch_flux_l_stmux_tx_txword_clk_mux_sel            = "SEL_XCVR_TXWORD_CLK"                      ,
        parameter ch_xcvrif_rx_ch_clk_static_mux                   = "SEL_SYS_CLK"                              ,
        parameter ch_xcvrif_tx_ch_clk_static_mux                   = "SEL_SYS_CLK"                           
        
)
(
        output          oflux_xoa_tx_n_l0_ux,
        output          oflux_xoa_tx_p_l0_ux,
        input           iflux_xia_rx_n_l0_ux,
        input           iflux_xia_rx_p_l0_ux,
        input   [79:0]  i_ss_async_pldif,        
        output  [49:0]  o_ss_async_pldif,        
        input   [79:0]  i_ss_async_pldif_pcie_mux,
        input   [19:0]  i_lavmm_addr,                       
        input   [3:0]   i_lavmm_be,
        input           i_lavmm_clk,
        input           i_lavmm_read,
        input           i_lavmm_rstn,
        input   [31:0]  i_lavmm_wdata,
        input           i_lavmm_write,
        output  [31:0]  o_lavmm_rdata,
        output          o_lavmm_rdata_valid,
        output          o_lavmm_waitreq,
        input           i_ft_rx_sclk_sync_ch,
        input           i_ft_tx_sclk_sync_ch,
        output          o_ft_rx_async_pulse_ch,
        output          o_ft_tx_async_pulse_ch,
        output          o_rxcdrlock2dataa,
        input           i_rst_ux_rx_sfrz,
        output          o_rst_flux0_cpi_cmn_busy,
        output          o_rst_oflux_rx_srds_rdy,
        output          o_rst_ux_all_synthlockstatus,
        output          o_rst_ux_rxcdrlockstatus,
        output          o_ux_tx_ch_ptr_smpl,                                                    //Check, Raised to PFE
        input           i_ick_sclk_tx,
        input           i_ick_sclk_rx,
        input           i_rst_pld_ux_tx_pma_rst_n,
        input           i_rst_pld_ux_rx_pma_rst_n,
        output  [31:0]  o_ch_lavmm_xcvrif_rdata,
        output          o_ch_lavmm_xcvrif_rdata_valid,
        output          o_ch_lavmm_xcvrif_waitreq,
        input   [19:0]  i_ch_lavmm_xcvrif_addr,
        input   [3:0]   i_ch_lavmm_xcvrif_be,
        input           i_ch_lavmm_xcvrif_clk,
        input           i_ch_lavmm_xcvrif_read,
        input           i_ch_lavmm_xcvrif_rstn,
        input   [31:0]  i_ch_lavmm_xcvrif_wdata,
        input           i_ch_lavmm_xcvrif_write,
//        input           i_pld_rx_lat_sclk_ch,             //In r10 Removed
//        input           i_pld_tx_lat_sclk_ch,             //In r10 Removed
        output          o_rx_latency_pulse,
        output          o_tx_latency_pulse,
        input   [42:0]  i_xcvrif_tx_mux_data,                        
        output  [42:0]  o_rx_data,
        output  [1:0]   o_tx_source_sel,  
        input   [6:0]   i_ch_eth_xcvrif_tx_async,
        input           i_ch_eth_xcvrif_tx_direct,
        output  [13:0]  o_ch_eth_xcvrif_rx_async,
        output          o_ch_eth_xcvrif_rx_direct,
        input           i_rstxcvrif_xcvrif_signal_ok,
        input           i_rstxcvrif_rx_xcvrif_sfrz_n,
        input           i_rstxcvrif_xcvrif_rx_rst_n,
        input           i_rstxcvrif_tx_xcvrif_sfrz_n,
        input           i_rstxcvrif_xcvrif_tx_rst_n,
        output          o_pma_rx_sf,
        output  [2:0]   o_rx_fifo_en_sel,
        output  [2:0]   o_tx_rst_source_sel,
        input           i_ch_xcvrif_rx_fifo_rd_en,
        output          o_ch_xcvrif_rx_fifo_rd_en,
        input           i_ch_xcvrif_tx_fifo_rd_en,
        output          o_ch_xcvrif_tx_fifo_rd_en,
//        input           i_xcvr_rx_ch_clk,                 In r10 Removed
//        input           i_xcvr_tx_ch_clk,                 In r10 Removed
        output  [1:0]   o_ux_rxuser1_sel,
        output  [1:0]   o_ux_rxuser2_sel,
        output  [1:0]   o_ux_txuser1_sel,
        output  [1:0]   o_ux_txuser2_sel,
        output          o_pcs_rxpostdiv,
        output          o_pcs_rxword,
        output          o_ux_txlc_clk,
        output          o_ock_pcs_txword,
        output  [2:0]   o_tx_xcvr_wordclk_sel,
        output  [1:0]   o_rx_xcvr_wordclk_sel,                                //NA in ch4_phy Sujoy RTL
        output          o_eth_rx_ch_clk,                                                   
        input           i_eth_rx_ch_clk,
//        input           i_eth_tx_ch_clk,                                                    //NA in ch4_phy Sujoy RTL
        input  [767:0]  uxwrap_bus_in  ,                 
        output [703:0]  uxwrap_bus_out ,        
        output [19:0]   o_lavmm_addr,
        output [3:0]    o_lavmm_be,
        output          o_lavmm_clk,
        output          o_lavmm_read,
        output          o_lavmm_rstn,
        output [31:0]   o_lavmm_wdata,
        output          o_lavmm_write,   
        input  [31:0]   i_lavmm_rdata, 
        input           i_lavmm_rdata_valid,
        input           i_lavmm_waitreq,    
        output          o_sclk_return_sel_rx,
        output          o_sclk_return_sel_tx,      
        output          o_ick_sclk_rx,           
        input   [4:0]   i_sync_common_control,          
        output          o_ft_rx_sclk_sync_ch,       
        output          o_ft_tx_sclk_sync_ch,       
        output          o_rst_ux_rx_pma_rst_n,      
        output          o_rst_ux_tx_pma_rst_n,       
        output          o_ick_pcs_txword,                   
        output          o_tx_dl_ch_bit,                     
        input           i_dat_pcs_measlatbit,               
        input           i_ft_rx_async_pulse_ch,
        input           i_ft_tx_async_pulse_ch,             
        input           i_rx_dl_ch_bit,                 
        input   [1:0]   i_ux_rxuser1_sel,
        input   [1:0]   i_ux_rxuser2_sel,                   
        input   [1:0]   i_ux_txuser1_sel,
        input   [1:0]   i_ux_txuser2_sel,                   
        output          o_octl_pcs_txstatus_a,              
        input           i_ictl_pcs_txenable_a,      
        input   [124:0] i_sync_cfg_data,                
        input   [249:0] i_sync_interface_control,         
        output  [79:0]  o_tx_data,                          
        input   [79:0]  i_rx_data,                      
        output  [319:0] o_sm_flux_ingress,              
        input   [256:0] i_sm_flux_egress,                       
        input           i_flux_cpi_int,                     
        input           i_flux_int,                     
        input           i_oflux_octl_pcs_txptr_smpl_lane,   
        output          o_ick_sclk_tx,                      
        input           i_flux_srds_rdy,                    
        input           i_pcs_rxword,                           
        input           i_pcs_rxpostdiv,                    
        input           i_ock_pcs_txword,            
        output          o_dat_pcs_measlatrndtripbit,            
//        input           i_dpma_refclk,            //Connected this from cnoc atom in phy_hal_coreip.sv
        output          o_ock_pcs_cdrfbclk,            
        output          o_ock_pcs_ref   ,
        output [39:0]   o_pcie_pcs,
        input [39:0]    i_pcie_pcs,
//New signals Added after r9
        input           i_sel_rxword_clk,
        input           i_xcvr_txword_clk,
        output          o_pcie_rxword_clk,
        output          o_eth_rxword_clk ,
        output          o_pcie_txword_clk,
        output          o_eth_txword_clk,
//New signals Added after r10   
        output           o_eth_tx_ch_clk,
//New Signals Added after r11       
//        input [5:0] ioack_ref_left_n_ux_bidir_in,
        input [5:0] ioack_ref_left_p_ux_bidir_in,
//        input ioack_hsref_left_n_ux_bidir_in,
        input ioack_hsref_left_p_ux_bidir_in,
//New Signals Added after r12
        input ioack_cdrdiv_left_ux_bidir_in,
        input ioack_synthdiv1_left_ux_bidir_in,
        input ioack_synthdiv2_left_ux_bidir_in,
        output ioack_cdrdiv_left_ux_bidir_out,
        output ioack_synthdiv1_left_ux_bidir_out,
        output ioack_synthdiv2_left_ux_bidir_out,

//KAHUAT_EDIT
        output [13:0] o_rxeq_best_eye_vala,
        output        o_rxeq_donea,
        output        o_rxmargin_nacka,
        output        o_rxmargin_statusa,
        output        o_rxsignaldetect_lfpsa,
        output        o_rxsignaldetecta,
        output [1:0]  o_rxmargin_status_gray,
        output        o_synthlcfast_postdiv,
        output        o_synthlcmed_postdiv,
        output        o_synthlcslow_postdiv,
        output        o_txdetectrx_acka,
        output        o_txdetectrx_statct,
        input         i_pcs_pipe_rstn,
        input         i_ux_ock_pma_clk,
        input         i_lfps_ennt,
        input  [1:0]  i_pcie_l1ctrla,
        input         i_pma_cmn_ctrl,
        input         i_pma_ctrl,
        input         i_pcie_pcs_rx_rst,
        input         i_pcie_pcs_tx_rst,
        input         i_rxeiosdetectstata,
        input  [2:0]  i_rxeq_precal_code_selnt,
        input         i_rxeq_starta,
        input         i_rxeq_static_ena,
        input         i_rxmargin_direction_nt,
        input         i_rxmargin_mode_nt,
        input         i_rxmargin_offset_change_a,     
        input  [6:0]  i_rxmargin_offset_nt,
        input         i_rxmargin_start_a,
        input  [2:0]  i_rxpstate,
        input  [3:0]  i_rxrate,
        input         i_rxterm_hiz_ena,
        input  [2:0]  i_rxwidth,
        input         i_tstbus_lane,
        input         i_txbeacona,
        input  [2:0]  i_txclkdivrate,
        input         i_txdetectrx_reqa,
        input  [5:0]  i_txdrv_levn,
        input  [4:0]  i_txdrv_levnm1,
        input  [2:0]  i_txdrv_levnm2,
        input  [4:0]  i_txdrv_levnp1,
        input  [3:0]  i_txdrv_slew,
        input  [3:0]  i_txelecidle,
        input  [2:0]  i_txpstate,
        input  [3:0]  i_txrate,
        input  [2:0]  i_txwidth,

        output o_rxstatusa,     //As per Kumaran Suggestion Connected this port to PLDIF i_ss_rst_ux_octl_pcs_rxstatus
        output o_txstatusa,      //As per Kumaran Suggestion Connected this port to PLDIF i_ss_rst_ux_octl_pcs_txstatus
        input  i_quartus_flux_s_to_ingress, //R24 Integration
        input  i_rstxcvrif_xcvrif_tx_rd_rst_n,
        input  i_rstxcvrif_xcvrif_tx_wr_rst_n,
        output o_tx_rst_rd_sync_rst_n,
        output o_tx_rst_wr_sync_rst_n       
);




  phy_hal_coreip
  # (
        .ch_l_xcvr_tx_preloaded_hardware_configs_atom           (ch_l_xcvr_tx_preloaded_hardware_configs_atom  ),
        .ch_l_xcvr_tx_protocol_hint_atom                        (ch_l_xcvr_tx_protocol_hint_atom               ),
        .ch_l_xcvr_tx_datarate_bps_atom                         (ch_l_xcvr_tx_datarate_bps_atom                ),
        .ch_l_xcvr_tx_prbs_gen_en_atom                          (ch_l_xcvr_tx_prbs_gen_en_atom                 ),
        .ch_l_xcvr_tx_prbs_pattern_atom                         (ch_l_xcvr_tx_prbs_pattern_atom                ),
        .ch_l_xcvr_tx_bond_size_atom                            (ch_l_xcvr_tx_bond_size_atom                   ),
        .ch_l_xcvr_tx_user_clk_only_mode_atom                   (ch_l_xcvr_tx_user_clk_only_mode_atom          ),
        .ch_l_xcvr_tx_width_atom                                (ch_l_xcvr_tx_width_atom                       ),
        .ch_l_xcvr_tx_word_clk_hz_atom                          (ch_l_xcvr_tx_word_clk_hz_atom                 ),
        .ch_l_xcvr_tx_dl_enable_atom                            (ch_l_xcvr_tx_dl_enable_atom                   ),
        .ch_l_xcvr_rx_preloaded_hardware_configs_atom           (ch_l_xcvr_rx_preloaded_hardware_configs_atom  ),
        .ch_l_xcvr_rx_protocol_hint_atom                        (ch_l_xcvr_rx_protocol_hint_atom               ),
        .ch_l_xcvr_rx_datarate_bps_atom                         (ch_l_xcvr_rx_datarate_bps_atom                ),    
        .ch_l_xcvr_rx_prbs_monitor_en_atom                      (ch_l_xcvr_rx_prbs_monitor_en_atom             ),
        .ch_l_xcvr_rx_prbs_pattern_atom                         (ch_l_xcvr_rx_prbs_pattern_atom                ),
        .ch_l_xcvr_rx_width_atom                                (ch_l_xcvr_rx_width_atom                       ),
        .ch_l_xcvr_rx_force_cdr_ltr_atom                        (ch_l_xcvr_rx_force_cdr_ltr_atom               ),
        .ch_l_xcvr_rx_adaptation_mode_atom                      (ch_l_xcvr_rx_adaptation_mode_atom             ),
        .ch_l_xcvr_rx_word_clk_hz_atom                          (ch_l_xcvr_rx_word_clk_hz_atom                 ),
        .ch_l_xcvr_rx_dl_enable_atom                            (ch_l_xcvr_rx_dl_enable_atom                   ),
        .ch_l_xcvr_cdr_f_ref_hz_atom                            (ch_l_xcvr_cdr_f_ref_hz_atom                   ),
        .ch_l_xcvr_cdr_f_vco_hz_atom                            (ch_l_xcvr_cdr_f_vco_hz_atom                   ),
        .ch_l_rx_postdiv_clk_en_atom                            (ch_l_rx_postdiv_clk_en_atom                   ),
        .ch_l_rx_postdiv_clk_divider_atom                       (ch_l_rx_postdiv_clk_divider_atom              ),
        .ch_l_tx_pll_f_ref_hz_atom                              (ch_l_tx_pll_f_ref_hz_atom                     ),
        .ch_l_tx_pll_f_out_hz_atom                              (ch_l_tx_pll_f_out_hz_atom                     ),
        .ch_l_tx_postdiv_clk_divider_atom                       (ch_l_tx_postdiv_clk_divider_atom              ),
        .ch_l_tx_pll_refclk_select_atom                         (ch_l_tx_pll_refclk_select_atom                ),
        .ch_l_loopback_mode_atom                                (ch_l_loopback_mode_atom                       ),
        .ch_flux_l_flux_mode_atom                               (ch_flux_l_flux_mode_atom                      ),
        .ch_flux_l_rx_protocol_hint_atom                        (ch_flux_l_rx_protocol_hint_atom               ),
        .ch_flux_l_tx_dl_enable_atom                            (ch_flux_l_tx_dl_enable_atom                   ),
        .ch_flux_l_rx_dl_enable_atom                            (ch_flux_l_rx_dl_enable_atom                   ),
        .ch_xcvrif_l_tx_dl_enable_atom                          (ch_xcvrif_l_tx_dl_enable_atom                 ),
        .ch_xcvrif_l_rx_dl_enable_atom                          (ch_xcvrif_l_rx_dl_enable_atom                 ),
        .ch_xcvrif_l_loopback_mode_atom                         (ch_xcvrif_l_loopback_mode_atom                ),
        .ch_xcvrif_l_tx_fifo_mode_atom                          (ch_xcvrif_l_tx_fifo_mode_atom                 ),
        .ch_xcvrif_l_rx_fifo_mode_atom                          (ch_xcvrif_l_rx_fifo_mode_atom                 ),
        .ch_xcvrif_l_tx_bond_size_atom                          (ch_xcvrif_l_tx_bond_size_atom                 ),
        .ch_flux_l_tx_bond_size_atom                            (ch_flux_l_tx_bond_size_atom                   ),
        .ch_xcvrif_l_rx_bond_size_atom                          (ch_xcvrif_l_rx_bond_size_atom                 ),
        .ch_l_xcvr_tx_en_atom                                   (ch_l_xcvr_tx_en_atom                          ),
        .ch_l_xcvr_rx_en_atom                                   (ch_l_xcvr_rx_en_atom                          ),
        .ch_l_duplex_mode_atom                                  (ch_l_duplex_mode_atom                         ),
        .ch_xcvrif_l_tx_en_atom                                 (ch_xcvrif_l_tx_en_atom                        ),
        .ch_xcvrif_l_rx_en_atom                                 (ch_xcvrif_l_rx_en_atom                        ),
        .ch_xcvrif_l_duplex_mode_atom                           (ch_xcvrif_l_duplex_mode_atom                  ),
        .ch_flux_l_rx_fec_type_used_atom                        (ch_flux_l_rx_fec_type_used_atom               ),
        .ch_l_sim_mode_atom                                     (ch_l_sim_mode_atom                            ),
        .ch_flux_l_rx_sim_mode_atom                             (ch_flux_l_rx_sim_mode_atom                    ),
        .ch_flux_l_tx_sim_mode_atom                             (ch_flux_l_tx_sim_mode_atom                    ),
        .ch_flux_l_dr_enabled_atom                              (ch_flux_l_dr_enabled_atom                     ),
        .ch_xcvrif_l_sup_mode_atom                              (ch_xcvrif_l_sup_mode_atom                     ),
        .ch_xcvrif_l_sim_mode_atom                              (ch_xcvrif_l_sim_mode_atom                     ),
        .ch_xcvrif_l_dr_enabled_atom                            (ch_xcvrif_l_dr_enabled_atom                   ),
        .ch_l_xcvr_tx_spread_spectrum_en_atom                   (ch_l_xcvr_tx_spread_spectrum_en_atom          ),
        .ch_l_xcvr_cdr_f_out_hz_atom                            (ch_l_xcvr_cdr_f_out_hz_atom                   ),
        .ch_l_xcvr_cdr_f_pfd_hz_atom                            (ch_l_xcvr_cdr_f_pfd_hz_atom                   ),
        .ch_l_cdr_l_counter_atom                                (ch_l_cdr_l_counter_atom                       ),
        .ch_l_cdr_m_counter_atom                                (ch_l_cdr_m_counter_atom                       ),
        .ch_l_cdr_n_counter_atom                                (ch_l_cdr_n_counter_atom                       ),
        .ch_l_tx_pll_f_pfd_hz_atom                              (ch_l_tx_pll_f_pfd_hz_atom                     ),
        .ch_l_tx_pll_f_vco_hz_atom                              (ch_l_tx_pll_f_vco_hz_atom                     ),
        .ch_l_tx_pll_k_counter_atom                             (ch_l_tx_pll_k_counter_atom                    ),
        .ch_l_tx_pll_l_counter_atom                             (ch_l_tx_pll_l_counter_atom                    ),
        .ch_l_tx_pll_m_counter_atom                             (ch_l_tx_pll_m_counter_atom                    ),
        .ch_l_tx_pll_n_counter_atom                             (ch_l_tx_pll_n_counter_atom                    ),
        .ch_l_tx_pll_fb_counter_atom                            (ch_l_tx_pll_fb_counter_atom                   ),
        .ch_l_tx_pll_postdiv_sel_atom                           (ch_l_tx_pll_postdiv_sel_atom                  ),
        .ch_l_tx_synthdiv_out_hz_atom                           (ch_l_tx_synthdiv_out_hz_atom                  ),
        .ch_l_tx_synthdiv_out_divider_atom                      (ch_l_tx_synthdiv_out_divider_atom             ),
        .ch_l_tx_postdiv_cdr_refclk_hz_atom                     (ch_l_tx_postdiv_cdr_refclk_hz_atom            ),
        .ch_l_tx_postdiv_cdr_refclk_divider_atom                (ch_l_tx_postdiv_cdr_refclk_divider_atom       ),
        .ch_l_rx_postdiv_clk_hz_atom                            (ch_l_rx_postdiv_clk_hz_atom                   ),
        .ch_l_rx_postdiv_clk_fractional_en_atom                 (ch_l_rx_postdiv_clk_fractional_en_atom        ),
        .ch_l_cdr_refclk_select_atom                            (ch_l_cdr_refclk_select_atom                   ),
        .ch_l_tx_postdiv_clk_hz_atom                            (ch_l_tx_postdiv_clk_hz_atom                   ),
        .ch_l_tx_postdiv_clk_fractional_en_atom                 (ch_l_tx_postdiv_clk_fractional_en_atom        ),
        .ch_flux_l_lc_postdiv_sel_atom                          (ch_flux_l_lc_postdiv_sel_atom                 ),
        .ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom            (ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom   ),
        .ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom            (ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom   ),
        .ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom            (ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom   ),
        .ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom            (ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom   ),
        .ch_xcvrif_l_tx_gb_width_atom                           (ch_xcvrif_l_tx_gb_width_atom                  ),
        .ch_xcvrif_l_rx_gb_width_atom                           (ch_xcvrif_l_rx_gb_width_atom                  ),
        .ch_xcvrif_l_tx_dynamic_mux_atom                        (ch_xcvrif_l_tx_dynamic_mux_atom               ),
        .ch_xcvrif_l_tx_word_clk_dynamic_mux_atom               (ch_xcvrif_l_tx_word_clk_dynamic_mux_atom      ),
        .ch_xcvrif_l_rx_word_clk_dynamic_mux_atom               (ch_xcvrif_l_rx_word_clk_dynamic_mux_atom      ),
        .ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom             (ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom    ),
        .ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom             (ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom    ),
        .ch_xcvrif_l_tx_rst_dynamic_mux_atom                    (ch_xcvrif_l_tx_rst_dynamic_mux_atom           ),
        .ch_l_clk_debug_select_0_enable_atom                    (ch_l_clk_debug_select_0_enable_atom           ),
        .ch_l_clk_debug_select_0_setting_atom                   (ch_l_clk_debug_select_0_setting_atom          ),
        .ch_l_clk_debug_select_1_enable_atom                    (ch_l_clk_debug_select_1_enable_atom           ),
        .ch_l_clk_debug_select_1_setting_atom                   (ch_l_clk_debug_select_1_setting_atom          ),
        .ch_l_xcvr_tx_eq_main_tap_atom                          (ch_l_xcvr_tx_eq_main_tap_atom                 ),
        .ch_l_xcvr_tx_eq_post_tap_1_atom                        (ch_l_xcvr_tx_eq_post_tap_1_atom               ),
        .ch_l_xcvr_tx_eq_pre_tap_1_atom                         (ch_l_xcvr_tx_eq_pre_tap_1_atom                ),
        .ch_l_xcvr_tx_eq_pre_tap_2_atom                         (ch_l_xcvr_tx_eq_pre_tap_2_atom                ),
        .ch_l_tx_pll_feed_forward_gain_atom                     (ch_l_tx_pll_feed_forward_gain_atom            ),
        .ch_l_xcvr_rx_termination_mode_atom                     (ch_l_xcvr_rx_termination_mode_atom            ),
        .ch_l_xcvr_rx_onchip_termination_setting_atom           (ch_l_xcvr_rx_onchip_termination_setting_atom  ),
        .ch_l_xcvr_rx_eq_vga_gain_atom                          (ch_l_xcvr_rx_eq_vga_gain_atom                 ),
        .ch_l_xcvr_x_eq_hf_boost_atom                           (ch_l_xcvr_x_eq_hf_boost_atom                  ),
        .ch_l_xcvr_rx_eq_dfe_tap_1_atom                         (ch_l_xcvr_rx_eq_dfe_tap_1_atom                ),
        .ch_l_xcvr_rx_external_couple_type_atom                 (ch_l_xcvr_rx_external_couple_type_atom        ),
        .ch_l_tx_pll_bw_sel_atom                                (ch_l_tx_pll_bw_sel_atom                       ),
        .ch_l_xcvr_tx_bonding_category_atom                     (ch_l_xcvr_tx_bonding_category_atom            ),
        .ch_l_xcvr_tx_master_pll_mode_atom                      (ch_l_xcvr_tx_master_pll_mode_atom             ),
        .ch_l_xcvr_rx_cdrdivout_en_atom                         (ch_l_xcvr_rx_cdrdivout_en_atom                ),
        .ch_xcvrif_l_tx_bonding_mode_atom                       (ch_xcvrif_l_tx_bonding_mode_atom              ),
        .ch_xcvrif_l_rx_bonding_mode_atom                       (ch_xcvrif_l_rx_bonding_mode_atom              ),
        .ch_l_speed_grade_atom                                  (ch_l_speed_grade_atom                         ),
        .ch_flux_l_sequencer_reg_en_atom                        (ch_flux_l_sequencer_reg_en_atom               ),
        .ch_usb_mode_atom                                       (ch_usb_mode_atom                              ),
        .ch_pcie_mode_atom                                      (ch_pcie_mode_atom                             ),
        .ch_l_ick_tx_word_clk_hz_atom                           (ch_l_ick_tx_word_clk_hz_atom                  ),
        .ch_l_pcs_ref_clk_hz_atom                               (ch_l_pcs_ref_clk_hz_atom                      ),
        .ch_l_lane_common_ref_clk_hz_atom                       (ch_l_lane_common_ref_clk_hz_atom              ),
        .ch_rx_invert_pin_atom                                  (ch_rx_invert_pin_atom                         ),
        .ch_tx_invert_pin_atom                                  (ch_tx_invert_pin_atom                         ),
        .ch_rx_dl_rx_lat_bit_for_async_atom                     (ch_rx_dl_rx_lat_bit_for_async_atom            ),
        .ch_rx_dl_rxbit_cntr_pma_atom                           (ch_rx_dl_rxbit_cntr_pma_atom                  ),
        .ch_rx_dl_rxbit_rollover_atom                           (ch_rx_dl_rxbit_rollover_atom                  ),
        .ch_eth_rx_clk_hz_atom                                  (ch_eth_rx_clk_hz_atom                         ),
        .ch_eth_tx_clk_hz_atom                                  (ch_eth_tx_clk_hz_atom                         ),
        .ch_clkrx_refclk_cssm_fw_control_atom                   (ch_clkrx_refclk_cssm_fw_control_atom              ),
        .ch_clkrx_refclk_sector_specifies_refclk_ready_atom     (ch_clkrx_refclk_sector_specifies_refclk_ready_atom),
        .ch_local_refclk_cssm_fw_control_atom                   (ch_local_refclk_cssm_fw_control_atom              ),
        .ch_local_refclk_sector_specifies_refclk_ready_atom     (ch_local_refclk_sector_specifies_refclk_ready_atom),
        .ch_flux_l_stmux_rx_demux_sel                           (ch_flux_l_stmux_rx_demux_sel                  ),
        .ch_flux_l_stmux_rx_rxword_clk_demux_sel                (ch_flux_l_stmux_rx_rxword_clk_demux_sel       ),
        .ch_flux_l_stmux_tx_txword_clk_demux_sel                (ch_flux_l_stmux_tx_txword_clk_demux_sel       ),
        .ch_flux_l_stmux_tx_mux_sel                             (ch_flux_l_stmux_tx_mux_sel                    ),
        .ch_flux_l_stmux_tx_txword_clk_mux_sel                  (ch_flux_l_stmux_tx_txword_clk_mux_sel         ),
        .ch_xcvrif_rx_ch_clk_static_mux                         (ch_xcvrif_rx_ch_clk_static_mux                ),
        .ch_xcvrif_tx_ch_clk_static_mux                         (ch_xcvrif_tx_ch_clk_static_mux                )
)
phy_hal_coreip_inst(
        .oflux_xoa_tx_n_l0_ux               (oflux_xoa_tx_n_l0_ux),
        .oflux_xoa_tx_p_l0_ux               (oflux_xoa_tx_p_l0_ux),
        .iflux_xia_rx_n_l0_ux               (iflux_xia_rx_n_l0_ux),
        .iflux_xia_rx_p_l0_ux               (iflux_xia_rx_p_l0_ux),
        .i_ss_async_pldif                   (i_ss_async_pldif        ),
        .o_ss_async_pldif                   (o_ss_async_pldif        ),
        .i_ss_async_pldif_pcie_mux          (i_ss_async_pldif_pcie_mux),
        .i_lavmm_addr                       (i_lavmm_addr),
        .i_lavmm_be                         (i_lavmm_be),
        .i_lavmm_clk                        (i_lavmm_clk),
        .i_lavmm_read                       (i_lavmm_read),
        .i_lavmm_rstn                       (i_lavmm_rstn),
        .i_lavmm_wdata                      (i_lavmm_wdata),
        .i_lavmm_write                      (i_lavmm_write),
        .o_lavmm_rdata                      (o_lavmm_rdata),
        .o_lavmm_rdata_valid                (o_lavmm_rdata_valid),
        .o_lavmm_waitreq                    (o_lavmm_waitreq),
        .i_ft_rx_sclk_sync_ch               (i_ft_rx_sclk_sync_ch),
        .i_ft_tx_sclk_sync_ch               (i_ft_tx_sclk_sync_ch),
        .o_ft_rx_async_pulse_ch             (o_ft_rx_async_pulse_ch),
        .o_ft_tx_async_pulse_ch             (o_ft_tx_async_pulse_ch),
        .o_rxcdrlock2dataa                  (o_rxcdrlock2dataa),
        .i_rst_ux_rx_sfrz                   (i_rst_ux_rx_sfrz),
        .o_rst_flux0_cpi_cmn_busy           (o_rst_flux0_cpi_cmn_busy),
        .o_rst_oflux_rx_srds_rdy            (o_rst_oflux_rx_srds_rdy),
        .o_rst_ux_all_synthlockstatus       (o_rst_ux_all_synthlockstatus),
        .o_rst_ux_rxcdrlockstatus           (o_rst_ux_rxcdrlockstatus),
        .o_ux_tx_ch_ptr_smpl                (o_ux_tx_ch_ptr_smpl),
        .i_ick_sclk_tx                      (i_ick_sclk_tx),
        .i_ick_sclk_rx                      (i_ick_sclk_rx),
        .i_rst_pld_ux_tx_pma_rst_n          (i_rst_pld_ux_tx_pma_rst_n),
        .i_rst_pld_ux_rx_pma_rst_n          (i_rst_pld_ux_rx_pma_rst_n),
        .o_ch_lavmm_xcvrif_rdata            (o_ch_lavmm_xcvrif_rdata),
        .o_ch_lavmm_xcvrif_rdata_valid      (o_ch_lavmm_xcvrif_rdata_valid),
        .o_ch_lavmm_xcvrif_waitreq          (o_ch_lavmm_xcvrif_waitreq),
        .i_ch_lavmm_xcvrif_addr             (i_ch_lavmm_xcvrif_addr),
        .i_ch_lavmm_xcvrif_be               (i_ch_lavmm_xcvrif_be),
        .i_ch_lavmm_xcvrif_clk              (i_ch_lavmm_xcvrif_clk),
        .i_ch_lavmm_xcvrif_read             (i_ch_lavmm_xcvrif_read),
        .i_ch_lavmm_xcvrif_rstn             (i_ch_lavmm_xcvrif_rstn),
        .i_ch_lavmm_xcvrif_wdata            (i_ch_lavmm_xcvrif_wdata),
        .i_ch_lavmm_xcvrif_write            (i_ch_lavmm_xcvrif_write),
//        .i_pld_rx_lat_sclk_ch               (i_pld_rx_lat_sclk_ch),
//        .i_pld_tx_lat_sclk_ch               (i_pld_tx_lat_sclk_ch),
        .o_rx_latency_pulse                 (o_rx_latency_pulse),
        .o_tx_latency_pulse                 (o_tx_latency_pulse),
        .i_xcvrif_tx_mux_data               (i_xcvrif_tx_mux_data),
        .o_rx_data                          (o_rx_data),
        .o_tx_source_sel                    (o_tx_source_sel),
        .i_ch_eth_xcvrif_tx_async           (i_ch_eth_xcvrif_tx_async),
        .i_ch_eth_xcvrif_tx_direct          (i_ch_eth_xcvrif_tx_direct),
        .o_ch_eth_xcvrif_rx_async           (o_ch_eth_xcvrif_rx_async),
        .o_ch_eth_xcvrif_rx_direct          (o_ch_eth_xcvrif_rx_direct),
        .i_rstxcvrif_xcvrif_signal_ok       (i_rstxcvrif_xcvrif_signal_ok),
        .i_rstxcvrif_rx_xcvrif_sfrz_n       (i_rstxcvrif_rx_xcvrif_sfrz_n),
        .i_rstxcvrif_xcvrif_rx_rst_n        (i_rstxcvrif_xcvrif_rx_rst_n),
        .i_rstxcvrif_tx_xcvrif_sfrz_n       (i_rstxcvrif_tx_xcvrif_sfrz_n),
        .i_rstxcvrif_xcvrif_tx_rst_n        (i_rstxcvrif_xcvrif_tx_rst_n),
        .o_pma_rx_sf                        (o_pma_rx_sf),
        .o_rx_fifo_en_sel                   (o_rx_fifo_en_sel      ),
        .o_tx_rst_source_sel                (o_tx_rst_source_sel   ),
        .i_ch_xcvrif_rx_fifo_rd_en          (i_ch_xcvrif_rx_fifo_rd_en),
        .o_ch_xcvrif_rx_fifo_rd_en          (o_ch_xcvrif_rx_fifo_rd_en),
        .i_ch_xcvrif_tx_fifo_rd_en          (i_ch_xcvrif_tx_fifo_rd_en),
        .o_ch_xcvrif_tx_fifo_rd_en          (o_ch_xcvrif_tx_fifo_rd_en),
//        .i_xcvr_rx_ch_clk                   (i_xcvr_rx_ch_clk   ),
//        .i_xcvr_tx_ch_clk                   (i_xcvr_tx_ch_clk   ),
        .o_ux_rxuser1_sel                   (o_ux_rxuser1_sel      ),
        .o_ux_rxuser2_sel                   (o_ux_rxuser2_sel      ),
        .o_ux_txuser1_sel                   (o_ux_txuser1_sel      ),
        .o_ux_txuser2_sel                   (o_ux_txuser2_sel      ),
        .o_pcs_rxpostdiv                    (o_pcs_rxpostdiv            ),
        .o_pcs_rxword                       (o_pcs_rxword               ),
        .o_ux_txlc_clk                      (o_ux_txlc_clk       ),
        .o_ock_pcs_txword                   (o_ock_pcs_txword           ),
        .o_tx_xcvr_wordclk_sel              (o_tx_xcvr_wordclk_sel ),
        .o_rx_xcvr_wordclk_sel              (o_rx_xcvr_wordclk_sel ),
        .i_eth_rx_ch_clk                    (i_eth_rx_ch_clk            ),
//        .i_eth_tx_ch_clk                    (i_eth_tx_ch_clk            ),       
        .uxwrap_bus_in                      (uxwrap_bus_in                      ),      
        .uxwrap_bus_out                     (uxwrap_bus_out                    ) ,
        .o_lavmm_addr                       (o_lavmm_addr                      ) ,
        .o_lavmm_be                         (o_lavmm_be                        ) ,
        .o_lavmm_clk                        (o_lavmm_clk                       ) ,
        .o_lavmm_read                       (o_lavmm_read                      ) ,
        .o_lavmm_rstn                       (o_lavmm_rstn                      ) ,
        .o_lavmm_wdata                      (o_lavmm_wdata                     ) ,
        .o_lavmm_write                      (o_lavmm_write                     ) ,
        .i_lavmm_rdata                      (i_lavmm_rdata                     ) ,
        .i_lavmm_rdata_valid                (i_lavmm_rdata_valid                ),
        .i_lavmm_waitreq                    (i_lavmm_waitreq                   ) ,
        .o_sclk_return_sel_rx               (o_sclk_return_sel_rx              ) ,
        .o_sclk_return_sel_tx               (o_sclk_return_sel_tx               ),
        .o_ick_sclk_rx                      (o_ick_sclk_rx                     ) ,
        .i_sync_common_control              (i_sync_common_control             ) ,
        .o_ft_rx_sclk_sync_ch               (o_ft_rx_sclk_sync_ch              ) ,
        .o_ft_tx_sclk_sync_ch               (o_ft_tx_sclk_sync_ch              ) ,
        .o_rst_ux_rx_pma_rst_n              (o_rst_ux_rx_pma_rst_n             ) ,
        .o_rst_ux_tx_pma_rst_n              (o_rst_ux_tx_pma_rst_n             ) ,
        .o_ick_pcs_txword                   (o_ick_pcs_txword                   ),
        .o_tx_dl_ch_bit                     (o_tx_dl_ch_bit                     ),
        .i_dat_pcs_measlatbit               (i_dat_pcs_measlatbit               ),
        .i_ft_rx_async_pulse_ch             (i_ft_rx_async_pulse_ch            ) ,
        .i_ft_tx_async_pulse_ch             (i_ft_tx_async_pulse_ch             ),
        .i_rx_dl_ch_bit                     (i_rx_dl_ch_bit                     ),
        .i_ux_rxuser1_sel                   (i_ux_rxuser1_sel                  ) ,
        .i_ux_rxuser2_sel                   (i_ux_rxuser2_sel                   ),
        .i_ux_txuser1_sel                   (i_ux_txuser1_sel                  ) ,
        .i_ux_txuser2_sel                   (i_ux_txuser2_sel                   ),
        .o_octl_pcs_txstatus_a              (o_octl_pcs_txstatus_a              ),
        .i_ictl_pcs_txenable_a              (i_ictl_pcs_txenable_a             ) ,
        .i_sync_cfg_data                    (i_sync_cfg_data                    ),
        .i_sync_interface_control           (i_sync_interface_control           ),
        .o_tx_data                          (o_tx_data                          ),
        .i_rx_data                          (i_rx_data                          ),
        .o_sm_flux_ingress                  (o_sm_flux_ingress                 ) ,
        .i_sm_flux_egress                   (i_sm_flux_egress                  ) ,
        .i_flux_cpi_int                     (i_flux_cpi_int                    ) ,
        .i_flux_int                         (i_flux_int                        ) ,
        .i_oflux_octl_pcs_txptr_smpl_lane   (i_oflux_octl_pcs_txptr_smpl_lane  ) ,
        .o_ick_sclk_tx                      (o_ick_sclk_tx                     ) ,
        .i_flux_srds_rdy                    (i_flux_srds_rdy                    ),
        .i_pcs_rxword                       (i_pcs_rxword                      ) ,
        .i_pcs_rxpostdiv                    (i_pcs_rxpostdiv                    ),
        .i_ock_pcs_txword                   (i_ock_pcs_txword                  ) ,
        .o_dat_pcs_measlatrndtripbit        (o_dat_pcs_measlatrndtripbit                  ) ,
//        .i_dpma_refclk                      (i_dpma_refclk                              ) ,   //Connected this from cnoc atom in phy_hal_coreip.sv
        .o_ock_pcs_cdrfbclk                 (o_ock_pcs_cdrfbclk                           ) ,
        .o_ock_pcs_ref                      (o_ock_pcs_ref                        ), 
        .o_pcie_pcs                         (o_pcie_pcs),
        .i_pcie_pcs                         (i_pcie_pcs),
        .i_sel_rxword_clk                   (i_sel_rxword_clk),
        .i_xcvr_txword_clk                  (i_xcvr_txword_clk),
        .o_pcie_rxword_clk                  (o_pcie_rxword_clk),
        .o_eth_rxword_clk                   (o_eth_rxword_clk),
        .o_pcie_txword_clk                  (o_pcie_txword_clk),
        .o_eth_txword_clk                   (o_eth_txword_clk),
        .o_eth_rx_ch_clk                    (o_eth_rx_ch_clk),
        .o_eth_tx_ch_clk                    (o_eth_tx_ch_clk),
        .ioack_ref_left_p_ux_bidir_in       (ioack_ref_left_p_ux_bidir_in),
        .ioack_hsref_left_p_ux_bidir_in     (ioack_hsref_left_p_ux_bidir_in),
        .ioack_cdrdiv_left_ux_bidir_in      (ioack_cdrdiv_left_ux_bidir_in),
        .ioack_synthdiv1_left_ux_bidir_in   (ioack_synthdiv1_left_ux_bidir_in),
        .ioack_synthdiv2_left_ux_bidir_in   (ioack_synthdiv2_left_ux_bidir_in),
        .ioack_cdrdiv_left_ux_bidir_out     (ioack_cdrdiv_left_ux_bidir_out),
        .ioack_synthdiv1_left_ux_bidir_out  (ioack_synthdiv1_left_ux_bidir_out),
        .ioack_synthdiv2_left_ux_bidir_out  (ioack_synthdiv2_left_ux_bidir_out),
        .i_quartus_flux_s_to_ingress        (i_quartus_flux_s_to_ingress),        
        .i_rstxcvrif_xcvrif_tx_rd_rst_n     (i_rstxcvrif_xcvrif_tx_rd_rst_n),        
        .i_rstxcvrif_xcvrif_tx_wr_rst_n     (i_rstxcvrif_xcvrif_tx_wr_rst_n),        
        .o_tx_rst_rd_sync_rst_n             (o_tx_rst_rd_sync_rst_n),        
        .o_tx_rst_wr_sync_rst_n             (o_tx_rst_wr_sync_rst_n),        

//KAHUAT_EDIT
        .o_rxeq_best_eye_vala               (o_rxeq_best_eye_vala),
        .o_rxeq_donea                       (o_rxeq_donea),
        .o_rxmargin_nacka                   (o_rxmargin_nacka),
        .o_rxmargin_statusa                 (o_rxmargin_statusa),
        .o_rxsignaldetect_lfpsa             (o_rxsignaldetect_lfpsa),
        .o_rxsignaldetecta                  (o_rxsignaldetecta),
        .o_rxmargin_status_gray             (o_rxmargin_status_gray),
        .o_rxstatusa                        (o_rxstatusa),
        .o_synthlcfast_postdiv              (o_synthlcfast_postdiv),
        .o_synthlcmed_postdiv               (o_synthlcmed_postdiv),
        .o_synthlcslow_postdiv              (o_synthlcslow_postdiv),
        .o_txdetectrx_acka                  (o_txdetectrx_acka),
        .o_txdetectrx_statct                (o_txdetectrx_statct),
        .o_txstatusa                        (o_txstatusa),
        .i_pcs_pipe_rstn                    (i_pcs_pipe_rstn),
        .i_ux_ock_pma_clk                   (i_ux_ock_pma_clk),
        .i_lfps_ennt                        (i_lfps_ennt),
        .i_pcie_l1ctrla                     (i_pcie_l1ctrla),
        .i_pma_cmn_ctrl                     (i_pma_cmn_ctrl),
        .i_pma_ctrl                         (i_pma_ctrl),
        .i_pcie_pcs_rx_rst                  (i_pcie_pcs_rx_rst),
        .i_pcie_pcs_tx_rst                  (i_pcie_pcs_tx_rst),
        .i_rxeiosdetectstata                (i_rxeiosdetectstata),
        .i_rxeq_precal_code_selnt           (i_rxeq_precal_code_selnt),
        .i_rxeq_starta                      (i_rxeq_starta),
        .i_rxeq_static_ena                  (i_rxeq_static_ena),
        .i_rxmargin_direction_nt            (i_rxmargin_direction_nt),
        .i_rxmargin_mode_nt                 (i_rxmargin_mode_nt),
        .i_rxmargin_offset_change_a         (i_rxmargin_offset_change_a),
        .i_rxmargin_offset_nt               (i_rxmargin_offset_nt),
        .i_rxmargin_start_a                 (i_rxmargin_start_a),
        .i_rxpstate                         (i_rxpstate),
        .i_rxrate                           (i_rxrate),
        .i_rxterm_hiz_ena                   (i_rxterm_hiz_ena),
        .i_rxwidth                          (i_rxwidth),
        .i_tstbus_lane                      (i_tstbus_lane),
        .i_txbeacona                        (i_txbeacona),
        .i_txclkdivrate                     (i_txclkdivrate),
        .i_txdetectrx_reqa                  (i_txdetectrx_reqa),
        .i_txdrv_levn                       (i_txdrv_levn),
        .i_txdrv_levnm1                     (i_txdrv_levnm1),
        .i_txdrv_levnm2                     (i_txdrv_levnm2),
        .i_txdrv_levnp1                     (i_txdrv_levnp1),
        .i_txdrv_slew                       (i_txdrv_slew),
        .i_txelecidle                       (i_txelecidle),
        .i_txpstate                         (i_txpstate),
        .i_txrate                           (i_txrate),
        .i_txwidth                          (i_txwidth)
);

endmodule

