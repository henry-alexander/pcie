// system_intel_pcie_gts_0_one_lane_pcie_hal_pldif_hal_2100_agcatrq.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_intel_pcie_gts_0_one_lane_pcie_hal_pldif_hal_2100_agcatrq #(
		parameter       ch_pldif_l_tx_en_atom                    = "TRUE",
		parameter       ch_pldif_l_rx_en_atom                    = "TRUE",
		parameter       ch_pldif_l_duplex_mode_atom              = "DUPLEX_MODE_DUPLEX",
		parameter       ch_pldif_l_tx_fifo_mode_atom             = "TX_FIFO_MODE_PHASE_COMP",
		parameter       ch_pldif_l_tx_fifo_width_atom            = "TX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH",
		parameter       ch_pldif_l_rx_fifo_mode_atom             = "RX_FIFO_MODE_PHASE_COMP",
		parameter       ch_pldif_l_rx_fifo_width_atom            = "RX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH",
		parameter       ch_pldif_l_tx_clkout1_divider_atom       = "TX_CLKOUT1_DIVIDER_DIV1",
		parameter       ch_pldif_l_tx_clkout2_divider_atom       = "TX_CLKOUT2_DIVIDER_DIV1",
		parameter       ch_pldif_l_rx_clkout1_divider_atom       = "RX_CLKOUT1_DIVIDER_DIV1",
		parameter       ch_pldif_l_rx_clkout2_divider_atom       = "RX_CLKOUT2_DIVIDER_DIV1",
		parameter       ch_pldif_l_dr_enabled_atom               = "DR_ENABLED_DR_DISABLED",
		parameter       ch_pldif_l_ptp_enable_atom               = "PTP_ENABLE_DISABLE",
		parameter       ch_pldif_l_tx_user1_clk_dynamic_mux_atom = "TX_USER1_CLK_DYNAMIC_MUX_UX",
		parameter       ch_pldif_l_tx_user2_clk_dynamic_mux_atom = "TX_USER2_CLK_DYNAMIC_MUX_UX",
		parameter       ch_pldif_l_rx_user1_clk_dynamic_mux_atom = "RX_USER1_CLK_DYNAMIC_MUX_UX",
		parameter       ch_pldif_l_rx_user2_clk_dynamic_mux_atom = "RX_USER2_CLK_DYNAMIC_MUX_UX",
		parameter       ch_pldif_l_sup_mode_atom                 = "SUP_MODE_USER_MODE",
		parameter       ch_pldif_l_tx_mac_en_atom                = "FALSE",
		parameter       ch_pldif_l_pld_channel_identifier_atom   = "PLD_CHANNEL_IDENTIFIER_PHIP",
		parameter[35:0] ch_pldif_rx_fifo_wr_clk_hz_atom          = 36'b000000010001111000011010001100000000,
		parameter[35:0] ch_pldif_tx_fifo_rd_clk_hz_atom          = 36'b000000010001111000011010001100000000,
		parameter       ch_pldif_l_rx_dyn_mux_atom               = "RX_DYN_MUX_XCVRIF",
		parameter       ch_pldif_l_tx_bond_location_atom         = "TX_BOND_LOCATION_FIRST",
		parameter       ch_pldif_l_rx_bond_location_atom         = "RX_BOND_LOCATION_UNUSED",
		parameter       ch_pldif_l_ehip_lb_tx_rx_atom            = "EHIP_LB_TX_RX_DISABLE",
		parameter       ch_pldif_l_ehip_lb_txmac_rx_atom         = "EHIP_LB_TXMAC_RX_DISABLE",
		parameter       ch_pldif_l_rx_pmadir_singlewidth_en_atom = "RX_PMADIR_SINGLEWIDTH_EN_DISABLE",
		parameter       ch_pldif_l_tx_pmadir_singlewidth_en_atom = "TX_PMADIR_SINGLEWIDTH_EN_DISABLE",
		parameter       ch_pldif_l_ehip_lb_txpcs_rx_atom         = "EHIP_LB_TXPCS_RX_DISABLE",
		parameter       ch_pcs_l_tx_bond_size_atom               = "TX_BOND_SIZE_X4",
		parameter       ch_pcs_l_rx_bond_size_atom               = "RX_BOND_SIZE_UNUSED",
		parameter       ch_vc_rx_pldif_wm_en_atom                = "VC_RX_PLDIF_WM_EN_DISABLE",
		parameter       ch_pldif_l_stmux_tx_demux_sel            = "SEL_PCIE",
		parameter       ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel  = "SEL_PCIE",
		parameter       ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel  = "SEL_PCIE",
		parameter       ch_pldif_l_stmux_rx_mux_sel              = "SEL_PCIE",
		parameter       ch_l_xcvr_rx_preloaded_hardware_configs  = "PCIE_GEN4",
		parameter       ch_l_xcvr_tx_preloaded_hardware_configs  = "PCIE_GEN4"
	) (
		input  wire [79:0] i_hio_txdata,                                       //                                       i_hio_txdata.data
		input  wire [9:0]  i_hio_txdata_extra,                                 //                                 i_hio_txdata_extra.data
		input  wire        i_hio_txdata_fifo_wr_en,                            //                            i_hio_txdata_fifo_wr_en.fifowriteenable
		output wire        o_hio_txdata_fifo_wr_empty,                         //                         o_hio_txdata_fifo_wr_empty.fifowritestatus
		output wire        o_hio_txdata_fifo_wr_pempty,                        //                        o_hio_txdata_fifo_wr_pempty.fifowritestatus
		output wire        o_hio_txdata_fifo_wr_full,                          //                          o_hio_txdata_fifo_wr_full.fifowritestatus
		output wire        o_hio_txdata_fifo_wr_pfull,                         //                         o_hio_txdata_fifo_wr_pfull.fifowritestatus
		output wire [79:0] o_hio_rxdata,                                       //                                       o_hio_rxdata.data
		output wire [9:0]  o_hio_rxdata_extra,                                 //                                 o_hio_rxdata_extra.data
		output wire        o_hio_rxdata_fifo_rd_empty,                         //                         o_hio_rxdata_fifo_rd_empty.fiforeadenable
		output wire        o_hio_rxdata_fifo_rd_pempty,                        //                        o_hio_rxdata_fifo_rd_pempty.fiforeadstatus
		output wire        o_hio_rxdata_fifo_rd_full,                          //                          o_hio_rxdata_fifo_rd_full.fiforeadstatus
		output wire        o_hio_rxdata_fifo_rd_pfull,                         //                         o_hio_rxdata_fifo_rd_pfull.fiforeadstatus
		input  wire        i_hio_rxdata_fifo_rd_en,                            //                            i_hio_rxdata_fifo_rd_en.fiforeadstatus
		input  wire        i_hio_ptp_rst_n,                                    //                                    i_hio_ptp_rst_n.data
		input  wire        i_hio_ehip_rx_rst_n,                                //                                i_hio_ehip_rx_rst_n.data
		input  wire        i_hio_ehip_tx_rst_n,                                //                                i_hio_ehip_tx_rst_n.data
		input  wire        i_hio_ehip_signal_ok,                               //                               i_hio_ehip_signal_ok.data
		input  wire        i_hio_sfreeze_2_r03f_rx_mac_srfz_n,                 //                 i_hio_sfreeze_2_r03f_rx_mac_srfz_n.data
		input  wire        i_hio_sfreeze_3_c2f_tx_deskew_srfz_n,               //               i_hio_sfreeze_3_c2f_tx_deskew_srfz_n.data
		input  wire        i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n,                 //                 i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n.data
		output wire        o_hio_rstepcs_rx_pcs_fully_aligned,                 //                 o_hio_rstepcs_rx_pcs_fully_aligned.status
		input  wire        i_hio_rstfec_fec_rx_rst_n,                          //                          i_hio_rstfec_fec_rx_rst_n.data
		input  wire        i_hio_rstfec_fec_tx_rst_n,                          //                          i_hio_rstfec_fec_tx_rst_n.data
		input  wire        i_hio_rstfec_fec_csr_ret,                           //                           i_hio_rstfec_fec_csr_ret.data
		output wire        o_hio_rstfec_fec_rx_rdy_n,                          //                          o_hio_rstfec_fec_rx_rdy_n.status
		input  wire        i_hio_rstfec_rx_fec_sfrz_n,                         //                         i_hio_rstfec_rx_fec_sfrz_n.data
		input  wire        i_hio_rstfec_tx_fec_sfrz_n,                         //                         i_hio_rstfec_tx_fec_sfrz_n.data
		input  wire        i_hio_rstxcvrif_xcvrif_rx_rst_n,                    //                    i_hio_rstxcvrif_xcvrif_rx_rst_n.data
		input  wire        i_hio_rstxcvrif_xcvrif_tx_rst_n,                    //                    i_hio_rstxcvrif_xcvrif_tx_rst_n.data
		input  wire        i_hio_rstxcvrif_xcvrif_signal_ok,                   //                   i_hio_rstxcvrif_xcvrif_signal_ok.data
		input  wire        i_hio_rstxcvrif_rx_xcvrif_sfrz_n,                   //                   i_hio_rstxcvrif_rx_xcvrif_sfrz_n.data
		input  wire        i_hio_rstxcvrif_tx_xcvrif_sfrz_n,                   //                   i_hio_rstxcvrif_tx_xcvrif_sfrz_n.data
		input  wire        i_hio_rst_pld_clrhip,                               //                               i_hio_rst_pld_clrhip.data
		input  wire        i_hio_rst_pld_clrpcs,                               //                               i_hio_rst_pld_clrpcs.data
		input  wire        i_hio_rst_pld_perstn,                               //                               i_hio_rst_pld_perstn.data
		input  wire        i_hio_rst_pld_ready,                                //                                i_hio_rst_pld_ready.status
		input  wire        i_hio_rst_pld_adapter_rx_pld_rst_n,                 //                 i_hio_rst_pld_adapter_rx_pld_rst_n.data
		input  wire        i_hio_rst_pld_adapter_tx_pld_rst_n,                 //                 i_hio_rst_pld_adapter_tx_pld_rst_n.data
		input  wire        i_hio_rst_ux_rx_pma_rst_n,                          //                          i_hio_rst_ux_rx_pma_rst_n.data
		input  wire        i_hio_rst_ux_rx_sfrz,                               //                               i_hio_rst_ux_rx_sfrz.data
		input  wire        i_hio_rst_ux_tx_pma_rst_n,                          //                          i_hio_rst_ux_tx_pma_rst_n.data
		output wire        o_hio_rst_flux0_cpi_cmn_busy,                       //                       o_hio_rst_flux0_cpi_cmn_busy.status
		output wire        o_hio_rst_oflux_rx_srds_rdy,                        //                        o_hio_rst_oflux_rx_srds_rdy.status
		output wire        o_hio_rst_ux_all_synthlockstatus,                   //                   o_hio_rst_ux_all_synthlockstatus.status
		output wire        o_hio_rst_ux_octl_pcs_rxstatus,                     //                     o_hio_rst_ux_octl_pcs_rxstatus.status
		output wire        o_hio_rst_ux_octl_pcs_txstatus,                     //                     o_hio_rst_ux_octl_pcs_txstatus.status
		output wire        o_hio_rst_ux_rxcdrlock2data,                        //                        o_hio_rst_ux_rxcdrlock2data.data
		output wire        o_hio_rst_ux_rxcdrlockstatus,                       //                       o_hio_rst_ux_rxcdrlockstatus.status
		output wire        o_ss_ehip_rx_rst_n,                                 //                                 o_ss_ehip_rx_rst_n.data
		output wire        o_ss_ehip_tx_rst_n,                                 //                                 o_ss_ehip_tx_rst_n.data
		output wire        o_ss_ehip_signal_ok,                                //                                o_ss_ehip_signal_ok.data
		output wire        o_ss_sfreeze_2_r03f_rx_mac_srfz_n,                  //                  o_ss_sfreeze_2_r03f_rx_mac_srfz_n.data
		output wire        o_ss_sfreeze_3_c2f_tx_deskew_srfz_n,                //                o_ss_sfreeze_3_c2f_tx_deskew_srfz_n.data
		input  wire        i_ss_rstepcs_rx_pcs_fully_aligned,                  //                  i_ss_rstepcs_rx_pcs_fully_aligned.status
		output wire        o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n,                  //                  o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n.data
		output wire        o_ss_rstfec_fec_rx_rst_n,                           //                           o_ss_rstfec_fec_rx_rst_n.data
		output wire        o_ss_rstfec_fec_tx_rst_n,                           //                           o_ss_rstfec_fec_tx_rst_n.data
		output wire        o_ss_rstfec_fec_csr_ret,                            //                            o_ss_rstfec_fec_csr_ret.data
		input  wire        i_ss_rstfec_fec_rx_rdy_n,                           //                           i_ss_rstfec_fec_rx_rdy_n.status
		output wire        o_ss_rstfec_rx_fec_sfrz_n,                          //                          o_ss_rstfec_rx_fec_sfrz_n.data
		output wire        o_ss_rstfec_tx_fec_sfrz_n,                          //                          o_ss_rstfec_tx_fec_sfrz_n.data
		output wire        o_ss_rstxcvrif_xcvrif_rx_rst_n,                     //                     o_ss_rstxcvrif_xcvrif_rx_rst_n.data
		output wire        o_ss_rstxcvrif_xcvrif_tx_rst_n,                     //                     o_ss_rstxcvrif_xcvrif_tx_rst_n.data
		output wire        o_ss_rstxcvrif_xcvrif_signal_ok,                    //                    o_ss_rstxcvrif_xcvrif_signal_ok.data
		output wire        o_ss_rstxcvrif_rx_xcvrif_sfrz_n,                    //                    o_ss_rstxcvrif_rx_xcvrif_sfrz_n.data
		output wire        o_ss_rstxcvrif_tx_xcvrif_sfrz_n,                    //                    o_ss_rstxcvrif_tx_xcvrif_sfrz_n.data
		output wire        o_ss_rst_ux_rx_pma_rst_n,                           //                           o_ss_rst_ux_rx_pma_rst_n.data
		output wire        o_ss_rst_ux_rx_sfrz,                                //                                o_ss_rst_ux_rx_sfrz.data
		output wire        o_ss_rst_ux_tx_pma_rst_n,                           //                           o_ss_rst_ux_tx_pma_rst_n.data
		input  wire        i_ss_rst_flux0_cpi_cmn_busy,                        //                        i_ss_rst_flux0_cpi_cmn_busy.status
		input  wire        i_ss_rst_oflux_rx_srds_rdy,                         //                         i_ss_rst_oflux_rx_srds_rdy.status
		input  wire        i_ss_rst_ux_all_synthlockstatus,                    //                    i_ss_rst_ux_all_synthlockstatus.status
		input  wire        i_ss_rst_ux_octl_pcs_rxstatus,                      //                      i_ss_rst_ux_octl_pcs_rxstatus.status
		input  wire        i_ss_rst_ux_octl_pcs_txstatus,                      //                      i_ss_rst_ux_octl_pcs_txstatus.status
		input  wire        i_ss_rst_ux_rxcdrlock2data,                         //                         i_ss_rst_ux_rxcdrlock2data.data
		input  wire        i_ss_rst_ux_rxcdrlockstatus,                        //                        i_ss_rst_ux_rxcdrlockstatus.status
		input  wire        i_hio_pld_reset_clk_row,                            //                            i_hio_pld_reset_clk_row.status
		input  wire [11:0] i_ss_eth_fec_rx_async,                              //                                        asyncdata_0.data
		input  wire        i_ss_eth_fec_rx_direct,                             //                                        asyncdata_1.data
		output wire [6:0]  o_ss_eth_fec_tx_async,                              //                                        asyncdata_2.data
		output wire        o_ss_eth_fec_tx_direct,                             //                                        asyncdata_3.data
		input  wire [13:0] i_ss_eth_mac_rx_async,                              //                                        asyncdata_4.data
		input  wire        i_ss_eth_mac_rx_direct,                             //                                        asyncdata_5.data
		output wire [13:0] o_ss_eth_mac_tx_async,                              //                                        asyncdata_6.data
		output wire        o_ss_eth_mac_tx_direct,                             //                                        asyncdata_7.data
		input  wire [13:0] i_ss_eth_pcs_rx_async,                              //                                        asyncdata_8.data
		input  wire        i_ss_eth_pcs_rx_direct,                             //                                        asyncdata_9.data
		output wire [7:0]  o_ss_eth_pcs_tx_async,                              //                                       asyncdata_10.data
		output wire        o_ss_eth_pcs_tx_direct,                             //                                       asyncdata_11.data
		input  wire [13:0] i_ss_eth_xcvrif_rx_async,                           //                                       asyncdata_12.data
		input  wire        i_ss_eth_xcvrif_rx_direct,                          //                                       asyncdata_13.data
		output wire [6:0]  o_ss_eth_xcvrif_tx_async,                           //                                       asyncdata_14.data
		output wire        o_ss_eth_xcvrif_tx_direct,                          //                                       asyncdata_15.data
		input  wire [87:0] i_ss_pcie_ctrl_rx_async,                            //                                       asyncdata_16.data
		input  wire [7:0]  i_ss_pcie_ctrl_rx_direct,                           //                                       asyncdata_17.data
		output wire [79:0] o_ss_uxquad_async,                                  //                                       asyncdata_20.data
		output wire [79:0] o_ss_uxquad_async_pcie_mux,                         //                                       asyncdata_21.data
		input  wire [49:0] i_ss_uxquad_async,                                  //                                       asyncdata_22.data
		input  wire [79:0] i_hio_uxquad_async,                                 //                                       asyncdata_23.data
		input  wire [79:0] i_hio_uxquad_async_pcie_mux,                        //                                       asyncdata_24.data
		output wire [49:0] o_hio_uxquad_async,                                 //                                       asyncdata_25.data
		input  wire [99:0] i_hio_txdata_async,                                 //                                       asyncdata_26.data
		input  wire [9:0]  i_hio_txdata_direct,                                //                                       asyncdata_27.data
		output wire [99:0] o_hio_rxdata_async,                                 //                                       asyncdata_28.data
		output wire [9:0]  o_hio_rxdata_direct,                                //                                       asyncdata_29.data
		output wire [31:0] o_hio_lavmm_rdata,                                  //                                     reconfig_lavmm.readdata
		output wire        o_hio_lavmm_rdata_valid,                            //                                                   .readdatavalid
		output wire        o_hio_lavmm_waitreq,                                //                                                   .waitrequest
		input  wire [20:0] i_hio_lavmm_addr,                                   //                                                   .address
		input  wire [3:0]  i_hio_lavmm_be,                                     //                                                   .byteenable
		input  wire        i_hio_lavmm_read,                                   //                                                   .read
		input  wire [31:0] i_hio_lavmm_wdata,                                  //                                                   .writedata
		input  wire        i_hio_lavmm_write,                                  //                                                   .write
		input  wire        i_hio_lavmm_clk,                                    //                                 reconfig_lavmm_clk.clk
		input  wire        i_hio_lavmm_rstn,                                   //                                 reconfig_lavmm_rst.reset
		input  wire [31:0] i_ss_lavmm_pcie_rdata,                              //                                      reconfig_pcie.readdata
		input  wire        i_ss_lavmm_pcie_rdata_valid,                        //                                                   .readdatavalid
		input  wire        i_ss_lavmm_pcie_waitreq,                            //                                                   .waitrequest
		output wire [16:0] o_ss_lavmm_pcie_addr,                               //                                                   .address
		output wire [3:0]  o_ss_lavmm_pcie_be,                                 //                                                   .byteenable
		output wire        o_ss_lavmm_pcie_read,                               //                                                   .read
		output wire [31:0] o_ss_lavmm_pcie_wdata,                              //                                                   .writedata
		output wire        o_ss_lavmm_pcie_write,                              //                                                   .write
		output wire        o_ss_lavmm_pcie_clk,                                //                                  reconfig_pcie_clk.clk
		output wire        o_ss_lavmm_pcie_rstn,                               //                                  reconfig_pcie_rst.reset
		output wire        o_hio_user_rx_clk1_clk,                             //                             o_hio_user_rx_clk1_clk.clk
		output wire        o_hio_user_rx_clk2_clk,                             //                             o_hio_user_rx_clk2_clk.clk
		output wire        o_hio_user_tx_clk1_clk,                             //                             o_hio_user_tx_clk1_clk.clk
		output wire        o_hio_user_tx_clk2_clk,                             //                             o_hio_user_tx_clk2_clk.clk
		input  wire        i_ux_chnl_refclk_mux,                               //                               i_ux_chnl_refclk_mux.clk
		output wire        o_hio_ux_chnl_refclk_mux,                           //                           o_hio_ux_chnl_refclk_mux.data
		input  wire        i_hio_pld_rx_clk_in_row_clk,                        //                        i_hio_pld_rx_clk_in_row_clk.clk
		input  wire        i_hio_pld_tx_clk_in_row_clk,                        //                        i_hio_pld_tx_clk_in_row_clk.clk
		input  wire        i_hio_det_lat_rx_dl_clk,                            //                            i_hio_det_lat_rx_dl_clk.clk
		input  wire        i_hio_det_lat_rx_mux_select,                        //                        i_hio_det_lat_rx_mux_select.muxsel
		input  wire        i_hio_det_lat_rx_sclk_flop,                         //                         i_hio_det_lat_rx_sclk_flop.clk
		input  wire        i_hio_det_lat_rx_sclk_gen_clk,                      //                      i_hio_det_lat_rx_sclk_gen_clk.clk
		input  wire        i_hio_det_lat_rx_trig_flop,                         //                         i_hio_det_lat_rx_trig_flop.clk
		input  wire        i_hio_det_lat_sampling_clk,                         //                         i_hio_det_lat_sampling_clk.clk
		input  wire        i_hio_det_lat_tx_dl_clk,                            //                            i_hio_det_lat_tx_dl_clk.clk
		input  wire        i_hio_det_lat_tx_mux_select,                        //                        i_hio_det_lat_tx_mux_select.muxsel
		input  wire        i_hio_det_lat_tx_sclk_flop,                         //                         i_hio_det_lat_tx_sclk_flop.clk
		input  wire        i_hio_det_lat_tx_sclk_gen_clk,                      //                      i_hio_det_lat_tx_sclk_gen_clk.clk
		input  wire        i_hio_det_lat_tx_trig_flop,                         //                         i_hio_det_lat_tx_trig_flop.clk
		output wire        o_hio_det_lat_rx_async_dl_sync,                     //                     o_hio_det_lat_rx_async_dl_sync.syncsignal
		output wire        o_hio_det_lat_rx_async_pulse,                       //                       o_hio_det_lat_rx_async_pulse.syncsignal
		output wire        o_hio_det_lat_rx_async_sample_sync,                 //                 o_hio_det_lat_rx_async_sample_sync.syncsignal
		output wire        o_hio_det_lat_rx_sclk_sample_sync,                  //                  o_hio_det_lat_rx_sclk_sample_sync.syncsignal
		output wire        o_hio_det_lat_rx_trig_sample_sync,                  //                  o_hio_det_lat_rx_trig_sample_sync.syncsignal
		output wire        o_hio_det_lat_tx_async_dl_sync,                     //                     o_hio_det_lat_tx_async_dl_sync.syncsignal
		output wire        o_hio_det_lat_tx_async_pulse,                       //                       o_hio_det_lat_tx_async_pulse.syncsignal
		output wire        o_hio_det_lat_tx_async_sample_sync,                 //                 o_hio_det_lat_tx_async_sample_sync.syncsignal
		output wire        o_hio_det_lat_tx_sclk_sample_sync,                  //                  o_hio_det_lat_tx_sclk_sample_sync.syncsignal
		output wire        o_hio_det_lat_tx_trig_sample_sync,                  //                  o_hio_det_lat_tx_trig_sample_sync.syncsignal
		output wire        o_hio_xcvrif_rx_latency_pulse,                      //                      o_hio_xcvrif_rx_latency_pulse.syncsignal
		output wire        o_hio_xcvrif_tx_latency_pulse,                      //                      o_hio_xcvrif_tx_latency_pulse.syncsignal
		output wire        o_ss_det_lat_rx_sclk_clk,                           //                           o_ss_det_lat_rx_sclk_clk.clk
		output wire        o_ss_det_lat_rx_sclk_sync,                          //                          o_ss_det_lat_rx_sclk_sync.syncsignal
		output wire        o_ss_det_lat_tx_sclk_clk,                           //                           o_ss_det_lat_tx_sclk_clk.clk
		output wire        o_ss_det_lat_tx_sclk_sync,                          //                          o_ss_det_lat_tx_sclk_sync.syncsignal
		input  wire        i_ss_det_lat_rx_async_pulse,                        //                        i_ss_det_lat_rx_async_pulse.syncsignal
		input  wire        i_ss_det_lat_tx_async_pulse,                        //                        i_ss_det_lat_tx_async_pulse.syncsignal
		input  wire        i_ss_xcvrif_rx_latency_pulse,                       //                       i_ss_xcvrif_rx_latency_pulse.syncsignal
		input  wire        i_ss_xcvrif_tx_latency_pulse,                       //                       i_ss_xcvrif_tx_latency_pulse.syncsignal
		input  wire        i_ux_tx_ch_ptr_smpl,                                //                                i_ux_tx_ch_ptr_smpl.syncsignal
		output wire        o_hio_ux_tx_ch_ptr_smpl,                            //                            o_hio_ux_tx_ch_ptr_smpl.syncsignal
		input  wire        i_deskew_rx_ch_clk,                                 //                                 i_deskew_rx_ch_clk.clk
		input  wire        i_deskew_tx_ch_clk,                                 //                                 i_deskew_tx_ch_clk.clk
		output wire        o_marker_found,                                     //                                     o_marker_found.status
		input  wire        i_marker_found_up,                                  //                                  i_marker_found_up.status
		input  wire        i_marker_found_dn,                                  //                                  i_marker_found_dn.status
		output wire [42:0] o_ch_pld_tx_deskewed_data,                          //                          o_ch_pld_tx_deskewed_data.data
		output wire [8:0]  o_ch_ptp_tx_deskewed_data,                          //                          o_ch_ptp_tx_deskewed_data.data
		input  wire [7:0]  i_ch_ptp_rx_data,                                   //                                   i_ch_ptp_rx_data.data
		input  wire        i_ch_tx_mac_ready,                                  //                                  i_ch_tx_mac_ready.status
		input  wire        i_ch_rx_mac_inframe,                                //                                i_ch_rx_mac_inframe.status
		output wire        o_ch_tx_mac_valid,                                  //                                  o_ch_tx_mac_valid.status
		input  wire        i_ptp_rx_dsk_marker,                                //                                i_ptp_rx_dsk_marker.status
		input  wire        i_ptp_mas_wm,                                       //                                       i_ptp_mas_wm.status
		input  wire [42:0] i_tx_pcs_data,                                      //                                      i_tx_pcs_data.data
		input  wire [42:0] i_tx_mac_data,                                      //                                      i_tx_mac_data.data
		output wire [19:0] o_lavmm_xcvrif_addr,                                //                                    reconfig_xcvrif.address
		output wire [3:0]  o_lavmm_xcvrif_be,                                  //                                                   .byteenable
		output wire        o_lavmm_xcvrif_read,                                //                                                   .read
		output wire [31:0] o_lavmm_xcvrif_wdata,                               //                                                   .writedata
		output wire        o_lavmm_xcvrif_write,                               //                                                   .write
		input  wire [31:0] i_lavmm_xcvrif_rdata,                               //                                                   .readdata
		input  wire        i_lavmm_xcvrif_rdata_valid,                         //                                                   .readdatavalid
		input  wire        i_lavmm_xcvrif_waitreq,                             //                                                   .waitrequest
		output wire        o_lavmm_xcvrif_clk,                                 //                                reconfig_xcvrif_clk.clk
		output wire        o_lavmm_xcvrif_rstn,                                //                                reconfig_xcvrif_rst.reset
		output wire [19:0] o_lavmm_emac_addr,                                  //                                      reconfig_emac.address
		output wire [3:0]  o_lavmm_emac_be,                                    //                                                   .byteenable
		output wire        o_lavmm_emac_read,                                  //                                                   .read
		output wire [31:0] o_lavmm_emac_wdata,                                 //                                                   .writedata
		output wire        o_lavmm_emac_write,                                 //                                                   .write
		input  wire [31:0] i_lavmm_emac_rdata,                                 //                                                   .readdata
		input  wire        i_lavmm_emac_rdata_valid,                           //                                                   .readdatavalid
		input  wire        i_lavmm_emac_waitreq,                               //                                                   .waitrequest
		output wire        o_lavmm_emac_clk,                                   //                                  reconfig_emac_clk.clk
		output wire        o_lavmm_emac_rstn,                                  //                                  reconfig_emac_rst.reset
		output wire [19:0] o_lavmm_epcs_addr,                                  //                                      reconfig_epcs.address
		output wire [3:0]  o_lavmm_epcs_be,                                    //                                                   .byteenable
		output wire        o_lavmm_epcs_read,                                  //                                                   .read
		output wire [31:0] o_lavmm_epcs_wdata,                                 //                                                   .writedata
		output wire        o_lavmm_epcs_write,                                 //                                                   .write
		input  wire [31:0] i_lavmm_epcs_rdata,                                 //                                                   .readdata
		input  wire        i_lavmm_epcs_rdata_valid,                           //                                                   .readdatavalid
		input  wire        i_lavmm_epcs_waitreq,                               //                                                   .waitrequest
		output wire        o_lavmm_epcs_clk,                                   //                                  reconfig_epcs_clk.clk
		output wire        o_lavmm_epcs_rstn,                                  //                                  reconfig_epcs_rst.reset
		output wire [19:0] o_lavmm_fec_addr,                                   //                                       reconfig_fec.address
		output wire [3:0]  o_lavmm_fec_be,                                     //                                                   .byteenable
		output wire        o_lavmm_fec_read,                                   //                                                   .read
		output wire [31:0] o_lavmm_fec_wdata,                                  //                                                   .writedata
		output wire        o_lavmm_fec_write,                                  //                                                   .write
		input  wire [31:0] i_lavmm_fec_rdata,                                  //                                                   .readdata
		input  wire        i_lavmm_fec_rdata_valid,                            //                                                   .readdatavalid
		input  wire        i_lavmm_fec_waitreq,                                //                                                   .waitrequest
		output wire        o_lavmm_fec_clk,                                    //                                   reconfig_fec_clk.clk
		output wire        o_lavmm_fec_rstn,                                   //                                   reconfig_fec_rst.reset
		output wire [19:0] o_lavmm_ux_addr,                                    //                                        reconfig_ux.address
		output wire [3:0]  o_lavmm_ux_be,                                      //                                                   .byteenable
		output wire        o_lavmm_ux_read,                                    //                                                   .read
		output wire [31:0] o_lavmm_ux_wdata,                                   //                                                   .writedata
		output wire        o_lavmm_ux_write,                                   //                                                   .write
		input  wire [31:0] i_lavmm_ux_rdata,                                   //                                                   .readdata
		input  wire        i_lavmm_ux_rdata_valid,                             //                                                   .readdatavalid
		input  wire        i_lavmm_ux_waitreq,                                 //                                                   .waitrequest
		output wire        o_lavmm_ux_clk,                                     //                                    reconfig_ux_clk.clk
		output wire        o_lavmm_ux_rstn,                                    //                                    reconfig_ux_rst.reset
		input  wire [10:0] i_ptp_tx_data,                                      //                                      i_ptp_tx_data.data
		output wire [9:0]  o_ch_ptp_rx_data,                                   //                                   o_ch_ptp_rx_data.data
		output wire [79:0] sm_pld_tx_demux_0_o_pcie,                           //                           sm_pld_tx_demux_0_o_pcie.data
		input  wire        sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp, // sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp.clk
		input  wire        sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp, // sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp.clk
		input  wire [79:0] sm_pld_rx_mux_0_i_pcie,                             //                             sm_pld_rx_mux_0_i_pcie.data
		input  wire        sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie,       //       sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie.clk
		input  wire        sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie,       //       sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie.clk
		input  wire [79:0] sm_pld_rx_mux_0_i_pcie_bond,                        //                        sm_pld_rx_mux_0_i_pcie_bond.data
		input  wire        sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top,   //   sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top.clk
		input  wire        sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top,   //   sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top.clk
		output wire [2:0]  k_user_rx_clk1_c0c1c2_sel,                          //                          k_user_rx_clk1_c0c1c2_sel.data
		output wire [2:0]  k_user_rx_clk2_c0c1c2_sel,                          //                          k_user_rx_clk2_c0c1c2_sel.data
		output wire [2:0]  k_user_tx_clk1_c0c1c2_sel,                          //                          k_user_tx_clk1_c0c1c2_sel.data
		output wire [2:0]  k_user_tx_clk2_c0c1c2_sel,                          //                          k_user_tx_clk2_c0c1c2_sel.data
		input  wire        i_ss_user_rx_clk1_clk,                              //                              i_ss_user_rx_clk1_clk.clk
		input  wire        i_ss_user_rx_clk2_clk,                              //                              i_ss_user_rx_clk2_clk.clk
		input  wire        i_ss_user_tx_clk1_clk,                              //                              i_ss_user_tx_clk1_clk.clk
		input  wire        i_ss_user_tx_clk2_clk,                              //                              i_ss_user_tx_clk2_clk.clk
		input  wire [42:0] i_ch_muxed_rx_data,                                 //                                 i_ch_muxed_rx_data.data
		output wire [2:0]  o_deskew_rx_source_sel                              //                             o_deskew_rx_source_sel.data
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (ch_pldif_l_tx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_duplex_mode_atom != "DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_fifo_mode_atom != "TX_FIFO_MODE_PHASE_COMP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_fifo_mode_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_fifo_width_atom != "TX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_fifo_width_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_fifo_mode_atom != "RX_FIFO_MODE_PHASE_COMP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_fifo_mode_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_fifo_width_atom != "RX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_fifo_width_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_clkout1_divider_atom != "TX_CLKOUT1_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_clkout1_divider_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_clkout2_divider_atom != "TX_CLKOUT2_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_clkout2_divider_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_clkout1_divider_atom != "RX_CLKOUT1_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_clkout1_divider_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_clkout2_divider_atom != "RX_CLKOUT2_DIVIDER_DIV1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_clkout2_divider_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_dr_enabled_atom != "DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_ptp_enable_atom != "PTP_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_ptp_enable_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_user1_clk_dynamic_mux_atom != "TX_USER1_CLK_DYNAMIC_MUX_UX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_user1_clk_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_user2_clk_dynamic_mux_atom != "TX_USER2_CLK_DYNAMIC_MUX_UX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_user2_clk_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_user1_clk_dynamic_mux_atom != "RX_USER1_CLK_DYNAMIC_MUX_UX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_user1_clk_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_user2_clk_dynamic_mux_atom != "RX_USER2_CLK_DYNAMIC_MUX_UX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_user2_clk_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_sup_mode_atom != "SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_sup_mode_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_mac_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_mac_en_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_pld_channel_identifier_atom != "PLD_CHANNEL_IDENTIFIER_PHIP")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_pld_channel_identifier_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_rx_fifo_wr_clk_hz_atom != 36'b000000010001111000011010001100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_rx_fifo_wr_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_tx_fifo_rd_clk_hz_atom != 36'b000000010001111000011010001100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_tx_fifo_rd_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_dyn_mux_atom != "RX_DYN_MUX_XCVRIF")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_dyn_mux_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_bond_location_atom != "TX_BOND_LOCATION_FIRST")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_bond_location_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_bond_location_atom != "RX_BOND_LOCATION_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_bond_location_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_ehip_lb_tx_rx_atom != "EHIP_LB_TX_RX_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_ehip_lb_tx_rx_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_ehip_lb_txmac_rx_atom != "EHIP_LB_TXMAC_RX_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_ehip_lb_txmac_rx_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_rx_pmadir_singlewidth_en_atom != "RX_PMADIR_SINGLEWIDTH_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_rx_pmadir_singlewidth_en_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_tx_pmadir_singlewidth_en_atom != "TX_PMADIR_SINGLEWIDTH_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_tx_pmadir_singlewidth_en_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_ehip_lb_txpcs_rx_atom != "EHIP_LB_TXPCS_RX_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_ehip_lb_txpcs_rx_atom_check ( .error(1'b1) );
		end
		if (ch_pcs_l_tx_bond_size_atom != "TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pcs_l_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch_pcs_l_rx_bond_size_atom != "RX_BOND_SIZE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pcs_l_rx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch_vc_rx_pldif_wm_en_atom != "VC_RX_PLDIF_WM_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_vc_rx_pldif_wm_en_atom_check ( .error(1'b1) );
		end
		if (ch_pldif_l_stmux_tx_demux_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_stmux_tx_demux_sel_check ( .error(1'b1) );
		end
		if (ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel_check ( .error(1'b1) );
		end
		if (ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel_check ( .error(1'b1) );
		end
		if (ch_pldif_l_stmux_rx_mux_sel != "SEL_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pldif_l_stmux_rx_mux_sel_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_preloaded_hardware_configs != "PCIE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_preloaded_hardware_configs_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_preloaded_hardware_configs != "PCIE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_preloaded_hardware_configs_check ( .error(1'b1) );
		end
	endgenerate

	system_intel_pcie_gts_0_pldif_hal_2100_uhebp5y #(
		.ch_pldif_l_tx_en_atom                    ("TRUE"),
		.ch_pldif_l_rx_en_atom                    ("TRUE"),
		.ch_pldif_l_duplex_mode_atom              ("DUPLEX_MODE_DUPLEX"),
		.ch_pldif_l_tx_fifo_mode_atom             ("TX_FIFO_MODE_PHASE_COMP"),
		.ch_pldif_l_tx_fifo_width_atom            ("TX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH"),
		.ch_pldif_l_rx_fifo_mode_atom             ("RX_FIFO_MODE_PHASE_COMP"),
		.ch_pldif_l_rx_fifo_width_atom            ("RX_FIFO_WIDTH_DOUBLE_DOUBLE_WIDTH"),
		.ch_pldif_l_tx_clkout1_divider_atom       ("TX_CLKOUT1_DIVIDER_DIV1"),
		.ch_pldif_l_tx_clkout2_divider_atom       ("TX_CLKOUT2_DIVIDER_DIV1"),
		.ch_pldif_l_rx_clkout1_divider_atom       ("RX_CLKOUT1_DIVIDER_DIV1"),
		.ch_pldif_l_rx_clkout2_divider_atom       ("RX_CLKOUT2_DIVIDER_DIV1"),
		.ch_pldif_l_dr_enabled_atom               ("DR_ENABLED_DR_DISABLED"),
		.ch_pldif_l_ptp_enable_atom               ("PTP_ENABLE_DISABLE"),
		.ch_pldif_l_tx_user1_clk_dynamic_mux_atom ("TX_USER1_CLK_DYNAMIC_MUX_UX"),
		.ch_pldif_l_tx_user2_clk_dynamic_mux_atom ("TX_USER2_CLK_DYNAMIC_MUX_UX"),
		.ch_pldif_l_rx_user1_clk_dynamic_mux_atom ("RX_USER1_CLK_DYNAMIC_MUX_UX"),
		.ch_pldif_l_rx_user2_clk_dynamic_mux_atom ("RX_USER2_CLK_DYNAMIC_MUX_UX"),
		.ch_pldif_l_sup_mode_atom                 ("SUP_MODE_USER_MODE"),
		.ch_pldif_l_tx_mac_en_atom                ("FALSE"),
		.ch_pldif_l_pld_channel_identifier_atom   ("PLD_CHANNEL_IDENTIFIER_PHIP"),
		.ch_pldif_rx_fifo_wr_clk_hz_atom          (36'b000000010001111000011010001100000000),
		.ch_pldif_tx_fifo_rd_clk_hz_atom          (36'b000000010001111000011010001100000000),
		.ch_pldif_l_rx_dyn_mux_atom               ("RX_DYN_MUX_XCVRIF"),
		.ch_pldif_l_tx_bond_location_atom         ("TX_BOND_LOCATION_FIRST"),
		.ch_pldif_l_rx_bond_location_atom         ("RX_BOND_LOCATION_UNUSED"),
		.ch_pldif_l_ehip_lb_tx_rx_atom            ("EHIP_LB_TX_RX_DISABLE"),
		.ch_pldif_l_ehip_lb_txmac_rx_atom         ("EHIP_LB_TXMAC_RX_DISABLE"),
		.ch_pldif_l_rx_pmadir_singlewidth_en_atom ("RX_PMADIR_SINGLEWIDTH_EN_DISABLE"),
		.ch_pldif_l_tx_pmadir_singlewidth_en_atom ("TX_PMADIR_SINGLEWIDTH_EN_DISABLE"),
		.ch_pldif_l_ehip_lb_txpcs_rx_atom         ("EHIP_LB_TXPCS_RX_DISABLE"),
		.ch_pcs_l_tx_bond_size_atom               ("TX_BOND_SIZE_X4"),
		.ch_pcs_l_rx_bond_size_atom               ("RX_BOND_SIZE_UNUSED"),
		.ch_vc_rx_pldif_wm_en_atom                ("VC_RX_PLDIF_WM_EN_DISABLE"),
		.ch_pldif_l_stmux_tx_demux_sel            ("SEL_PCIE"),
		.ch_pldif_l_stmux_rx_fifo_wr_clk_mux_sel  ("SEL_PCIE"),
		.ch_pldif_l_stmux_tx_fifo_rd_clk_mux_sel  ("SEL_PCIE"),
		.ch_pldif_l_stmux_rx_mux_sel              ("SEL_PCIE"),
		.ch_l_xcvr_rx_preloaded_hardware_configs  ("PCIE_GEN4"),
		.ch_l_xcvr_tx_preloaded_hardware_configs  ("PCIE_GEN4")
	) pldif_hal_top (
		.i_hio_txdata                                       (i_hio_txdata),                                       //   input,   width = 80,                                       i_hio_txdata.data
		.i_hio_txdata_extra                                 (i_hio_txdata_extra),                                 //   input,   width = 10,                                 i_hio_txdata_extra.data
		.i_hio_txdata_fifo_wr_en                            (i_hio_txdata_fifo_wr_en),                            //   input,    width = 1,                            i_hio_txdata_fifo_wr_en.fifowriteenable
		.o_hio_txdata_fifo_wr_empty                         (o_hio_txdata_fifo_wr_empty),                         //  output,    width = 1,                         o_hio_txdata_fifo_wr_empty.fifowritestatus
		.o_hio_txdata_fifo_wr_pempty                        (o_hio_txdata_fifo_wr_pempty),                        //  output,    width = 1,                        o_hio_txdata_fifo_wr_pempty.fifowritestatus
		.o_hio_txdata_fifo_wr_full                          (o_hio_txdata_fifo_wr_full),                          //  output,    width = 1,                          o_hio_txdata_fifo_wr_full.fifowritestatus
		.o_hio_txdata_fifo_wr_pfull                         (o_hio_txdata_fifo_wr_pfull),                         //  output,    width = 1,                         o_hio_txdata_fifo_wr_pfull.fifowritestatus
		.o_hio_rxdata                                       (o_hio_rxdata),                                       //  output,   width = 80,                                       o_hio_rxdata.data
		.o_hio_rxdata_extra                                 (o_hio_rxdata_extra),                                 //  output,   width = 10,                                 o_hio_rxdata_extra.data
		.o_hio_rxdata_fifo_rd_empty                         (o_hio_rxdata_fifo_rd_empty),                         //  output,    width = 1,                         o_hio_rxdata_fifo_rd_empty.fiforeadenable
		.o_hio_rxdata_fifo_rd_pempty                        (o_hio_rxdata_fifo_rd_pempty),                        //  output,    width = 1,                        o_hio_rxdata_fifo_rd_pempty.fiforeadstatus
		.o_hio_rxdata_fifo_rd_full                          (o_hio_rxdata_fifo_rd_full),                          //  output,    width = 1,                          o_hio_rxdata_fifo_rd_full.fiforeadstatus
		.o_hio_rxdata_fifo_rd_pfull                         (o_hio_rxdata_fifo_rd_pfull),                         //  output,    width = 1,                         o_hio_rxdata_fifo_rd_pfull.fiforeadstatus
		.i_hio_rxdata_fifo_rd_en                            (i_hio_rxdata_fifo_rd_en),                            //   input,    width = 1,                            i_hio_rxdata_fifo_rd_en.fiforeadstatus
		.i_hio_ptp_rst_n                                    (i_hio_ptp_rst_n),                                    //   input,    width = 1,                                    i_hio_ptp_rst_n.data
		.i_hio_ehip_rx_rst_n                                (i_hio_ehip_rx_rst_n),                                //   input,    width = 1,                                i_hio_ehip_rx_rst_n.data
		.i_hio_ehip_tx_rst_n                                (i_hio_ehip_tx_rst_n),                                //   input,    width = 1,                                i_hio_ehip_tx_rst_n.data
		.i_hio_ehip_signal_ok                               (i_hio_ehip_signal_ok),                               //   input,    width = 1,                               i_hio_ehip_signal_ok.data
		.i_hio_sfreeze_2_r03f_rx_mac_srfz_n                 (i_hio_sfreeze_2_r03f_rx_mac_srfz_n),                 //   input,    width = 1,                 i_hio_sfreeze_2_r03f_rx_mac_srfz_n.data
		.i_hio_sfreeze_3_c2f_tx_deskew_srfz_n               (i_hio_sfreeze_3_c2f_tx_deskew_srfz_n),               //   input,    width = 1,               i_hio_sfreeze_3_c2f_tx_deskew_srfz_n.data
		.i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n                 (i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n),                 //   input,    width = 1,                 i_hio_t03f_sfreeze_1_tx_pcs_sfrz_n.data
		.o_hio_rstepcs_rx_pcs_fully_aligned                 (o_hio_rstepcs_rx_pcs_fully_aligned),                 //  output,    width = 1,                 o_hio_rstepcs_rx_pcs_fully_aligned.status
		.i_hio_rstfec_fec_rx_rst_n                          (i_hio_rstfec_fec_rx_rst_n),                          //   input,    width = 1,                          i_hio_rstfec_fec_rx_rst_n.data
		.i_hio_rstfec_fec_tx_rst_n                          (i_hio_rstfec_fec_tx_rst_n),                          //   input,    width = 1,                          i_hio_rstfec_fec_tx_rst_n.data
		.i_hio_rstfec_fec_csr_ret                           (i_hio_rstfec_fec_csr_ret),                           //   input,    width = 1,                           i_hio_rstfec_fec_csr_ret.data
		.o_hio_rstfec_fec_rx_rdy_n                          (o_hio_rstfec_fec_rx_rdy_n),                          //  output,    width = 1,                          o_hio_rstfec_fec_rx_rdy_n.status
		.i_hio_rstfec_rx_fec_sfrz_n                         (i_hio_rstfec_rx_fec_sfrz_n),                         //   input,    width = 1,                         i_hio_rstfec_rx_fec_sfrz_n.data
		.i_hio_rstfec_tx_fec_sfrz_n                         (i_hio_rstfec_tx_fec_sfrz_n),                         //   input,    width = 1,                         i_hio_rstfec_tx_fec_sfrz_n.data
		.i_hio_rstxcvrif_xcvrif_rx_rst_n                    (i_hio_rstxcvrif_xcvrif_rx_rst_n),                    //   input,    width = 1,                    i_hio_rstxcvrif_xcvrif_rx_rst_n.data
		.i_hio_rstxcvrif_xcvrif_tx_rst_n                    (i_hio_rstxcvrif_xcvrif_tx_rst_n),                    //   input,    width = 1,                    i_hio_rstxcvrif_xcvrif_tx_rst_n.data
		.i_hio_rstxcvrif_xcvrif_signal_ok                   (i_hio_rstxcvrif_xcvrif_signal_ok),                   //   input,    width = 1,                   i_hio_rstxcvrif_xcvrif_signal_ok.data
		.i_hio_rstxcvrif_rx_xcvrif_sfrz_n                   (i_hio_rstxcvrif_rx_xcvrif_sfrz_n),                   //   input,    width = 1,                   i_hio_rstxcvrif_rx_xcvrif_sfrz_n.data
		.i_hio_rstxcvrif_tx_xcvrif_sfrz_n                   (i_hio_rstxcvrif_tx_xcvrif_sfrz_n),                   //   input,    width = 1,                   i_hio_rstxcvrif_tx_xcvrif_sfrz_n.data
		.i_hio_rst_pld_clrhip                               (i_hio_rst_pld_clrhip),                               //   input,    width = 1,                               i_hio_rst_pld_clrhip.data
		.i_hio_rst_pld_clrpcs                               (i_hio_rst_pld_clrpcs),                               //   input,    width = 1,                               i_hio_rst_pld_clrpcs.data
		.i_hio_rst_pld_perstn                               (i_hio_rst_pld_perstn),                               //   input,    width = 1,                               i_hio_rst_pld_perstn.data
		.i_hio_rst_pld_ready                                (i_hio_rst_pld_ready),                                //   input,    width = 1,                                i_hio_rst_pld_ready.status
		.i_hio_rst_pld_adapter_rx_pld_rst_n                 (i_hio_rst_pld_adapter_rx_pld_rst_n),                 //   input,    width = 1,                 i_hio_rst_pld_adapter_rx_pld_rst_n.data
		.i_hio_rst_pld_adapter_tx_pld_rst_n                 (i_hio_rst_pld_adapter_tx_pld_rst_n),                 //   input,    width = 1,                 i_hio_rst_pld_adapter_tx_pld_rst_n.data
		.i_hio_rst_ux_rx_pma_rst_n                          (i_hio_rst_ux_rx_pma_rst_n),                          //   input,    width = 1,                          i_hio_rst_ux_rx_pma_rst_n.data
		.i_hio_rst_ux_rx_sfrz                               (i_hio_rst_ux_rx_sfrz),                               //   input,    width = 1,                               i_hio_rst_ux_rx_sfrz.data
		.i_hio_rst_ux_tx_pma_rst_n                          (i_hio_rst_ux_tx_pma_rst_n),                          //   input,    width = 1,                          i_hio_rst_ux_tx_pma_rst_n.data
		.o_hio_rst_flux0_cpi_cmn_busy                       (o_hio_rst_flux0_cpi_cmn_busy),                       //  output,    width = 1,                       o_hio_rst_flux0_cpi_cmn_busy.status
		.o_hio_rst_oflux_rx_srds_rdy                        (o_hio_rst_oflux_rx_srds_rdy),                        //  output,    width = 1,                        o_hio_rst_oflux_rx_srds_rdy.status
		.o_hio_rst_ux_all_synthlockstatus                   (o_hio_rst_ux_all_synthlockstatus),                   //  output,    width = 1,                   o_hio_rst_ux_all_synthlockstatus.status
		.o_hio_rst_ux_octl_pcs_rxstatus                     (o_hio_rst_ux_octl_pcs_rxstatus),                     //  output,    width = 1,                     o_hio_rst_ux_octl_pcs_rxstatus.status
		.o_hio_rst_ux_octl_pcs_txstatus                     (o_hio_rst_ux_octl_pcs_txstatus),                     //  output,    width = 1,                     o_hio_rst_ux_octl_pcs_txstatus.status
		.o_hio_rst_ux_rxcdrlock2data                        (o_hio_rst_ux_rxcdrlock2data),                        //  output,    width = 1,                        o_hio_rst_ux_rxcdrlock2data.data
		.o_hio_rst_ux_rxcdrlockstatus                       (o_hio_rst_ux_rxcdrlockstatus),                       //  output,    width = 1,                       o_hio_rst_ux_rxcdrlockstatus.status
		.o_ss_ehip_rx_rst_n                                 (o_ss_ehip_rx_rst_n),                                 //  output,    width = 1,                                 o_ss_ehip_rx_rst_n.data
		.o_ss_ehip_tx_rst_n                                 (o_ss_ehip_tx_rst_n),                                 //  output,    width = 1,                                 o_ss_ehip_tx_rst_n.data
		.o_ss_ehip_signal_ok                                (o_ss_ehip_signal_ok),                                //  output,    width = 1,                                o_ss_ehip_signal_ok.data
		.o_ss_sfreeze_2_r03f_rx_mac_srfz_n                  (o_ss_sfreeze_2_r03f_rx_mac_srfz_n),                  //  output,    width = 1,                  o_ss_sfreeze_2_r03f_rx_mac_srfz_n.data
		.o_ss_sfreeze_3_c2f_tx_deskew_srfz_n                (o_ss_sfreeze_3_c2f_tx_deskew_srfz_n),                //  output,    width = 1,                o_ss_sfreeze_3_c2f_tx_deskew_srfz_n.data
		.i_ss_rstepcs_rx_pcs_fully_aligned                  (i_ss_rstepcs_rx_pcs_fully_aligned),                  //   input,    width = 1,                  i_ss_rstepcs_rx_pcs_fully_aligned.status
		.o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n                  (o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n),                  //  output,    width = 1,                  o_ss_t03f_sfreeze_1_tx_pcs_sfrz_n.data
		.o_ss_rstfec_fec_rx_rst_n                           (o_ss_rstfec_fec_rx_rst_n),                           //  output,    width = 1,                           o_ss_rstfec_fec_rx_rst_n.data
		.o_ss_rstfec_fec_tx_rst_n                           (o_ss_rstfec_fec_tx_rst_n),                           //  output,    width = 1,                           o_ss_rstfec_fec_tx_rst_n.data
		.o_ss_rstfec_fec_csr_ret                            (o_ss_rstfec_fec_csr_ret),                            //  output,    width = 1,                            o_ss_rstfec_fec_csr_ret.data
		.i_ss_rstfec_fec_rx_rdy_n                           (i_ss_rstfec_fec_rx_rdy_n),                           //   input,    width = 1,                           i_ss_rstfec_fec_rx_rdy_n.status
		.o_ss_rstfec_rx_fec_sfrz_n                          (o_ss_rstfec_rx_fec_sfrz_n),                          //  output,    width = 1,                          o_ss_rstfec_rx_fec_sfrz_n.data
		.o_ss_rstfec_tx_fec_sfrz_n                          (o_ss_rstfec_tx_fec_sfrz_n),                          //  output,    width = 1,                          o_ss_rstfec_tx_fec_sfrz_n.data
		.o_ss_rstxcvrif_xcvrif_rx_rst_n                     (o_ss_rstxcvrif_xcvrif_rx_rst_n),                     //  output,    width = 1,                     o_ss_rstxcvrif_xcvrif_rx_rst_n.data
		.o_ss_rstxcvrif_xcvrif_tx_rst_n                     (o_ss_rstxcvrif_xcvrif_tx_rst_n),                     //  output,    width = 1,                     o_ss_rstxcvrif_xcvrif_tx_rst_n.data
		.o_ss_rstxcvrif_xcvrif_signal_ok                    (o_ss_rstxcvrif_xcvrif_signal_ok),                    //  output,    width = 1,                    o_ss_rstxcvrif_xcvrif_signal_ok.data
		.o_ss_rstxcvrif_rx_xcvrif_sfrz_n                    (o_ss_rstxcvrif_rx_xcvrif_sfrz_n),                    //  output,    width = 1,                    o_ss_rstxcvrif_rx_xcvrif_sfrz_n.data
		.o_ss_rstxcvrif_tx_xcvrif_sfrz_n                    (o_ss_rstxcvrif_tx_xcvrif_sfrz_n),                    //  output,    width = 1,                    o_ss_rstxcvrif_tx_xcvrif_sfrz_n.data
		.o_ss_rst_ux_rx_pma_rst_n                           (o_ss_rst_ux_rx_pma_rst_n),                           //  output,    width = 1,                           o_ss_rst_ux_rx_pma_rst_n.data
		.o_ss_rst_ux_rx_sfrz                                (o_ss_rst_ux_rx_sfrz),                                //  output,    width = 1,                                o_ss_rst_ux_rx_sfrz.data
		.o_ss_rst_ux_tx_pma_rst_n                           (o_ss_rst_ux_tx_pma_rst_n),                           //  output,    width = 1,                           o_ss_rst_ux_tx_pma_rst_n.data
		.i_ss_rst_flux0_cpi_cmn_busy                        (i_ss_rst_flux0_cpi_cmn_busy),                        //   input,    width = 1,                        i_ss_rst_flux0_cpi_cmn_busy.status
		.i_ss_rst_oflux_rx_srds_rdy                         (i_ss_rst_oflux_rx_srds_rdy),                         //   input,    width = 1,                         i_ss_rst_oflux_rx_srds_rdy.status
		.i_ss_rst_ux_all_synthlockstatus                    (i_ss_rst_ux_all_synthlockstatus),                    //   input,    width = 1,                    i_ss_rst_ux_all_synthlockstatus.status
		.i_ss_rst_ux_octl_pcs_rxstatus                      (i_ss_rst_ux_octl_pcs_rxstatus),                      //   input,    width = 1,                      i_ss_rst_ux_octl_pcs_rxstatus.status
		.i_ss_rst_ux_octl_pcs_txstatus                      (i_ss_rst_ux_octl_pcs_txstatus),                      //   input,    width = 1,                      i_ss_rst_ux_octl_pcs_txstatus.status
		.i_ss_rst_ux_rxcdrlock2data                         (i_ss_rst_ux_rxcdrlock2data),                         //   input,    width = 1,                         i_ss_rst_ux_rxcdrlock2data.data
		.i_ss_rst_ux_rxcdrlockstatus                        (i_ss_rst_ux_rxcdrlockstatus),                        //   input,    width = 1,                        i_ss_rst_ux_rxcdrlockstatus.status
		.i_hio_pld_reset_clk_row                            (i_hio_pld_reset_clk_row),                            //   input,    width = 1,                            i_hio_pld_reset_clk_row.status
		.i_ss_eth_fec_rx_async                              (i_ss_eth_fec_rx_async),                              //   input,   width = 12,                                        asyncdata_0.data
		.i_ss_eth_fec_rx_direct                             (i_ss_eth_fec_rx_direct),                             //   input,    width = 1,                                        asyncdata_1.data
		.o_ss_eth_fec_tx_async                              (o_ss_eth_fec_tx_async),                              //  output,    width = 7,                                        asyncdata_2.data
		.o_ss_eth_fec_tx_direct                             (o_ss_eth_fec_tx_direct),                             //  output,    width = 1,                                        asyncdata_3.data
		.i_ss_eth_mac_rx_async                              (i_ss_eth_mac_rx_async),                              //   input,   width = 14,                                        asyncdata_4.data
		.i_ss_eth_mac_rx_direct                             (i_ss_eth_mac_rx_direct),                             //   input,    width = 1,                                        asyncdata_5.data
		.o_ss_eth_mac_tx_async                              (o_ss_eth_mac_tx_async),                              //  output,   width = 14,                                        asyncdata_6.data
		.o_ss_eth_mac_tx_direct                             (o_ss_eth_mac_tx_direct),                             //  output,    width = 1,                                        asyncdata_7.data
		.i_ss_eth_pcs_rx_async                              (i_ss_eth_pcs_rx_async),                              //   input,   width = 14,                                        asyncdata_8.data
		.i_ss_eth_pcs_rx_direct                             (i_ss_eth_pcs_rx_direct),                             //   input,    width = 1,                                        asyncdata_9.data
		.o_ss_eth_pcs_tx_async                              (o_ss_eth_pcs_tx_async),                              //  output,    width = 8,                                       asyncdata_10.data
		.o_ss_eth_pcs_tx_direct                             (o_ss_eth_pcs_tx_direct),                             //  output,    width = 1,                                       asyncdata_11.data
		.i_ss_eth_xcvrif_rx_async                           (i_ss_eth_xcvrif_rx_async),                           //   input,   width = 14,                                       asyncdata_12.data
		.i_ss_eth_xcvrif_rx_direct                          (i_ss_eth_xcvrif_rx_direct),                          //   input,    width = 1,                                       asyncdata_13.data
		.o_ss_eth_xcvrif_tx_async                           (o_ss_eth_xcvrif_tx_async),                           //  output,    width = 7,                                       asyncdata_14.data
		.o_ss_eth_xcvrif_tx_direct                          (o_ss_eth_xcvrif_tx_direct),                          //  output,    width = 1,                                       asyncdata_15.data
		.i_ss_pcie_ctrl_rx_async                            (i_ss_pcie_ctrl_rx_async),                            //   input,   width = 88,                                       asyncdata_16.data
		.i_ss_pcie_ctrl_rx_direct                           (i_ss_pcie_ctrl_rx_direct),                           //   input,    width = 8,                                       asyncdata_17.data
		.o_ss_uxquad_async                                  (o_ss_uxquad_async),                                  //  output,   width = 80,                                       asyncdata_20.data
		.o_ss_uxquad_async_pcie_mux                         (o_ss_uxquad_async_pcie_mux),                         //  output,   width = 80,                                       asyncdata_21.data
		.i_ss_uxquad_async                                  (i_ss_uxquad_async),                                  //   input,   width = 50,                                       asyncdata_22.data
		.i_hio_uxquad_async                                 (i_hio_uxquad_async),                                 //   input,   width = 80,                                       asyncdata_23.data
		.i_hio_uxquad_async_pcie_mux                        (i_hio_uxquad_async_pcie_mux),                        //   input,   width = 80,                                       asyncdata_24.data
		.o_hio_uxquad_async                                 (o_hio_uxquad_async),                                 //  output,   width = 50,                                       asyncdata_25.data
		.i_hio_txdata_async                                 (i_hio_txdata_async),                                 //   input,  width = 100,                                       asyncdata_26.data
		.i_hio_txdata_direct                                (i_hio_txdata_direct),                                //   input,   width = 10,                                       asyncdata_27.data
		.o_hio_rxdata_async                                 (o_hio_rxdata_async),                                 //  output,  width = 100,                                       asyncdata_28.data
		.o_hio_rxdata_direct                                (o_hio_rxdata_direct),                                //  output,   width = 10,                                       asyncdata_29.data
		.o_hio_lavmm_rdata                                  (o_hio_lavmm_rdata),                                  //  output,   width = 32,                                     reconfig_lavmm.readdata
		.o_hio_lavmm_rdata_valid                            (o_hio_lavmm_rdata_valid),                            //  output,    width = 1,                                                   .readdatavalid
		.o_hio_lavmm_waitreq                                (o_hio_lavmm_waitreq),                                //  output,    width = 1,                                                   .waitrequest
		.i_hio_lavmm_addr                                   (i_hio_lavmm_addr),                                   //   input,   width = 21,                                                   .address
		.i_hio_lavmm_be                                     (i_hio_lavmm_be),                                     //   input,    width = 4,                                                   .byteenable
		.i_hio_lavmm_read                                   (i_hio_lavmm_read),                                   //   input,    width = 1,                                                   .read
		.i_hio_lavmm_wdata                                  (i_hio_lavmm_wdata),                                  //   input,   width = 32,                                                   .writedata
		.i_hio_lavmm_write                                  (i_hio_lavmm_write),                                  //   input,    width = 1,                                                   .write
		.i_hio_lavmm_clk                                    (i_hio_lavmm_clk),                                    //   input,    width = 1,                                 reconfig_lavmm_clk.clk
		.i_hio_lavmm_rstn                                   (i_hio_lavmm_rstn),                                   //   input,    width = 1,                                 reconfig_lavmm_rst.reset
		.i_ss_lavmm_pcie_rdata                              (i_ss_lavmm_pcie_rdata),                              //   input,   width = 32,                                      reconfig_pcie.readdata
		.i_ss_lavmm_pcie_rdata_valid                        (i_ss_lavmm_pcie_rdata_valid),                        //   input,    width = 1,                                                   .readdatavalid
		.i_ss_lavmm_pcie_waitreq                            (i_ss_lavmm_pcie_waitreq),                            //   input,    width = 1,                                                   .waitrequest
		.o_ss_lavmm_pcie_addr                               (o_ss_lavmm_pcie_addr),                               //  output,   width = 17,                                                   .address
		.o_ss_lavmm_pcie_be                                 (o_ss_lavmm_pcie_be),                                 //  output,    width = 4,                                                   .byteenable
		.o_ss_lavmm_pcie_read                               (o_ss_lavmm_pcie_read),                               //  output,    width = 1,                                                   .read
		.o_ss_lavmm_pcie_wdata                              (o_ss_lavmm_pcie_wdata),                              //  output,   width = 32,                                                   .writedata
		.o_ss_lavmm_pcie_write                              (o_ss_lavmm_pcie_write),                              //  output,    width = 1,                                                   .write
		.o_ss_lavmm_pcie_clk                                (o_ss_lavmm_pcie_clk),                                //  output,    width = 1,                                  reconfig_pcie_clk.clk
		.o_ss_lavmm_pcie_rstn                               (o_ss_lavmm_pcie_rstn),                               //  output,    width = 1,                                  reconfig_pcie_rst.reset
		.o_hio_user_rx_clk1_clk                             (o_hio_user_rx_clk1_clk),                             //  output,    width = 1,                             o_hio_user_rx_clk1_clk.clk
		.o_hio_user_rx_clk2_clk                             (o_hio_user_rx_clk2_clk),                             //  output,    width = 1,                             o_hio_user_rx_clk2_clk.clk
		.o_hio_user_tx_clk1_clk                             (o_hio_user_tx_clk1_clk),                             //  output,    width = 1,                             o_hio_user_tx_clk1_clk.clk
		.o_hio_user_tx_clk2_clk                             (o_hio_user_tx_clk2_clk),                             //  output,    width = 1,                             o_hio_user_tx_clk2_clk.clk
		.i_ux_chnl_refclk_mux                               (i_ux_chnl_refclk_mux),                               //   input,    width = 1,                               i_ux_chnl_refclk_mux.clk
		.o_hio_ux_chnl_refclk_mux                           (o_hio_ux_chnl_refclk_mux),                           //  output,    width = 1,                           o_hio_ux_chnl_refclk_mux.data
		.i_hio_pld_rx_clk_in_row_clk                        (i_hio_pld_rx_clk_in_row_clk),                        //   input,    width = 1,                        i_hio_pld_rx_clk_in_row_clk.clk
		.i_hio_pld_tx_clk_in_row_clk                        (i_hio_pld_tx_clk_in_row_clk),                        //   input,    width = 1,                        i_hio_pld_tx_clk_in_row_clk.clk
		.i_hio_det_lat_rx_dl_clk                            (i_hio_det_lat_rx_dl_clk),                            //   input,    width = 1,                            i_hio_det_lat_rx_dl_clk.clk
		.i_hio_det_lat_rx_mux_select                        (i_hio_det_lat_rx_mux_select),                        //   input,    width = 1,                        i_hio_det_lat_rx_mux_select.muxsel
		.i_hio_det_lat_rx_sclk_flop                         (i_hio_det_lat_rx_sclk_flop),                         //   input,    width = 1,                         i_hio_det_lat_rx_sclk_flop.clk
		.i_hio_det_lat_rx_sclk_gen_clk                      (i_hio_det_lat_rx_sclk_gen_clk),                      //   input,    width = 1,                      i_hio_det_lat_rx_sclk_gen_clk.clk
		.i_hio_det_lat_rx_trig_flop                         (i_hio_det_lat_rx_trig_flop),                         //   input,    width = 1,                         i_hio_det_lat_rx_trig_flop.clk
		.i_hio_det_lat_sampling_clk                         (i_hio_det_lat_sampling_clk),                         //   input,    width = 1,                         i_hio_det_lat_sampling_clk.clk
		.i_hio_det_lat_tx_dl_clk                            (i_hio_det_lat_tx_dl_clk),                            //   input,    width = 1,                            i_hio_det_lat_tx_dl_clk.clk
		.i_hio_det_lat_tx_mux_select                        (i_hio_det_lat_tx_mux_select),                        //   input,    width = 1,                        i_hio_det_lat_tx_mux_select.muxsel
		.i_hio_det_lat_tx_sclk_flop                         (i_hio_det_lat_tx_sclk_flop),                         //   input,    width = 1,                         i_hio_det_lat_tx_sclk_flop.clk
		.i_hio_det_lat_tx_sclk_gen_clk                      (i_hio_det_lat_tx_sclk_gen_clk),                      //   input,    width = 1,                      i_hio_det_lat_tx_sclk_gen_clk.clk
		.i_hio_det_lat_tx_trig_flop                         (i_hio_det_lat_tx_trig_flop),                         //   input,    width = 1,                         i_hio_det_lat_tx_trig_flop.clk
		.o_hio_det_lat_rx_async_dl_sync                     (o_hio_det_lat_rx_async_dl_sync),                     //  output,    width = 1,                     o_hio_det_lat_rx_async_dl_sync.syncsignal
		.o_hio_det_lat_rx_async_pulse                       (o_hio_det_lat_rx_async_pulse),                       //  output,    width = 1,                       o_hio_det_lat_rx_async_pulse.syncsignal
		.o_hio_det_lat_rx_async_sample_sync                 (o_hio_det_lat_rx_async_sample_sync),                 //  output,    width = 1,                 o_hio_det_lat_rx_async_sample_sync.syncsignal
		.o_hio_det_lat_rx_sclk_sample_sync                  (o_hio_det_lat_rx_sclk_sample_sync),                  //  output,    width = 1,                  o_hio_det_lat_rx_sclk_sample_sync.syncsignal
		.o_hio_det_lat_rx_trig_sample_sync                  (o_hio_det_lat_rx_trig_sample_sync),                  //  output,    width = 1,                  o_hio_det_lat_rx_trig_sample_sync.syncsignal
		.o_hio_det_lat_tx_async_dl_sync                     (o_hio_det_lat_tx_async_dl_sync),                     //  output,    width = 1,                     o_hio_det_lat_tx_async_dl_sync.syncsignal
		.o_hio_det_lat_tx_async_pulse                       (o_hio_det_lat_tx_async_pulse),                       //  output,    width = 1,                       o_hio_det_lat_tx_async_pulse.syncsignal
		.o_hio_det_lat_tx_async_sample_sync                 (o_hio_det_lat_tx_async_sample_sync),                 //  output,    width = 1,                 o_hio_det_lat_tx_async_sample_sync.syncsignal
		.o_hio_det_lat_tx_sclk_sample_sync                  (o_hio_det_lat_tx_sclk_sample_sync),                  //  output,    width = 1,                  o_hio_det_lat_tx_sclk_sample_sync.syncsignal
		.o_hio_det_lat_tx_trig_sample_sync                  (o_hio_det_lat_tx_trig_sample_sync),                  //  output,    width = 1,                  o_hio_det_lat_tx_trig_sample_sync.syncsignal
		.o_hio_xcvrif_rx_latency_pulse                      (o_hio_xcvrif_rx_latency_pulse),                      //  output,    width = 1,                      o_hio_xcvrif_rx_latency_pulse.syncsignal
		.o_hio_xcvrif_tx_latency_pulse                      (o_hio_xcvrif_tx_latency_pulse),                      //  output,    width = 1,                      o_hio_xcvrif_tx_latency_pulse.syncsignal
		.o_ss_det_lat_rx_sclk_clk                           (o_ss_det_lat_rx_sclk_clk),                           //  output,    width = 1,                           o_ss_det_lat_rx_sclk_clk.clk
		.o_ss_det_lat_rx_sclk_sync                          (o_ss_det_lat_rx_sclk_sync),                          //  output,    width = 1,                          o_ss_det_lat_rx_sclk_sync.syncsignal
		.o_ss_det_lat_tx_sclk_clk                           (o_ss_det_lat_tx_sclk_clk),                           //  output,    width = 1,                           o_ss_det_lat_tx_sclk_clk.clk
		.o_ss_det_lat_tx_sclk_sync                          (o_ss_det_lat_tx_sclk_sync),                          //  output,    width = 1,                          o_ss_det_lat_tx_sclk_sync.syncsignal
		.i_ss_det_lat_rx_async_pulse                        (i_ss_det_lat_rx_async_pulse),                        //   input,    width = 1,                        i_ss_det_lat_rx_async_pulse.syncsignal
		.i_ss_det_lat_tx_async_pulse                        (i_ss_det_lat_tx_async_pulse),                        //   input,    width = 1,                        i_ss_det_lat_tx_async_pulse.syncsignal
		.i_ss_xcvrif_rx_latency_pulse                       (i_ss_xcvrif_rx_latency_pulse),                       //   input,    width = 1,                       i_ss_xcvrif_rx_latency_pulse.syncsignal
		.i_ss_xcvrif_tx_latency_pulse                       (i_ss_xcvrif_tx_latency_pulse),                       //   input,    width = 1,                       i_ss_xcvrif_tx_latency_pulse.syncsignal
		.i_ux_tx_ch_ptr_smpl                                (i_ux_tx_ch_ptr_smpl),                                //   input,    width = 1,                                i_ux_tx_ch_ptr_smpl.syncsignal
		.o_hio_ux_tx_ch_ptr_smpl                            (o_hio_ux_tx_ch_ptr_smpl),                            //  output,    width = 1,                            o_hio_ux_tx_ch_ptr_smpl.syncsignal
		.i_deskew_rx_ch_clk                                 (i_deskew_rx_ch_clk),                                 //   input,    width = 1,                                 i_deskew_rx_ch_clk.clk
		.i_deskew_tx_ch_clk                                 (i_deskew_tx_ch_clk),                                 //   input,    width = 1,                                 i_deskew_tx_ch_clk.clk
		.o_marker_found                                     (o_marker_found),                                     //  output,    width = 1,                                     o_marker_found.status
		.i_marker_found_up                                  (i_marker_found_up),                                  //   input,    width = 1,                                  i_marker_found_up.status
		.i_marker_found_dn                                  (i_marker_found_dn),                                  //   input,    width = 1,                                  i_marker_found_dn.status
		.o_ch_pld_tx_deskewed_data                          (o_ch_pld_tx_deskewed_data),                          //  output,   width = 43,                          o_ch_pld_tx_deskewed_data.data
		.o_ch_ptp_tx_deskewed_data                          (o_ch_ptp_tx_deskewed_data),                          //  output,    width = 9,                          o_ch_ptp_tx_deskewed_data.data
		.i_ch_ptp_rx_data                                   (i_ch_ptp_rx_data),                                   //   input,    width = 8,                                   i_ch_ptp_rx_data.data
		.i_ch_tx_mac_ready                                  (i_ch_tx_mac_ready),                                  //   input,    width = 1,                                  i_ch_tx_mac_ready.status
		.i_ch_rx_mac_inframe                                (i_ch_rx_mac_inframe),                                //   input,    width = 1,                                i_ch_rx_mac_inframe.status
		.o_ch_tx_mac_valid                                  (o_ch_tx_mac_valid),                                  //  output,    width = 1,                                  o_ch_tx_mac_valid.status
		.i_ptp_rx_dsk_marker                                (i_ptp_rx_dsk_marker),                                //   input,    width = 1,                                i_ptp_rx_dsk_marker.status
		.i_ptp_mas_wm                                       (i_ptp_mas_wm),                                       //   input,    width = 1,                                       i_ptp_mas_wm.status
		.i_tx_pcs_data                                      (i_tx_pcs_data),                                      //   input,   width = 43,                                      i_tx_pcs_data.data
		.i_tx_mac_data                                      (i_tx_mac_data),                                      //   input,   width = 43,                                      i_tx_mac_data.data
		.o_lavmm_xcvrif_addr                                (o_lavmm_xcvrif_addr),                                //  output,   width = 20,                                    reconfig_xcvrif.address
		.o_lavmm_xcvrif_be                                  (o_lavmm_xcvrif_be),                                  //  output,    width = 4,                                                   .byteenable
		.o_lavmm_xcvrif_read                                (o_lavmm_xcvrif_read),                                //  output,    width = 1,                                                   .read
		.o_lavmm_xcvrif_wdata                               (o_lavmm_xcvrif_wdata),                               //  output,   width = 32,                                                   .writedata
		.o_lavmm_xcvrif_write                               (o_lavmm_xcvrif_write),                               //  output,    width = 1,                                                   .write
		.i_lavmm_xcvrif_rdata                               (i_lavmm_xcvrif_rdata),                               //   input,   width = 32,                                                   .readdata
		.i_lavmm_xcvrif_rdata_valid                         (i_lavmm_xcvrif_rdata_valid),                         //   input,    width = 1,                                                   .readdatavalid
		.i_lavmm_xcvrif_waitreq                             (i_lavmm_xcvrif_waitreq),                             //   input,    width = 1,                                                   .waitrequest
		.o_lavmm_xcvrif_clk                                 (o_lavmm_xcvrif_clk),                                 //  output,    width = 1,                                reconfig_xcvrif_clk.clk
		.o_lavmm_xcvrif_rstn                                (o_lavmm_xcvrif_rstn),                                //  output,    width = 1,                                reconfig_xcvrif_rst.reset
		.o_lavmm_emac_addr                                  (o_lavmm_emac_addr),                                  //  output,   width = 20,                                      reconfig_emac.address
		.o_lavmm_emac_be                                    (o_lavmm_emac_be),                                    //  output,    width = 4,                                                   .byteenable
		.o_lavmm_emac_read                                  (o_lavmm_emac_read),                                  //  output,    width = 1,                                                   .read
		.o_lavmm_emac_wdata                                 (o_lavmm_emac_wdata),                                 //  output,   width = 32,                                                   .writedata
		.o_lavmm_emac_write                                 (o_lavmm_emac_write),                                 //  output,    width = 1,                                                   .write
		.i_lavmm_emac_rdata                                 (i_lavmm_emac_rdata),                                 //   input,   width = 32,                                                   .readdata
		.i_lavmm_emac_rdata_valid                           (i_lavmm_emac_rdata_valid),                           //   input,    width = 1,                                                   .readdatavalid
		.i_lavmm_emac_waitreq                               (i_lavmm_emac_waitreq),                               //   input,    width = 1,                                                   .waitrequest
		.o_lavmm_emac_clk                                   (o_lavmm_emac_clk),                                   //  output,    width = 1,                                  reconfig_emac_clk.clk
		.o_lavmm_emac_rstn                                  (o_lavmm_emac_rstn),                                  //  output,    width = 1,                                  reconfig_emac_rst.reset
		.o_lavmm_epcs_addr                                  (o_lavmm_epcs_addr),                                  //  output,   width = 20,                                      reconfig_epcs.address
		.o_lavmm_epcs_be                                    (o_lavmm_epcs_be),                                    //  output,    width = 4,                                                   .byteenable
		.o_lavmm_epcs_read                                  (o_lavmm_epcs_read),                                  //  output,    width = 1,                                                   .read
		.o_lavmm_epcs_wdata                                 (o_lavmm_epcs_wdata),                                 //  output,   width = 32,                                                   .writedata
		.o_lavmm_epcs_write                                 (o_lavmm_epcs_write),                                 //  output,    width = 1,                                                   .write
		.i_lavmm_epcs_rdata                                 (i_lavmm_epcs_rdata),                                 //   input,   width = 32,                                                   .readdata
		.i_lavmm_epcs_rdata_valid                           (i_lavmm_epcs_rdata_valid),                           //   input,    width = 1,                                                   .readdatavalid
		.i_lavmm_epcs_waitreq                               (i_lavmm_epcs_waitreq),                               //   input,    width = 1,                                                   .waitrequest
		.o_lavmm_epcs_clk                                   (o_lavmm_epcs_clk),                                   //  output,    width = 1,                                  reconfig_epcs_clk.clk
		.o_lavmm_epcs_rstn                                  (o_lavmm_epcs_rstn),                                  //  output,    width = 1,                                  reconfig_epcs_rst.reset
		.o_lavmm_fec_addr                                   (o_lavmm_fec_addr),                                   //  output,   width = 20,                                       reconfig_fec.address
		.o_lavmm_fec_be                                     (o_lavmm_fec_be),                                     //  output,    width = 4,                                                   .byteenable
		.o_lavmm_fec_read                                   (o_lavmm_fec_read),                                   //  output,    width = 1,                                                   .read
		.o_lavmm_fec_wdata                                  (o_lavmm_fec_wdata),                                  //  output,   width = 32,                                                   .writedata
		.o_lavmm_fec_write                                  (o_lavmm_fec_write),                                  //  output,    width = 1,                                                   .write
		.i_lavmm_fec_rdata                                  (i_lavmm_fec_rdata),                                  //   input,   width = 32,                                                   .readdata
		.i_lavmm_fec_rdata_valid                            (i_lavmm_fec_rdata_valid),                            //   input,    width = 1,                                                   .readdatavalid
		.i_lavmm_fec_waitreq                                (i_lavmm_fec_waitreq),                                //   input,    width = 1,                                                   .waitrequest
		.o_lavmm_fec_clk                                    (o_lavmm_fec_clk),                                    //  output,    width = 1,                                   reconfig_fec_clk.clk
		.o_lavmm_fec_rstn                                   (o_lavmm_fec_rstn),                                   //  output,    width = 1,                                   reconfig_fec_rst.reset
		.o_lavmm_ux_addr                                    (o_lavmm_ux_addr),                                    //  output,   width = 20,                                        reconfig_ux.address
		.o_lavmm_ux_be                                      (o_lavmm_ux_be),                                      //  output,    width = 4,                                                   .byteenable
		.o_lavmm_ux_read                                    (o_lavmm_ux_read),                                    //  output,    width = 1,                                                   .read
		.o_lavmm_ux_wdata                                   (o_lavmm_ux_wdata),                                   //  output,   width = 32,                                                   .writedata
		.o_lavmm_ux_write                                   (o_lavmm_ux_write),                                   //  output,    width = 1,                                                   .write
		.i_lavmm_ux_rdata                                   (i_lavmm_ux_rdata),                                   //   input,   width = 32,                                                   .readdata
		.i_lavmm_ux_rdata_valid                             (i_lavmm_ux_rdata_valid),                             //   input,    width = 1,                                                   .readdatavalid
		.i_lavmm_ux_waitreq                                 (i_lavmm_ux_waitreq),                                 //   input,    width = 1,                                                   .waitrequest
		.o_lavmm_ux_clk                                     (o_lavmm_ux_clk),                                     //  output,    width = 1,                                    reconfig_ux_clk.clk
		.o_lavmm_ux_rstn                                    (o_lavmm_ux_rstn),                                    //  output,    width = 1,                                    reconfig_ux_rst.reset
		.i_ptp_tx_data                                      (i_ptp_tx_data),                                      //   input,   width = 11,                                      i_ptp_tx_data.data
		.o_ch_ptp_rx_data                                   (o_ch_ptp_rx_data),                                   //  output,   width = 10,                                   o_ch_ptp_rx_data.data
		.sm_pld_tx_demux_0_o_pcie                           (sm_pld_tx_demux_0_o_pcie),                           //  output,   width = 80,                           sm_pld_tx_demux_0_o_pcie.data
		.sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp), //   input,    width = 1, sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_eth_or_ptp.clk
		.sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp), //   input,    width = 1, sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_eth_or_ptp.clk
		.sm_pld_rx_mux_0_i_pcie                             (sm_pld_rx_mux_0_i_pcie),                             //   input,   width = 80,                             sm_pld_rx_mux_0_i_pcie.data
		.sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie       (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie),       //   input,    width = 1,       sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie.clk
		.sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie       (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie),       //   input,    width = 1,       sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie.clk
		.sm_pld_rx_mux_0_i_pcie_bond                        (sm_pld_rx_mux_0_i_pcie_bond),                        //   input,   width = 80,                        sm_pld_rx_mux_0_i_pcie_bond.data
		.sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top   (sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top),   //   input,    width = 1,   sm_hssi_pld_chnl_rx_fifo_wr_clk_mux_0_i_pcie_top.clk
		.sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top   (sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top),   //   input,    width = 1,   sm_hssi_pld_chnl_tx_fifo_rd_clk_mux_0_i_pcie_top.clk
		.k_user_rx_clk1_c0c1c2_sel                          (k_user_rx_clk1_c0c1c2_sel),                          //  output,    width = 3,                          k_user_rx_clk1_c0c1c2_sel.data
		.k_user_rx_clk2_c0c1c2_sel                          (k_user_rx_clk2_c0c1c2_sel),                          //  output,    width = 3,                          k_user_rx_clk2_c0c1c2_sel.data
		.k_user_tx_clk1_c0c1c2_sel                          (k_user_tx_clk1_c0c1c2_sel),                          //  output,    width = 3,                          k_user_tx_clk1_c0c1c2_sel.data
		.k_user_tx_clk2_c0c1c2_sel                          (k_user_tx_clk2_c0c1c2_sel),                          //  output,    width = 3,                          k_user_tx_clk2_c0c1c2_sel.data
		.i_ss_user_rx_clk1_clk                              (i_ss_user_rx_clk1_clk),                              //   input,    width = 1,                              i_ss_user_rx_clk1_clk.clk
		.i_ss_user_rx_clk2_clk                              (i_ss_user_rx_clk2_clk),                              //   input,    width = 1,                              i_ss_user_rx_clk2_clk.clk
		.i_ss_user_tx_clk1_clk                              (i_ss_user_tx_clk1_clk),                              //   input,    width = 1,                              i_ss_user_tx_clk1_clk.clk
		.i_ss_user_tx_clk2_clk                              (i_ss_user_tx_clk2_clk),                              //   input,    width = 1,                              i_ss_user_tx_clk2_clk.clk
		.i_ch_muxed_rx_data                                 (i_ch_muxed_rx_data),                                 //   input,   width = 43,                                 i_ch_muxed_rx_data.data
		.o_deskew_rx_source_sel                             (o_deskew_rx_source_sel)                              //  output,    width = 3,                             o_deskew_rx_source_sel.data
	);

endmodule
