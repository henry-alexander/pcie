// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
iOsd2bkaVS9bg0WW2jl/YCprz3KqG5rQ5p/I/GQF5j+rz6KffVW32b3X5Qqm
2RhzIX9F/FY2whxS/l40EOV4e+ggQ2zXLeSp+PRaOQmAM659fLjLL76PMEeP
SdG8AJU3ymF9W6R5qJ+eS35KQvmAEDgvpLHxsFz0rMkoC05xWiGl0S2jZZTw
uCSHQwSyjeGdFYH5EMIQTng0zMidVPbRlJabNS/SakDjT7QDlw4ogPncr0mY
jiUDtgtiJK+YoClW+QwyPXm1PgbOVh+J/aZR7w96vn0Yw86KKw1uydk4TbI5
EVNt82degjTjEKvkkDpzldvWyPeoHF8LA8PZ1lEO/Q==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hKLykUaecCLxI+p/G5Gp/++4AfnY35EiJN7dIzczJVrN6kIQZAmilAywzBp3
UPNOf1koFwDyKbch3lJkGtWNwG9l2d1s2y5g/4v6J0AUemll/BJTCM8kLMPn
ezTuJijfHmVy6daoQXOlRGQ+rcGMiruJOgpinCotZp3WSr/3ZlPPlbQnU9HZ
di3sb3ZMnse1JqmO/NtaTrQWxThT1M6zMhApT1AJzf35ibM8L7hjWhxQQh2E
HJIrEbixVVR1yMWzpXIx+lt4BICqAbjP9JNmJekCkJu+BgrECE7RCO/JeBjt
WOrCG+zPjtzeLNzOP5uwf4jAOrVzOsy7VThgTntueg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
qecXaZDbgZxZDlQr9ypVgCZ/n9YtMDEKfLUClZAPd+19nbHLwAltcifR/czW
iDmeHKHojwgl4WWVdxlPFAHT9qwUYvRMgpzdmSgUS1c2tPFxxs6DftCVNIkq
1djSg9xdSeftdakC9JL0NgvX4fjanMO56xO4H6Mo2iwoqWEwAgHeTeZrRjSr
CJ+tQHuT0SfIXZ1U/AVUW6Ks/lej39Af+IZp5xWvb/KXjA1rsQ1eb6hND3mn
TbiH3fdNF5W5iTyoZD6yyNlVlhyg7GHDGPs+Up4cdVhAIkcJQ30ScyC9vjyp
iZYs6K+9ot2J3mpcZizhfeV1LjGXLTUU2RVicToSIg==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
QgTaMJ3Zlzvh/RbIRe4qlbKwc773+Ux8868ppBI8QzB9cxg95O68W07oEbiK
1h/1bWzmdI3L0vNpr56meO5nviJGL2CMo6v4ri8MXW2+x9TPheuB+0LbH6Dz
LMbIPSwgqECqmOxp3qAIGFTYjeeMON6JUUwQF2X9poSMwCY7NKs=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
vwjQSptIAjq0qjGT3Y0GQn2l9cASHlhgJ2gCYUtO/hlUKYRLplRmbycPil0e
4IV2IX2EQFM+6FU3k8HjqgrhjNTCQI+IyHKbnUMwrvuxFJHIa6TjXZne42mZ
b4H8N39+ws9qywnz3ei8O60OUm72vF6cXXa8OGLBEZzmOYHtgu0qxDt17e5i
Nl52DJ9e1084EvkTaZglN7WYWLXF7hOU9x3ywDrWYfF//u/a8vOvNE/DdkMH
pozyKOTfVkKKn9wLnWnVeQ6gLCvcWtdFWtwhSZoQdpbVSQXOXO9AT4jr6u6y
HlF2b3DrzNl84soI3XkrDvNs72yupbR+RBy1jfsaKwwgUMHPiPBJJA/M+J9P
17wvvQyv91sjKRJP9Z3QoNmVA+hkeVsvN15mtIrDgVmqzf9dEhb33Db+JhV9
KUc9opw/BLFCn5lozexCZXpAwy3boZDKSy4h9z8MQK2x2Y1C+mtfduI9N2fM
Iaf4dPelLLQRecH2ADKNUxp+Izab6Crr


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bpCPhipLtMtX8gV1mvSTyQycC0RJYYe7k/VCURHrogv5+l1bfn1+PtPNCYpV
GYcuOeXs+i5hGNEDbDdGenUcr3BtTuw6vG8qMb9CyoxbDNdFkbtR8d61FrrE
NPr1/MY5hryzmwbb8iGrkt+OL/P5DWdqwW5cisN3rZIeF6gMELw=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
iJ3eONPCYnMoiegccTpsCdIwcMxo4aX8BLH9p2F4dL6OBIkdtNQPMbBe5vAq
IlVN9nocJmF9RaqAf+8jLaptOGwe+BFpcpRgxDiYNJLBevC2KWjDGfLoGxwH
Tomo3Jam6sf7bKbOIFlX42jHG/u3ePyB0+5kSBlaj1MMwKugRmo=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4736)
`pragma protect data_block
vwkav2L81GG6a6/ZF20ssc2hcsSwdNYHCJWrQBJqRcdTlRinJzSJlGGfM+9b
aA+f2sndXkmB99rScOIyjyDHAZp7LbQ7zU9WN2CLVqyt7of1IGYAocGZ/WPx
q1iMqAni2I9yf7aZ/s9U0irqbvlFbvFd77ui4Ie10tFJ3RPHSFXe8VRUBPIJ
bMq3+41eIB0GCTNwEEufSweMtFsWWV1JQv6Xputzzy7SY1ug8mpwKFVqr+GP
HjvkfSBn+uCWlYaqskhR9F0TuFK6GbwDO9N85pgvMy7Jz6mEVdES8RwKaG9v
SP807fpo0FKPLfl8Qg2JoUA01XBRnWrrT7OOHe+nQKK7/QIPGR7tUQqt+hx1
p9oCd8+f5VGgbOonX91XXEK9kYsuElSh5uWqxennIN/AsdukxQKSW81JWfzN
yzMmZlelzOaoOVZ5LgON8o1dcy/+gZBHNwFAzRNKIOyzKebN5pJpVqUAL8uH
b84yZk/xHMU/Y/v9PrjDvhsIdydGKwg4IFBgOWBTrgz4srojPaaE/+fA8r/R
CST0osZjvjTsx+NbuQi5MFL3er6mg1YjaJUCvVj+Imw5NmP7/gPo3dRyFYax
Xv+WJjZ7XVc6gbUzokWkj7g5zMcA7/gEF4w3xmXDBo3eN7bX7ypDXXg8hy+Z
tPmWI+5UgyggqLYXSJL3ncKUHwSZUS89lvkpjsrwaeojWHv8UXK5YzTegqbg
FTxE7xDriqDcUv8cwQGYbFGv0gpblqcTIf3w3fOwwVU2Q4FWwWtyxCFdm0Tb
PxQC3BtzaBLbA1MRhjeM5saFmNwd6PqhJhqglRcOnc0q3st7m/686mKzbkWL
hCAq3wAoWLJU0ae//FA1TFIMOINE3ok0YhlzPOGYaAzQAq84DvWXeTJaqbfe
PJwxyDC5urqM0+H+HQ3tPOugJWKe3R/oiiehfBRDtLkKasfdQ1t4C7Vm8jH1
yB7b5zj3akfo4+IGNGONt8V2TOFE44D5VYmgjmxnU34FagLJ6KN1bu+rxEcr
3O626uHrETsvleWL0zZAhdOK4TiOx1z0bpKzwHix5bF/dPsmO9txebG2i4nU
hufZend7Bg8Q0CRHrWU59QdpUY3HhYure10m/qmwxWNbukOLJMqGhqmC+PFn
vi7MFD3sljOJipiQHRMSX0yHZO6eJ4RHKJOiZJhgkEzelTBUE9eAwzqxkjVt
d0Oz/HJlcvjwttnnHyldqb0vz9yMlZ8UMlJzumtTfXzAlktdOxcab8m/F2Vy
OYSfo20kHy+NTf796q1mj45onKze2BsP+B0MeuuqprQPeRIEMwTdB5FYiszt
lmIRjVaZeCLc3HvdIr54u9XLN6Cvht6ErCIHGaXxczMRMHGxf/e7G23/mB1B
aPUARBmU/2uiPhdccAKAB8G3mCFXpywhG2iyPIS3pQ4SySarXfcXcI6Y8FXG
O62Iz9RNf45aw1WJxrHcx758mkDFHNFvwEhEzmrZeWDyQkqiWEpmzqSvPm10
gK6k2L3r+rvmQD3c6g4sku01pZ5Ve89UMNC/9mF+CP34Y9CON7AjgXDvdQDQ
KBGV1yevVPp3hGKpt5QPLoAyhzZMAuPjiN/Cvht/HtKqy4aA9wgILf+/DXz6
GEv5ejrhkhFRd02y3aVLfju+IAzEHLyxa3CWVzdzp1jw2EhbYbGRu3HCYlPi
3Fvgix16r5HXWcw4qwCTX5sJDpRC3NsVx4aPRVkWJbWrkDeG5K7cANJsbS9v
L7x6YhbDN+fsCcFChuLyKpQCpJDUbYbH6y1Elv5V6XDIWKu3KKv+a75y50zv
+yKo+cyZSuJf6RvkvODOEeGYCLQ3V3NI/cg10HjMmV4IRvHhI6RaMA3lLqva
yZnZ9b2dQ7pM5NCBOjYWCM9RqOd2Z6vZBUn/pK7i/idMMvFNKOeWW/4zZ0DE
DrPdQ5W7mv0lQ7CVh/fs/jO3mT50PEcUCfGkDnYXpOMmbDSbqf7fO967WYY7
tufULtI/2oS+BmQddUM0NW/fhSvIwyi0PHDv+njXIQocCtH52RAsdMxUF+Yx
C5K2uobIOek+DFCCYITs7j25Aaa3BxGZqCE19YDn+57MShMNj/hkkuulhiz+
eiwHJadEHtv7fDbO1+EuyXwhUtrBNdxQ0gt85/Q5QMYp9ttb/PidydPHrGn/
iL/yHSHOb4JLwCVUycpO3Yals5Wwd62cZZRIARfJM6FVmiR9bUe8Lw8mx0Rh
ISuAyFJ66qFdJxB1mbLNlL2xlv4Xatj02EZMYex9Iohipv5DRdtm13E6G7Zh
5tn7grYH2mN1QbPokU97iFcocqOmLJMLqBpYsxTp+Ulu67yBaJATU/RVnseg
CEo365CpCh8l0M7DPg+rtGXl0HeH/KffQ8qsc4lPYA8gjQXCwgGo+jeu04At
p0qlSEFp3O/gQAVjJJZ6gfmdzC7R4VYB1TcT1AHn4cbzL8/tlNlPEv44OP9R
G6qaOqiY52Vvvf43WIrGRKoD38FZ2xVqu40NrGgTfDlBlKE48jqn7n8X3ca/
/mlASBP1q3AiV4va/+smigOfzn41goKpl8xJiYf5tfSw5rypR87CxPTvLLMX
1sgVUJZHYE7reR/GVQ/jjnSqeWKUTA5sp06/yyn5/sXF5HAV0LN7iA15hWoP
2uqhBGAThXQxXwx5dWtpsp1HFT6a+IbrpTn0bkcbHUCmvCtiQuNNG6UPiksR
cb0no7VDlktK/PYFZI9u6lqOEqEoLZ1qaBJjNplfW1lWTS634t/wwh2vcp6v
OC7Op8esVbVTetGFZgxHz4QLaXVgdMW3NbDXKQRXDgV9pXA8c84yppRrtY5m
p3sk5ai91/LuerZb3rh7F785cxyi16e/cQGqa+RoNf3GH37EULpd3r21fXUE
PBrokX1DlwrQrnvZzDruKu8vL0Z3Q63Brn0b1ock25EZxOz3yMlOagA3Qfs9
EbsaGDIrpHgZ9iE+p6A9TtpDxp3C36L+KMnwl5rIrWdnbYqWFDNLSzr3yiJM
iAUDt8OuUOSEENUvpvJ7+EPiB7uwy4SIoxhwVc3URM13mfoBAoCtm1DHdWEb
q0UMaM9U4MF+VU3vlUTEQd0gHtEhlHCUrE9SuZmpc8z2TPMv3p/qj0TFxxJe
kdRajNXpJRuh5HTesSwOEjMl0Pal4CFyp7UFaKzS9PgNH87C/jKz3Z/KmoYC
X+gC0OaKomCzrp8WmksA+XnVB1AWpk1q1MCRVdlimdmTeACz4DI4q14I201C
URXkx9XGFmEpCdwc4TPlAxBCE8ZsHrJ7Ns3t3Nkp0QYeDgOxxPzJJhrC2wGo
SzySlRsuvz2UsWfISsSPkvBVbouHUQJNpogcf9XixrUJfnDXYjEBTYc1nGe9
m1XNIR8IytmUkuyo4VxkYtYja+IUWjf/EHr0o7qFlY5KsyCQ3P9wVEUnlBZC
9HXNEztI4hwE8FvmxxkKA66Yz+HWz3coABuiJDOxUft6o52IieIA13bm86hG
M9Ulvgc7WiVqUoFzLqygEcf4LQ8HppX0x4/NWUz7sxlHPhvMHS0J/Nj/J9VE
2pU4i/2DLvYyyMUUPO1EKWBYB+K4wh51p+LrizSci6jt1KgP3KpflEVGy6Eb
zrAcQul8d5lZt5np7FeSQCHjotyHL/VX6k/QzyyB0JULuWuLuh6hKp4Lpfsk
1VSin0F7jF4YGO+RpRs7qMXuEHlRDoWGoUO4PC9WrKjsEdRFGiuYYRcxjE1u
jRDDldplhkuIPmsZGFW/iZlcRFiTlzW30i+CFy9DyL2rDaEQCVl6Bs04yy3N
AdLX7ST4eiFWWxZ3Z5I0Hi3lCzxDCiIZyqKo2RBnpENE91LL9HgiAXngn++z
sGHGoZP3CSzY4RUja5kn41kmfYcbY8t9GxwiY9kW7L4qIcmJkt4dDWTpM37R
3v22su0rv6kvqqL+8IaReFEMOBnCYqdqGs0fVVeRtun1JtRGU2+Zy9SxkhgT
ObY6KJ7W8CX93wJ9wY8HDiIIVvDgnzyOJ0M74yLi5V2gvoExCF51Asjuo/hT
ZrLzvre/th8rUWCyS4axxksNSeK0n2MzMsvp5zAVStcewfxk5Qco497ckFrz
D81AKKKMmjt6bgBrN0cnq3+hFbBDnVX8WXIzCWBG1vQNQ/KHgREfyYpMFb0h
IAtI5D+EHhSjAq0VNL/UwUXPNCD4QGQ+B1K+ueh6L0xi2Wi1kTxqZTjV+9Tc
gyKZ0Ws+MSaAa8E0J8v1H0R/pMX/Gvwnl38lOzXEEeFD6eZmEHTIir6sQIIB
cIaohsGPGJccf34522bke6skkBiV8EdSbULvNUItkwDUB2ID5ZRnKJyK73sS
qgxrdaIPSgzfYxgjT2EYsEEPCkz2xom9+bj148HQAXwlmqglPU9FoI+U0qGn
d4AYXK2+UJPp+mzg3UmiLeMUtPWPad6zk6736M2OZijBOWJu1M4H5bAS3d5e
WXMw0YTUHNG7l+w2zRhFee1mD4ap2iOqgS+2gI0Y/Il9mMpDfxia85ULIATi
lPPVjJzTVVswKFgyjNcDExAN1t/Fkw9GDTqL+g6KMRRwPvD0F/eobFrf1jfx
VziQWCYA+6htU1f0+2LLJqakzS9IHSdFYm+TRZISb7Y7sE5YtYsVL0xW7any
H1/7CWyU0Ec0G63D8Y6jWV8o36vWo7TKzddcTpnqPx3Vof8GafwYMOSKPA1x
Mlxu+rSpUferJpzBeNlrZuDEcOfe8ZhS1NwrQ2QBNn1rTMTqccXz4A4/S0IF
ZCiG7rWw1oE8YKOVmE0sZt/CqUI88iL5lcnugKCSMI8FnDeGaoMpW8HPpZQ9
P6xuqHbdSeJXc8dj7GUCF9kCi54qhQGYjmZdF716BJqdmVYSIUhVnHAzPSv+
hPHPkP0OsarYIUhk1wu62LkqYeffnqEusyZsAKuf2r8z7brt9pluYSN9nf3t
8KmZuK10xOPr59JSbmSiwW4BFsCqYL338tMOa7zJQZIZxeHhhBWzgBKMNl7J
vGmyt5Xfi6AKigF6T1YfgzIiqsHILW8uhQTV07p1CvSc8nv5DarHQ7vhSTKQ
QY8Xhol7Vh8rDYkNl+Obc+/qaOT0npwL1j3FU0fo4Ae1iJNroTp8+x7YhTO5
XvtMxcBngfRv7p6f9uBEyNC4Erj0B2VmuGUA4cHPEE/q3ktND0KQH3VgohjA
Lre9ialaeVynR/V+LWs2GZmhKYrCqloDKtxzgdMppQTAPpf1260grbKsTnAM
INI1RKusuY5xvjWaU9T6bL9Z/rpscR0yxQGJVvOEGMJa7nUwJWjidwLnyQvw
dRYw9N7mp0PdKhgWcLOXzy1PUTxsIIq9pVIrI8Q29IIyNDHHxN1iRp5DI5Ed
UrJSD8B7wGucj1yPHAbTL9Qtlg5DRVVSGpCFdn8Qzh4X2LXw6+rk2A6+c7BY
aJ735OtycT5EJwNEulXTf8qfBWPURXOUTahoiis+rNLtM6H14Ztew3n9TgAz
752DQcOihKyW9vSeEwNFf9Olj1cK7hAaIFmVuC2+52n86lSCIR7c8OBQLW3R
ohVFKO5/7imSXc5MTRqJbju4cHjPqCaRok6usuER3k9xEeJH42yHQFG4vqfH
yXjYqfe0fcTlOP9l8CuXw1elYOcejtNYNrNEnHf/ZC1cElzgei3DSzu85irI
DfyT7I6Z5StOeNpjAXUIe+ICQCSd93Mdlc5lnYBmwYW33sUbYdymxWcexNc9
fydN49pRQHBrY9sl42NSBa/NNgbQLq9CXFdVreakXVdHZh57JuL2x1Lv7zgA
82tDWzUnSekKik3NYUiDcbLy/Ee5qQQJFaR/FHUijZZAM9iq7vlw2P+Zm378
7qUrIw01iyup4Vi7P4nh9IClaMGdPR6JFaLRB9sX17z6hapCoQ9NsmohCZFz
7BZJD2OjeIIP4oW4AZhImD/8wr51yd/kQZDToMtIMHhKh3w3Hq+vlyQcoVJo
kSwp7LVsAcCHbKyM/l+VQF+CmyRE3nfLWhKN37sEJ8dbKcfOynt9si2qCcRA
1XLgWJUNmmQ1IDxFZlyhu5S9+THgWMJmwnu9kAXPZeq2r/V0ncJhQiGY8RHR
pqLE/nFAbgCkbVVBxcJU0bvqGQmlzocbM5DtVqkSC16Tdn4pFuqUrml/prs1
UE2HCZQArIiRwC0O4S70ilmTk4NcOLHX32RsIQ0Nem9kMgBzaYSz5c6Q1V/D
zfwXVqlW2HUlkKdEqlM/FJ4Qk2U/G9ZrdCVa5sj2deBVT8HaeH2mrPXOUbJG
Dxu+xQyfqJVhDNJH1bg/aM+pI0o3G3BtUDNRpH2TViEe9DR10igxDgwGrDHn
RgdIPw7rggQq45U=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfSTpfx5CD/baKe4UO8zVCCXXMXv6UAB/AxiMk/sZbijNlpTZZWKis5gVXRLLAbkKMd9a2ZxRHMrll/2kR8yZnDUX1MB3YVDSjlQKgxokDenYx+uf0o+qpZTKvfMgEKi5OZEFLY6g2GPVpjWnTgVJ71dmFgWQL8Vv4z976ox/wM3R6PLTWrDCquR1F/QaDq2zO0ZpYoB6Io1lhvJLvpPEUT/C5oAuPogWpQVxwiNetUdeFmt9Does8k+Sc7sR08i/27JGHCWPLeUsRpaO8ZUzgpPi2mX8AxnhFj8fM95SU8PIxVdy6C617FMAxd+os5EcxLgxMmUOvYkmXhsdI81eKMUIXmspDRuegZih7N1WnYglVJJALmyslrv/KZkSwK0kW6KKHGmm9KZwdM26/NzgmWf7lOgLLlKwAVGW54HaO6eKYX2/K2KehXNp0cDsjE/CGnun6a004Rw1si0ZCxg/gHanYIINmEWVuFy4lnH2TpVQNa7efNdcXaqRgWS4VatIkPpX238W9A567gnoO1NLKv7Vc8L8KxIEAg7ex5NecWtAl39OZw6GNDBf6/HhRByO0i8WnGE18X8c94PJJnL9GEaH+okGTD9JoTb1zrdh7WEs/aNTUe33nKuf1/Ckeha9SKAtQg9vyfb0erwWxLfaBwHd/2TaoHWrGUUOZlgeGK4iH/ZdkGbRvv8mkEcxblIZF4tWWSJzeYOQpPoSZcHO3HzUtMmXPHTsjmvU50juMhQOBVA+Lm2/Q3Ll0Y3nyptKID8IdcR0d748OPhen2pT8iM"
`endif