//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O8XBX7v0Nvl7F7OOhFWb4+q5UhWMokYfG/4NSAku+8ck5rvVihJoOJElc1RQ
NtuOeSHdck9ZhSeZHAvLIhbmVH2O30ASAetgE0+UGUfggfscdY0w3upFrBGB
oYtZgvTCPr31+jn2xrA5OlfT8wzHXyhGeRhhQz2NqqaafHet+/PGgAf0CSEu
pr7V8/BSMgepltgfGehAxJFj6oCGFc2VRUCX17328JbnjSDMkZ/t/tnv8Ihp
fIFT7MmRianMDNwrnXGcbCN5muS73Iq6UM31rdtb6/IfEVpv8B/an9zVZJ79
oegv7rzuhch0GCtCgLiB7Aa2BK5S3veGq/Q4hNIIBQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lPWn0McrCB7wjoUostnOYchZ9+3wXHfPQkyaXkz0QXfCKoQWEi7rXl8gZMyG
VKLlM0eiGdms83AfDbh8g7Bn7XoKHGG2Pdqt7DnMBlx0KN+NbZXk+GlAD9HC
a6bMD9HZh4Ualsg6g6NJym7OsB2gtSdMZrRKATaCma3riSoZXpeHiY85cor8
QaQU0Q6/VY5UyUZK+bJ9E0+1ruCHhsujoL4eciRGsSwLEnb6dLUG9A/S86cM
61HTGuUki53ibdKEpN8l5JXb9BYtgrB0pGuTIKCRGj8wjDPa+Uj+bdIM+lpV
79CIwclJEWFBYOGkwrkYA+mWOj/AHkVHHf2TKocx9g==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Dx1MmrnVwcZs2oGlw0GTIPvidgVYEXlsE2+3r5IgCKiLWx69lPQ5sV9/tQMg
bMkJAsUxSTemH73Kt6UgDC6qpnLEM342BrmYwzeph2B5Dl1Wq/O2YFl4ZAEr
3iBfdE4Oqko40PI56QhiNObmySWoay3KvM5vFEnqNsDfyEQsScguRmlqPzyG
9Jk089Pgn0m1Np4xaRXmqqrJVbCItFkYLDtnCIFgAq7hpN6dCpjiwLXKmNiT
I7ETXJWdsEDHY0Bg5fl0clulYORyPi1249nuM2vUeOHL97QsqMIe4vgo4m69
2iPJkskTIHEw8IYh8iDeBpZoTM0ATU18k6DpUj+GPQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pXg4OBai8ii7MQ5YTfGswH7So0zwQJhtA3mOrPMZquwjGLduoS7mx9Qwadyz
jNTLIOyQXtFYPHC2F74WAoR4ejAttxx5KFE+XarlDg9VIWnXhg9HwQUnxhiG
9wlNtFqOyXpWy9Ge461gcVwLtK8Ye/Z1FmwLjQJYD4LiK5aqa8k=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
atJg0Qjou888gpjBJS4jupCspJLz0UjtzVQwGBqu8hedOoee28Jp8GX0lekz
tfdwFwFt06KN/HogEmQf0sXEmdY7MAk6LwYi+HNmgCeY/KY19V2MjmGgFQoH
i7Bz1F9/DOqhkkCXT20Rve85KsNGurJeZx4CR1bNsYW0pQe9KOPrV/UnZRT4
CGbPwFuVifFI3ZCgn00warSHdq8iUpqsg9ubx6ykl2/1p6rbt6nHDGnfeWhZ
n++NgyD2lBBfSaWTq0C5Hehx2sNVXMn737zukrinorHNww1C6bY4V1SDyDqk
t0jIhYxDuBzSof+8xRzIjIqr29+P2gCZYzpoD6hR2ZgmYxxzggPJn+VTGCC+
zVI7n19MAZBzm3N3z7k8OwixzCvBd2vNbyBm6UwmGnDXKFX52BFdGOKWdQSY
k5IpwPmJq0Kr5qsZb8fALS1BDhjP4CdTE/e4L4k5YLIRfWb4rjqWIQaEVJZ7
1FO5AYBUUE1YVfjtauGCEcP7sDJrgyZE


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
NJZjrgplIc51/Tgb1J1k3YtxCrI2tKnHSu8RJebeJ00cIN6OZ55YnUQl+Vrt
Bpd9tXcCOcKcHrSOEA/6isNtISrK5xTZkdPQa9C0k2Gwam+unwBDpGJjse4z
n92SSSqWntanpVBgu+f3Imo6FvFPByavGtVmm+lH8ghNNsfNb8M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
uuNjz8T6pWFEwJSqKSqdydxG6m0uciL8DEZ1PirRaWSBE3Vi6wcWPkWp92si
fkIE9f3VOnhOoBTVMnaTokcec0i4c1g/geToiq2fgLHZSMFQUWTuun2iLGZv
En7n783nQ1/Q/4sxHEAYGcYFaWLMROoz+YtUtTqO3HLXKkvmZFI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2672)
`pragma protect data_block
8aTfHBBrjOb3aWyG7XrMvySVG4SWC92iLvBnD0CYURXIwsaVJao6Pv2+E4s2
G8tpHV/C8IDxuAhaW3CMVrIyOmY7jRz0MIDrP0wnyQNAGkG9+OD/j+mCZuSy
2McsUSSeZJJgXBoK+2fbNnvmqBHx7S+bm8sTFy5+s93k5Epy4KU3m/hHIbov
fPEAGjygyXV0XgTaTzIGpaUUwzoMcYYOTOk+/kcANNiryoErChsJ+bUXJpjb
yyq6WmQADufbSynw2WFJo0enUb6ZOAP1ILjRGgKQPhTYBd/XHfywWf9It18Y
oB3wrvZKjBp4FqMnH2Gtj7G97GwV63dWahOCMzFUW/v7xZJwVNY+AEpfF8W0
045IUn6uWznvoFny2BEBDVDoxSJAuTt6o78hQAX/lBwYvT7y8YxE6Vy2aI1r
UWU+elSLO1hzh8oqmBWvr8OfumuxXhjZ4l3KcxDyxbpyxYUXER4s9lcjNQbW
qtvwto2JId8s7YIl+4XkBFTys7KgE5iuxTZQxS61EyzO1uhIFfz7Y6RPYB49
3qGhS/mUHBDfjgX/T+UihU4eMgHVM6IbIU6ChngQvxiSItETxoNic0jzy1eK
YQqye4nKe/lRZoBr9pyokgVPDI8Xj8ToqfPelp9HQ2/TUccGlq+/iPc0IQ8n
Jp3KUv0wjiOApvkE7ovpcWxFxCt7wzFPyaGv6JceEBGRLmsYGuVHXAYLJh5b
bp2rF6bWcEMyfNos11attpn4JY0luQsM9HFsXPVI0S7Cu4a8wKicr9InzJqS
JbCAoi7WQIbtsBP3f5x3C0bYGOB/BdRLkVjVtb6ZFtdAhL1jftUP/+O1biX5
K8mNeUNnPYOEUwekcmPu7M7gceKRCUQhtebe4igjjaqtsC0a90GmqZtcSWLP
/wrLXY7RJ2QDXOyK5SF4GIih4Ct6hiRFg/LD1F1O78Jjd3iotgWW6SEbMJsc
4tpcx4GV1tOpRoEOStB++VUnOPjGeM0+mUerjyq41IBMoff/a7A/olPFjgo4
tIEsj8a0U9pQZ6kOhcSxbrKpb283edVl8kilRiBLtjAkLFhBtlCJ1Lb0E5uK
+d4U7VbB7ZV5PRs44xjNF+jeot4sAlsV80IMRzbsqRYuQBgBV20xPEXng3V4
Wo7H2lDuRX1sBeRBidEtsmnR0NXlnmEY+zWRHgTPGpLwue55XvPa9MBqtDdq
EWurgdFHOyFj8j7RrjgauJeGdXcTwcEl8YRZ3qxv2yUxrvgj79NBNFOwrBLE
JUbnHY4J6y0xikxXLXTqMTanZk6Xyja3QE0ExH1RaZhBjzBx7Yz22iKvXC4u
WmDwO2x5VA3tB5DZbOJw3+H5kBCncKyDny0Uj6CBgjEV1RJLTptoyb18tm0i
jPBj6UOKeWUhGLosnuF6+Npdrkivll/avqEluFCnnGTg+k/elG2jdLKmuK3Q
Q0kzDgxfzrcUZQd+3f4ww8ejmgV4Vy9okLPIzVK+1eFZpgsyTyUbwQjk7WK9
aGZn7yG0fsIHWlC/P2EWbT1m+ZpTJRaYR7owkA71QwHOOpL+5F6XpX/22tfR
cRzYa8rHSVrjZ+sC+pU9xnRmGkkj3+epKlfYzQnvQk41rIPbFjdqwttNiLuM
ua3XP3CGI/lck8nUZSpXhqVKq0mGy0YuXnpjDRBFx3WMYK1g6huFvjBSbUfT
5VkyPMMWvsrKNeCJfjNKPoIYg5MRATFJH1VIR3kyu2uTvhr0bA0xTzqc33iG
6EOZLt0p+cxdS5pA3C9K+gzaG2yemboINLt8jyPb+OtHFIlMwuZShUzNFL1t
17q4wYJ1EMZNMq84i5l0J4SQN9tytupsTWKdliIe5eXfJmQBc3rxhmmkXf5H
wcj4OiAEX2v53konkFTJSowMakCclXlA3pa2TaJ35i0AWgP8iYOgmtD4dPhx
oEjqq0vkjWcBmbv5tjPq/TBGmLIMWGkCVup5Sw0RqQ21fWy4zMNjdjLwMdQM
GBNCCYefnK6HAg0Ijb4Ih5he5npLgZFN0cWYI/UPx8RsbJJcedREfmHYSJLS
oOEvJsqtgTAjvoN5YioQ0/D7gS2vApdv7k1FMpwa3t3TOOdyo0hkCO2pBvBH
0j4Bxfzjipqn0fSAOpN5QX6/GJX0ee9Vevugf3aTn3Kfkd7RIxLoocJ8i7bZ
rHWBLpYGhPnSQJ9vx94XUbKA8DFgCNsO5srmKndUiCCna4Vov/j1J7dQsnnS
7yhaft5FUAYtO0Fk1pgMcmzEdqnrb/+8g9CS6WvrqLZwDCVl4FLPxrbi+s6Q
RqnpRtbqKYSpK6yHYJ1K0FIWScTfm/3hWNSSicJrc2rsyocK6pFEmGF5GQBy
cbCX1PLcR5EebkLbMfh8maFcqMejjj5PwEp0otLW6toD/ctGcPOLlfbkFNpt
ChSwypxkA/EFs0SgAINm8xVn/AQiAL2inTZedntq3s44kIdadIxr1Zoy0jeF
Ec8qZjL874+0DTwfdfNpMMSVT5HLUYmg8Jvk8dmHb6gtp26foRsIAAMWex8r
ilJSUuNqQyILOMMag6hi4qTor6K8G6Bf9kJyh7nduSj2NOb99tdZh1uu15P9
F6hNIMNIOoPbn9EStMjSJZZFNWj7S7c7tjydUxMyfQzXYkjDEGq9zp/JjACG
2c+IPzHZDaYG9kQXBG+ge7G6wfL4qvTnUwv/phCQOZjYvy2J4VzchgDdq871
kD5FdehJm3hvhWDgVz1G86seEwx54uPxlmfREuhlYetCqpI6ptB6YvF7sd2Y
b+moqYVGJicQXFx2kKDhi2rYK8QHJYgXcKmz1kfKPAWE9HByAaG6QDP7GbBr
QPpJP2XAGzgEJysVkvOHrkTaVIlJpTIg1tx/bzE/aPYrDEPxzfiDoesJlcnd
9lIYsciHImLwkAB5rVxGbLuxSmtdGvUqR+5dS2Yis7eOdmFozEI64DhtNLMy
m5+WLZRf/zniyFXyhYXAiH2Jq+2vZ+WIwZxSq/hOMvEDUe93IuJwggm4ZTFv
eisVQo02ev1g0DFcrtfgC6Pl68DTMF3/K8Lt8+CQ5yrcbpExRfmB+isClQnB
sPHixmfusb+DMBs4JGEzTV0h0Mpq+NVEOe1rKwe9Osn72mehdodObgzTgu/l
T4tXM8HYP4BYb0g6ghQMsDKYO02xv63qeSE3I8B7b6n3r3iSC5dnc8BJVY5z
sR0dxAk4Hn3nKMsBUADXm9TgJnQG+1Rf4+gG8eFXlFXvupnN3bdy7LAxEq/x
kAOvSv891xNP5AVuGx5XxVQuZLqoqVqtOyVVWy2hL1pxW25gOJYMloHh7Ulh
b1x87IeKq90yNxIGvefeDEzR/cu4XEyxval/14/3lY/pSGBwjXjbwBkC782C
p6AhyXh1ox3h8C5dMKn1XN1ZhWZvENue3zVxlfdYkzbfFfaggGFQNKZwYHBL
eYqiXGGGwLtd3AqXBCdcvs8j+tJddo4onsgL1EciwyYdsRArJb+piXraIaiP
9w8FsWBNgL3+mOu8cDnQiT7Eii0gvn7E41FnmCwEstYY5rhgZNgHx8bkpmSA
XWiiEr7m8ddPFSIZYNthfXw=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+nS643waPJK2Hb51CIZ3G9lgwuyxLdENvFaC6W+4xqYH/RpF+3HubU02A1Keb02bhR3juFfjCS8v/MMbqUL1PymqfUy2v0bxLGwydxKn9UZejmzeAfhDaXe4M7KVeso3UmMp40Bil4UCUWBQt/jbzZ/P3wLclm+uWttHeaWsDcAzLXWsxwtaE6VMn6tMMiAbH8jPHcCHCy7mGbaBu+4Wnr5mENRVm5EQRNebvjGlDLPqmXTN2HZZfu1HLZurS7fKbIPEYohMW9kSqL89fMYtD38QZGUp/C5DqJ6gh2DCgqDS6lil7ws/we5vqSebiWDYDlI/Nu6GCZX8q1kAMmejqRsAlcGu03actkVKgQxJQiVfgncUSdsqarPer4m0vqCYQ207Ju5i7Sj1eoxxsODK+cJFyqtYcKqvjlMKBSHRj+pgf/U2XzU0D2WwOgkQVvjpV2HyWEE2BSS8YboiLFYHT/P1v2WU9GSrdEsp4yL5oNhyRCLnglIKXQufQaTz8CMfV3sZrok8DoZXJFyz7jTdSTZfcI7QAxNGEyEkjQZVKGqSv+5sStKbGfI/nTPJpDrx0rAQeoQ2Y/vXFPBLPWGBG4K5LGfOp8kSlHn5clCmW9RX9VKdtWGR3k54EP7WByygjMNKkM55pT7Fa084BLs6gJysu3v3CEoS3ZJ7eQDEgLy1srkrm0FYgsBrL2NUv49UYSwYUygtMbyIsMbfngi3fqBGbzQnlKYx7OmsAuhlti5XLjPkGlDEYzyEXZM8nsHgpYMRjhKW4HuaPRZYcuqbozR"
`endif