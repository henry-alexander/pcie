// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Fd5tM/yvH6PiD1OQOzpi/n7bgqaCQH+JALSWJZxr9p9kpiL3b0PESFGg68S1
gRT2/HUCXyzEirBRZb3wjQtQS3IrT0oblzAKLDeOVKi7pORtsqgAWC6yYDnR
opKFjd//L2lxunvw8iQZxa/fdYn1CsU9yi+U7cMqSn9OayyIZLQNz6uNufNR
6ng7zE1qNWRTGUlyfLUz95V02tkeBHmL8qeMvrSIzzSGV4Z7izsZtYB1D758
fRjVqHnIB/oGOO2Hpc06Y/0OoX3ywOgqBIgD7DYcC7CAq+Ua7Cpz/K0TmBS4
u3I8/bIgcD/FRF+dIZ2rWbykTQDwBm+UD45KhrZTKQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
RX5TaKcbaEZjyf5TgJQD0AzWA3LPqzZFT5BfRGUSkJV0JMpHpbR6uDB4j3Qo
Q51eeOJ2kvxcjUFplCKTP2HH6/DANSSTCzsCqWmRQ+k0NbgslhVdpb6Jm2kr
ceUhzj+TmQreVIf6o66msDvkOEktqVMETUwDDsQ+RZHVTK3L0OaF+zpA9LbT
X295ePrzgKVYsiFlOeCemomrD6RvXwGD4C4Vgp8ETW9+UfvAaU6guKH2CSC/
KskFfQ84HRA4Bh6bwIpADS4moAs00r3If3TfcSf8yBwLVkVdA/CB6D7zy3/h
FE3UVns1sJISbQM9fNkEj4Rt6Lttp0CBV+R8OrTAEA==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
lsqSMmRig3WdMrHAcTCJkhIFrSckCvsyiFvcuLziArPrdtDlXCBP1xGfKCN2
n/oLveB+gSkP6jXSPCCzbRZl/1J5SNnLOwKtzvl2FWVjnz6hyp4c/RYPpZsX
djzguQAdFSh2U7jNBSeTV0SRyGX+OKErYv+mijZ0T6iStVaLYn8VOllYkM66
zyBG9lmqpi28CbXqe4BwaYFSXNwLQiqlUSFrd4f5C6t7gjJL6CeuJNpQ72GI
knK93jBXOgR8d7Zkypa9e8yHw0XSWgyTJAk0bcogNFvaHopv3CqlPctD7w3x
6L+ykSBEyw9dPcF2ZjK3a+g5jJ5BdbiXKJ5NnCDlsA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Ihnmvu0/XkyBbXf8ebz82LJgFdAmfhMn/b5XAiLtFIwxd1nm7rb4hF6ZMWoF
P3V4zAWo9/N2pdXpFVtVIEfkpgY1ye+u0LFZOUc9S31sLjiqXnb4QZMBCjv/
8MOTSw+pfsj2kCkPGmlvWOnsBKoF2AfKCOP5QujKlHKr5HR8RTY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
oRMM4q4YyfYiMOuXpQzZakAUOVZxjV3Dqt2GdWD/edajKLbLDnx8jSIsE1yJ
eqdabrzTYCK50Hm429Iatl64u7Cp/yO5lXfgD765LYkIfjUHQU66si/FBmcp
pXb2N20GNlzaEGbz/6lsiPbTJKEuD9sumaqlpgexGM92TKJufPl+BGNt46Fc
yZ5YPz/Qvn8S3FItWZO8QmLvurpQVe0Vz2HjRrhtVymccj4poeYJutzxJFVI
47GKluZc5dmlSRFKSTX+WahXFz3U8EXcihPqsrDItDihVlT1v8MaBIz4E3nC
PBTnaw1bydpBI7lhAXXYIyFdmcSpkflopkocsIzNF/TJQkMfD9l6q+MDs14h
acBQMPi+Yjm76d9s+d2AFeyTBMYzzrs3fw5TW7hwyDOLJQFX4kin3gStHAR1
fMLeH1arNgAzQ/45GGzBREFXsAW5c0tRV1Nrb/+PPmeXte6w76l83ILTVqGS
YPe3Q/SCPQ8O/QlJKIiNTQWD84PjWpdB


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
gGe22WMXASkDvftaC/XS9SsIR5Wnrpf9GXQZ0XLkurmKUbCQh1Yv8sY1UG8o
wc4rYRn9V3HB/isIVZU+J0rGKvH6X5sLJaL1QNniPaBY3wy5YAQoSAU7f3um
torFT2gl2DwiRq13XgNGijwWikAj3WuXGUAqJre+IVscBn6IFI0=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
bmxPtUI4ZDpM0Sv8ONtOmeTBsy2WnbbprspYOFu5R1XMcgtZa9jh4b0Pketu
5KJkMxKzAqQLuY9A5j4da3uJ0xOqHB3AhRqDERWnjNm+raAwCbyVW3mkjraM
7XByonlVhHut79C8qY15laGx/YcBbxTfQV2IUZ+vxv3g6VC33b8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6224)
`pragma protect data_block
LtLARYDSoKBFdc8Bj4NRXTVNzKY8BeD2QY3rZfJUQEauu3P2F1fN7rv7wzOv
he5CDOvk6WnQU5OKXbVYU/N8WiNILFX329lj8nPPTwu/qrCs3PBgMCLczljg
DnuDrepiU3HYiJkhFrODZPCoui+c38HS1Vg6W6urqJUkMINbdLCjqG4UlM9V
5ioH/M0+rV6AJYTCNRqI6h7lEkxdjXR6hg8pPru8gqr/kVbzd/LvhwO7hrsl
spO5XujcdP4SocR1OKhZco8JefMSPIi0aDARcC/qO7+RQwazFoiUx2zhCtut
3LsGg+2adBlVVv5khP1Tw+Twb1EAGZKI3WVcFTsKj19HoIE54ikoblWpC62A
1Pj7R3FNJ/6AJdklYm/FCH1SvnT3b3gjBa2JOGHRgvNbZsFupblaEHTA5P8u
Psv40qyE/SoXuX9V6aXHvNeG0HYvGKITehDSypEaiN6Q1h7HU7gLE837qaJU
u4HoDnmtrQfDEieNdicDf9bIud6A0davh+kTgxNtLrr41dPNhFJN0gP9Nkt/
8ecvqbrOeqcC/K+Qn/zMmTCQ4PI26Qr3XwxHiSEGuYTt2iWChf6Jg49dxXBs
DWJ5Uo5vox4iKvN3PnNS+maSWmPdXOWwBjlScB2M63KVSfF2fvFWNCjTB5yA
Mw78YcW/TGv//tr2GdkXVNia3sicS9gBQI3eRc+JL+GYqRl5XbydNniOwVsl
Qb0pr0eIq3HG+XKVZSWJn42iglY7CrkwW9qJhfsr36n2VmKGBoOVZmXAzk+t
vA+7pSt0Hf5Lrmg01IlV2zDSEHU71G/dYGv0yVBmB5hsMxDznveynJdZpXPZ
Xn0jBBgP4I/dkEK+1SDNxLWQQ0UBH4NGTyo13gDwxXkBfFGM5n/BcQDgt91F
UW0Xeof0pXhThLlHGTPfUhRCkK6kYaAx+AcmUGgD+oFhfw0Uo5uZO1jK5fIK
YZblbj6VKlwh8lTraNVx0edHs9U8xKofcnKzxLNjI4/CC6i5MWw+ApYF3tuh
lKvgP+r6Q9W8aF58KXuWkYm6CX3Oj7abxLQnDNJgV9xEUxxHx85JmlTu0Qif
t10eipRYPSzDhJv4rDVuILRWKJIKbfYcYs6eDvxNKf/g7Rrivnv/CPYxaDYn
5TH9kERZBDFUoeOIQ+O93rwQkgUjJUM6HHtWWzESZYnkDKUNwTgmmMxbsndj
sjDri/OGRr5GHyu2ysnIt9va8mzdBl0bnPruVTWOF3PuoAcYi0Z4FL3lvMPA
5jkHP/+iili3N56R/5jt1W3rdvdFlWLiGNis6FafgOLrkNcteKxAAYpA2j/6
X/Xhgn1tIk0wXhJXUV7YKrqbtE8pX2Mj24LV2na4lhdMbx9CPvD5fL6swpE0
FraSp6QBW46AA4rgUHCGkWSjAmI+CPEDVktpCOeBZcsWUKlGSWDY8QT8wf2a
JZhb9me6AteYdkBo2w8mAiYJs2yLXLGUShY9OlLH+bTsgAoiPxk8sjmoQTmW
aZiN0MdBEZp9QIipTT19GV7Du9/KP39ab4KFHhaA1/Xc/hKUDHTWoYG/96cJ
ys79pEHQR7gFbAuIj0xECQwaxnw1E67G+ITlVWs+R6xllv0KCn7mF4ggiGa5
XFXmx2bWdz9ZOIi32ImjxImwzzCbbKH3acBGFf4Z/QLuB+snLdDZX4eyQnL2
767WP4VxNSkSLndTr2gwynwBUpciYQ2bNjDkIRCndnm1WOK3fR+ZR2tzkuo7
neX30+q5i7hUVPfsV8YS6i3Lg7o59lXc4+TywVPd22wjRisPdn8JgGsESgdn
YMNbnaFLAwwP5HwS07vLkkHRXUeL81hQTksU7MMr1Hdnvx67z/AwyIxxzWnU
lX1efVd70zyOyRSZYsumeBwDwxJM2wfzu0HQrzOGPKnz23Z2hM0eG83P7Wfp
eohJ59MTxggweWwdraiKEmwy4VceDXnHFPFDsowC8fyPzpv62tvuLyKhCgev
P/MNW7yBvoCsP6EU4r1uv0zzydgG7YCdEMnNMjYeSviCJYdf8ccAbL+5KRGe
v/qS6q9u5a8hhojwKat9AJuSqHSjvz1CK2XGf3byl0Br/T4odjVplbRUb9wY
YPRXv/1Km8rMEye3SDimOpwr5iqTdPvr3HwFGKL9L0Ka3gHdwlL34Bm6zm0v
3LwR3wpRHjWAfQeHr/RklNg3Tl94Jr6qd5AvyYMFvSTM6wqkGdvXeAlfoqYQ
h+ci9Ug+szdiG1xuOgzjTT1h9DDUV095zJ3KN/x4lDutU3xsiqxeYon3VzSw
D0AG6fOEGYAiGRGUpS2xaqcv8NaliMlNimhRClqc01QbLpzqGhyyxDq435mu
tx1YZFwxVRuIcTpNKdxQxMbu2bpzOmTqj2jTHu09qI/wUPl9LpFiFxl+/no/
N7mJM0t15Oi2fe6laj5Ih7P5STVicutnZeiqwgfk8KnPajtBlcya8i31drxY
Y8Eg0oQ/4mpYnC1lRouy5ChEjzGPAZN/34QT8yx2PBHaL8L2Usv5TM2ytcF7
zCynO1DYIZc1pwQDyZrdqyfwP/bL/ic01QKSL0Nbg1z7zM7dUVbQtlNgI+Rx
jS/lur+uT/REMiBK5SoVEVFDckvrXHc/LwzU3Kv8FrsukVmPAq0P+XMKVmE6
d4xE0v96r1p5waJy3MSYaYC8qFl4JSNZDBwdD9RwOGI9Mv+gev/xsDPhhZNo
q0prG2b++c+tW1SEQDkOh9lMtQoZa9/4Wx78d9U1ndxLZyxpwsMqq9QsWDpE
M0tLhhLcxnPZH7tbC1jOLI++FIasPzXMpXV3g1de46lVnaEv61FQSaa0iwpv
zqHaAKJ9Xs4NFWUzIQeVoL9eKrOD5/3yN6JG1hWfRxVE7R4xlYEzrkl0Rg9j
wSfq13rYUmQiYkGYOPgV/Xj3z8LrhV2H5pAsGl7eqX36ZsFzlfkrdxNdS+X+
9GjcIY5RaPPiNF8TOlEr0OxqOp9QVEpsFwJwHNXY2mPR7KMZ4xvSi8iZaC/d
dCUAPTi9T/eX1EN6ZMCtrMCXpnj7WJK3wonHItWkJmQ0F6WquddCwJgRmLVR
3jRRiaRK3hR6QGLVL894wusp8Y9s4zziDYy8l6mMt4gz2Fv8mYO6sStPWy4b
FOeL2ZvjkuvIuRbCeYn1twfeH7xRLrGjdcjCFcniT5/n+tROF8aA9qx+HWGS
zUQWnfuLcp3x16CiWtvOCzmqMGeb/BP6Kg/pmpynImEw7KTXibjqe5i2iTkG
6con7COiKbTyZhMwfhl7gtFwk/8T/0i+pJeRwzgZUDb9GecXtovMcLNWkjyY
PUjsDQHSYcm2nXcnGEBE0TestFlKAUWBT8V66+6nXfTALYMcthq2VZfSNHr8
kOHM1hDrrrkWae/KvoMN+OU6tlB3Zkj7oeUbgaUaxUBNcc5aH080HVwiYjFt
Q7NCbjYHUmOjLGi5HMEh086xXX5grg3IZ3vPVnSZSv7PbGkx0Voxu7OGuvI2
E8O+IAmrzvYLu8Z9N3SzGXhFeokd2SYjiHJGX1X2iHniN2JpG8sAJGhuU9l1
q2k9e4qLj+sxY4D8FE6lCmw+1KlTEkwTNrhzcMu7Kx8IMiaiOmFlVYclsKi1
vF9a89DGwJz6lrDv9WqukyaSQryIhEtqzDjWHbYXbpmei4wdaVlVXR21Br5U
3fRjND9gcU/jo0+6aocJcTvUfwCh6A6ZHQ1iBvU8xdjFYCotuGT2xWV4Nfq3
O+UGm9NPcf6vfQjOfovUk5LVdWVkz9VM0DacR79HuK7WoyaZeLwovyLbIund
sILEvSmRj4Ms/MxYr0Wc2cYAGIrPJqSDlJu6dE+eT2qLNv6wQxY4BwH0acHZ
2fTtbqIcwex1OsN/tyczIfEheSqUR0E5xYmnAbHS6PgZi2JT6usgxUw7B3bs
C4VINBhZaVlxOPWd7zDDtWvB+9LMzLMBvsJ2TmjI7mJk/nCB+wbXm5wZMYoJ
KWzRrymgDRdNIp2g7ITsud/kKht8y1K/2dihZwxTcRl/FLjlGM70zrMeT2T/
PlALUZigiyfpsmuVMHk2rSvbsy+9rpJ01ReapjqZbcHGGyaVUpj9BhFyFTOx
OaSynoeXq9t+znXhSz2XMISsl8dSoeM7ma0NSskFXn0DCd6wEFxSg4ubQrMK
NhCiK/XGV0MgFR32vMl2bmjhkV/BPp9D1muL3cUQDGcDx0WHWf1HA/Vd2svX
t3iQ//HMUu9DDNzi0kKvsnXazNaLDptkdb5cqDfl1UlUc6kmDLerk6oMjdrG
AJppNFyhzz6C7L7w0uJBkx+JWnK9OhmxXyFPaWUqOwvl/8prN5DriMfv7nSS
FgK4HfL+r/Cy5W9MdjyXMpC6vCewLssCbSWy2YgmzjLj7RAzlt66JChLFWDq
uk9jQHyO2hrEOrFee44hhYGROJdwR7TnLXJGZoZ2stNoMX2sxUaLx7xalZ5I
34ESorWGMcdCw9u40w4LWCjBLONNUP8Gbk+l0qKpMAJ47jAuOJ9i3NQa519B
D+tFeRfWteFxYezJsVML6myDsYg6XWqQ6aSVn5xnATvtjZDDNXQp1YqoqxUe
TvQ2g6n3PbXC5n0II5vklqNDjcQFekn0KvcUe4GeSVP4H9akcKbMmO2zvDcr
Nr+HFeW8ooqNDjmTvYmH+XfGY5A5VUlr8Wcaiv2ahxNeR8Ixj8EME+mAGeO+
0HqE1qLowK+cniU7dHvZYNlKwqyvr53kTpUehWpCqsPpLc2pRIWsRmi09XvI
9+Fhx9W18j7wR6ahdqsAp9AhpYkpN9t/XwBVMqjdx2vXkIm6asXjKLboJVEK
jeI40EUmtEcj36B4LrH7ZR8Bq7k4F76K2d0CBaEYauJMUA3VlEWbW0QwdE6z
L3M79WqHa/OHJ/laJfhgLqvw6K/DFwxbxpn7qYeFk3xix+QMLzKUGbxGyNKl
9OJrD56GnDTiE95bAoWuvMoUUzXUbSPZu6okp5OZQHzFolKXHAMOfN2oeLzm
GMR4qWkFZrjtuMWw/DJnuz+ulLKt/zbu9eyZbhQHam/vKFkcicK89O9VhtTH
zr18pE++Q4Ioiz1JMkyJ53+PyQCrdss0AUZj7H8zH6cO7ygUY40EP2aNijRd
WUPCY4btUtctC/J/AO31dJAdsbbLkV9fLEWKyB7H2q7lOnQzpoiyklPGeWmq
K10UXuek1+wlY0pQVSFJz4ZEWtTY25yM+++lzNFQEuUpZCk7YCZdJIaUkJ0r
zjy2qzO4YS9lrnrw/LwAMD0Rdute9ORsylQ9Ki5g5MnBETHrNctW9SH4Y3v5
nsPpjkfbMMkScDMM5INtnwzTXlFjGYjT46NZ5DFQ6n44BDks62YX8diU3mJo
pTTgyru29XUF2vjNc0aSIbgQn7qxZdXc9kZhgSrRS/CZb7UyQyMYvivsM47U
5sq2VW1dKxK8APY3XIyd2f+/TDj0Uo3NpW4SA/BpfNkTV6DpXhKM1s5q9tC1
ghsxgXcAJbx0FzWBGMH8XGHgzVL5+1co6NRSH/a3+4A+jde8slGBLq9Z0W4z
JGPKLnOdVm2GYcrDJXdx2QqrQKgxmthBTiwixk0C6UbdDhB3FwKH7X7a7cst
nVvsKx9I0ktOZPSga0m0n6qRElddt+HWbG4Nmw3cxXfBiZl8hFtmcFJ1PC+L
W1p8DZz4Gwv8c4pxFqV7nHJWsA62r2JpR9zsLgUcpTUmwLeqripLrBY0DjR4
z90rxkKyjEjfxao2LcP3I0jOEl9Th6CouGybkBw7krNVWLKCWXhB9MjGUjpY
mAeglC2KaIOXEj+IsW5ks/8MY6VH7GTaRsK9ODWv6klauD/O/M8b4q+D2NWU
PJ5IlvwwlKaXylbV2TvDAaEn1kwSeus891u9MhYLuHZ2ST/DyVHv9pG90B7G
0tSL3VM8IiUyFWNauW2bS7zpwURMVspX7MLeoJIKxregwCKfH+SibRO9CTiW
GpxTir1lLoAnuXkxNSvEWyXsSLsCRvge6Ll/hABJr9firee8cfk5kXWZ64ra
a6Wm4si/zziDRfKQScNTxxdUlQ8s6CNhPAY5iIRqrGcgovFMmvpex6DUEDn3
RkhJmncur/IGLyRXH3YAP8XH2uhv/mZzkMxW6AcwoH0+JJhgDUTXtrX/S9fK
7JIyxr6p/eg0n2AigQ3DMwu/gy0HqoEadvAAJ6pLc6bVSJS709z85+LxoSK5
Ns5969t59Hvp6XenUi7MFLcQulBTJ145TVAfxobpzT0P6WXrMqPXb8xwVTUl
QfJhKciZsl6sw2kx9QR8/+6IR230aiBfoS57FHeTnkJXwXUlQnKV0wBQpoZL
xxWDxX1R/xfQL/D/wgI3DOasdaEU0OB+9iSWNVu3qEpr/Kaw50bO0v2KPjgL
zzF1AsT6BlKFiOkiMzEqK8hHFJNgC3w0sLV3DcQqL4JHDsqy0sWxvlJUoD62
P/TOYv1sqWWmDHfgwyQV7hFTZpUCkD0mv6kjmbMZP+M7Au5UdGGdtqu7RAC7
ElUsXcwHMoPh36z3nW0N6UBoPmaIFmXWcHQPOME6q7ITyq5c+emflz/GBnJz
qWwfvX0RjtGafInn+EaYM6Eu1HvSMKpTQ5wGgp/Q2KVf9XkUdBHmb9B+S/h5
/FnmvsWDS72UTjzThpnZ7MkbyFfaS9PdMGPGFcrbo9OkmXrgtGH8k/EwkOOv
MasEST+HGK0MzMnq2vyMqOsQZhev/ITHk+cuqVI2Odc63DSI3qcg0IKqX5Oz
0vOcR4B3LUHdzkUvX+X8RGhtNCoTbFLPqql1x9kBggE1jMjfqlObQMrtmFsx
kyIHCJB7kRXPBSFY0fENHxl5/7NM2WlOk+DOHDQRIxkV3cXAcmUjyBOFnjud
QpA0/mrbo98gTqPOVgQJHOJ09wVltL+DvsWQ0cwT9rKrI4Met1uRlHGWSyB7
Ujp4S/lBvLFZ2vK8gsaOyl7j1weO9BvTNZTPIb2crx9rfpxC36XHwIrYB41d
KePK8wrSbk5hr0kR9CmexH6UmRGsoWNO+Xw/m2LFu804xchISQfO/MJk52Hi
lATTw55vMvcJtkqwVl7Yzkqm6S1vxeCedsbW+B5MPNzB50HjmIx7y3Ohsd7+
nJenTru43DUMDvF1LxvrwwyyV++SJ/Y4zy1cEK1uxeApwoSM3oJ534IYzA0l
P6K3gzTWUSbCgtng4eUqyh6Dz6/nUbHa++dlzEv17qUaKS1KpmAbm1X0g2TS
XgEw+g7M3kTdJzH69bSnQtB5yXyn+FLEmYgYNBVRK5R6A6R1wwJ2sdp79V+X
SQdXxcKn6edHUDaG0grki/p+pEsqy+PqXVwQ2Gs3msIEY0FQIeYNsGYR+XH5
WK0ILaZzHJFROmne+hABtsnHCPbFOKRA9PkicaKjvXtH4FCF2LRODQmwbB0n
VgAYLzEOPjc3Y/VHvsp4dqYFHfQ2N4EPq+gW5/Lj5ExFxWuTKfMgJvGjvPGy
KOsMEqke+Rxh2QYPVbA6bWOVE4pTwhl1zoNDp5k3Wo4geI0DB0qbfUkxpAnb
BT9DmQp+Uz6J5W27pojbcITFBvuGEkL3PZvlVp9QUrjKCt3LpxpAlqDtDqmQ
zgfmGnFde1BQR88fwnrcircKZKmc2vlit0dVMOQ7jWws0UH/bqSUDwqob+3W
rfh+7byOiAxfYhOJLRh41ArdD7FKwkqNmWfyf2XEaaCMCl5ai8vJdFnbfcbd
7eqXUULqRLMI8lcnV59AbN/NSMvZa3EDryzIIJxyGb+ln9CnBk7+AOlDGGfY
81mD9fxHuDjOrGczgVloMUCkrLuxAfYQJJaDaKRCNPwSlpjWf0M5+bBFqJVG
XFkkGPWHgKkMxKw3xzWgeo/bOs96FUgfF9fKcKvsfDHNyhX8qJ27Y0Nu/vDQ
UqUcquyXV7y4etVVFhHgNFf4DQ1K66baJxkjnR0sGyYyfqJyd6/AUWnFVn1e
WvexZFC5f8de3IFRrFW1DlrD/aSXb3KM0+KmAfIcqzmFmKogl7jM/ncFqEg+
jaSO+lPKBWfvIbbITJBsT5BZ60kYGmNIhCyn/ZWirNQfLLnLMzIUcY48gCEL
E5XhMEBUoIYNvN2Qrb0uyJo7lNGAxypD6sVpMqiCNdTgUDzb6rjRGcwX/HQw
4JPYEt9m5bfkQVWH+IOo5j22piUOKAFQsTI697FFCi+JcVS87CxQwnDG5MuA
fe4khssJCGNQjc0Ln8KW7RmHIIYEGt+b64CGIlQeecZt4l2+7DunUcDNZtIK
g1d4VO29iHV2UWhHh27dL+UTOnAi8zWcYXaChr85ym/ZLRudk7lmuH0X3zSp
5+JmU1LLURo67Mzquq4=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfSFuqG6aRUGyhWNDtlHJdON5toktsrjyikIizlPrCpHSO176vO7qCyh+WTzq9mLB3kIrmjO0oXFbTUu7lQVbCABMGfAWrH+S9/4vIQ4pCHf0Oqoqu/83fBMsU7wXFaWVR7EOIli+/wnG5uHtYhP40Nut8snCr9pYACscwvhete0YgEhgNUynwkQusAtXqsua4l7UF2i237Yz2DrwgGuGZ1E5QrFZmjQBYhJ4sa+l7xRD3bKKH/w5z6h0ZlY2rsC7YUqGx0I1hsw8VPV7zkipjZX3Dx73KnH5npO4UPcpwfnw6xzX8P4TxkE5giM8DCJUAMYbMnHf1fsjK14oiGvSmZpsu7VqttVvzzfFBVBm6iHJ0bmBx+wHSv6B+HHS4ij4N3QQi0wRm8++/MnThvhh8mZz4k5XqCLj9PiWEo9zIuLL5M6UrE7wdrl9rhvEJLMVC4YdMZYDwA6BszpwEKEVsWwGdFQ/olxovEU07PKj7eFGEqC1vsT5jZDQcXMQCc7iBcZxhrWE65MUbY9V/Y0U2mr4b8xhpNWQllUyPIviP22xhHXs647zm6H/FsdXt6F/l0/dw+Sggfm0/Qlnv6TzCeDNSffLD/q1O6+2nTSO1F6IGL8A/CECZdKnDgvejDqUQncQA59hkWNVy32VkMTFwPjvnmQsnJ+XbswpEryCSZGuNne6ZBQUL0h+Qw4nIeHobxKm0SHP/x5jl78pEOf7mueshCAQEMA8pMdaVXjjvf5nekDBtUjj8SMaxDnRE7Q1jRhcebRAZFvj8qTqfljpN0M"
`endif