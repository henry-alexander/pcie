// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
O10CBU5v6A8XLetyDYTlnXKauV7f2qFmJlPEf9YE9UFcr+wm+z09GN+qht1e
NtpOwDkF+6Z+ZxMGk2Yv6KNA9jYCxDNKoNGSkqj1Q8BwXNn4TVrmlODlL/Nj
e5w5Q3qEoZRp1epnDGQ+2v3afaRJ2Ve+exTp+/biVbV1JTnRwDHQeWa8owhb
igFmHD1jOA1xHniKYe/RpVM4khD2JOwj3+5p8GHZTSvjNEGIbiewqWrxVKy9
f3tz3HDVN9tsK1vzZj55FE3rrejdPsU6K5/AlWIA0WfF4RJ0y9tycGTjrhUU
buCBSOc53yf/JYc1l8oLBI9ziYx7nj+LiKLpzJWfRA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fjecauUAvAns/NaNfCOcv9cTNB7eYY2ViF6IM9Lh9Kc+jucod/+v5CsKYUvP
ZCKAUQIQI2H5CfimIhpkghznxnMDnsrJKZR7DaEKs0EM5d/w4tU9LaOSnbw5
mCOHD9su1mU/9ISmAFuBxzC7KaowFhYYrzcCGw4tKrjYkq7e+iVujelpm2+b
Lkl7/cGRpYeqO4I45NwZlEt2VpeDwfVzG4JRGSCFfDla1rKrBPTB/NzXuz++
SWZ1QfusSQw75yRMXRFNna2uUD2mlm1RxGSZiFnHfvBAOiVK3ymC8Dzijf7N
q5XaWSyvzX6IMEheCr2Y6eOv5nMVQ1DM619/OzZbLg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cglbib2eXP8aL9LIJLdjIKcbH/8AbzZhPhq9YrmViwvfN9QqPEeWetJBrxRU
LBfPYEMEGmAUeNXLS2sMbmt2+g0oViL0U6dERWYQdWaCpXpsFdjwzusp/jRq
j8luKZ4+3tnbb8ynkzgXqj5QRuY08kyAkhu66XRHfY+VSIe66C6FYOSxtTAW
4DHxwiRsEafEUx+6ekZZOTzCXxUcQMyAvZuHz5iH4t0/M3THmBZEyOTKhD9c
3KyQf4YLPRuzqbW55ritbUVqP34BwN3ETiVIXRYVYmFtfolNsFHHbc6FMm+m
/RBik/iA+UznCqpQhtxRkJ/uiEsFL39t0vZy7vPcVA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
exIXpqIK3OVH96b/K6fIZMSC3SWbbvPQz9CXhC4jt9hPY4Dc977k2svsETzu
dUoC7fsUdAWRK5EnNMzcRZGfgLePs0RQxhwBOsJmTYoNlaj/d2CmdHz1x0n7
PrOxXk2LyGKL0Z3+z1eY1LWTOflBX96R4s9Ncd2821HMdMsyqjk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
eWOdTwsi/rbpgJkL4eR3ZZdOSpQ0hc9nS+H7WfKM6G2A9TxBpazveUTP+bEd
RtszNKrRdO+3Ybw7R7bHJgbcjHFdkDn99vADoJf1S5KV9w22RlVo2eKHZhyV
ghihIlo4+2Bp7Ys53W8HQqSztpe4cBEbIyYwcRrF3tov9usk6A7kcGnYpPxj
z1Bi5QAP7Pc7SaDbeerOgfqv+9q1KZGB7Hk7GWI+egWRnfgMvPGbzkW2iGyd
USJO0gXduHkUasRsMbn/2fEu1XQZNrj1upG227rVUzeQ7vz4iNQiI/coVpfL
cgZbohUF62zRUgIYRaUXJYY9HYYrtEX37M0tsQXb/I5I0WTo8wyOmVsii2k1
jtAarALL/N67XA3jtk6wJr5I55hYSWjex1cK/gJPhMWGBZz2aNFSgGtn4NsH
02i92YsdNkRVQmHC7h5Ic9Ga0JvAalV+YliChVF6ErN4Km9d8IkWOKDaTeCQ
xbSwY2NjV/j9qG9f4Qiex14wJT2zPhXk


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
VGmSlYNDWnkGMEkdCRlXNZPICIaCSdYLXFtJaOz0HaU17YCARCVJdFYpxUgw
4HImeT4siSDL/49Ripu5aZ7qcrFEpSElhewd1VgE/R3M/uZWjpPJsiQpY3kD
YKvjXWT7CJj0zTzV6mpxTRcoWizG0uSfUEkXdi2xzWsb07yMBr8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Bli8brbaBgLtXzxuHuKbUUgYcSY0jFxiYSp6Orf3vdRpl6u+N2CyEllv+UM3
ANRLoPy72LanuSwaGomaLchwTysisFaCCyiiN1XXHKEErpI+EG1a9B2MdSHy
xar/kb/5OVPgoGX/+Hg1BoJcKE1W4AiJR1SAgEqk4+YVGpI+MCc=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2160)
`pragma protect data_block
lt/Pqnz0rdD+LWY34kXaKldHPeBa5XomCVRb//ZRHcVeccAMLx/IBmahTmGG
zbH9PUrMU832DA7GcS1+J2YDkaXpkRehM9ugtGtD/VNicFsnoa6iiwM7ubfJ
7AGoXWICyeJ3QiZKGd37d9Esjzt5oon3TRuNy91pBjE2gsSBmWp0mn5uEPoP
WTe/aC9nYs2CYZeTQ2jVgvCeNpBRtuh3EqIsvYjzZakDptYCg2jrQU2/bALK
+xQTcOfq8CSVnOPHKkVlx9ReVuCMlN+qJdm+NN+OrsOZ0ecNkErcdGOD3K69
uH0f/BYqpuIzxuQpDLqBfTDC+93muyB7gE8kUwWw747kQNVg9ypETeTBQ7Pz
iXS28yPw74kT+BfM84382iU6bA2FzF+rCxCyzBegZNNIW5zyZyKQgQ67qeHV
T7SU1WvjPeF3a6d3Q5eyCL6K2shQD+DIZcDxRrz1AdpWPdWS5Ou9a0asCUa0
lDww0mqF6qzFYl8BQnjCEzqAkz44ny9NM51qXxiBzYP3h7bDnF36IArb1gvt
gZ1gpA0ex2l5YLL0gkmCzQOmpzbHyKXeLM8tWTeQyXYGhy0qr06KiM98rXh0
XpObqlbwOPMrfQWGM434pjZj1ISEcn86wm6hWogljYkYyp6s4nplFJM84utt
IsM+0MUgxEjgjN/GuKL2h3CS6JkSoOYJF+Ls0EvLC0I+eJ2pJ/G4Skfl+oqZ
8ii8OlfUZO36eBWCfXsS2qjLuw9odkTeldWSZXlXqwxEtuL2ypjqz+k8ONWw
tuL5ZpjDSwZ7tfB6xLA+qJvidLMQ4ximSi+iJTi1/v7P3msLiC/9eqTxuwha
CWjYxnhyYwJNLkgOE4yKH9eh0HQPjqgPGBTe2VQdCT10rnDe3zt2WopNCvLR
FqeWHZ8n3RFOkBXisBhPkA6W7xAM0NIuJqS/arthe7HZ+bAvgWeRaPP19/8O
4tXX3Ek2WwNqz2wD4H7nZOg1L8uU47INjl1hOB64+YG7X+8VkyfWBtiCuG9c
gbgbdRyUx9VNNKDuFA9iv7BGpJ1dJopW+OZPbFxkL8mRlY28SEhIWYZG7JCu
MUFVMoNWs7mDAhGDMXqhdFiDHlKgj4htXKPC3kO5ivKAzk2jvTb/iW8lztV9
7uzUwcX2pqprYXux7/zmZNKygwWHo4J1F5sp56Awa7X7FWatt3oDcrcCqgk9
bX05rOVRZ53m/bhbM45EcfCfwdIlKjVAx40Wo04acCYvTTToAvF7rpZhDPLl
5tnG5co97zcqKn/3W5AL5zPR/uk+qPwy5jk/cDY6+DsP5MfXFiORxQ3RILyA
YucBpjXIKkx1LnblLKgG+67x3l1uWMZsnB/7MnSun38UZTw9RKKccoYbTN8Q
Fw0J2KeBAp3F3pCpffmhUYt+0klJFqNxVL0t/4BhSzKJ5datQX8edbCXh7um
ky1AHsIz6KOrXz4lrDBwD0vmRgW3zi1dVIpc/fmIv6stv4TMtd6OeYAOOXz9
54RWieXFPSnCVaBDKuW4R/YvbBgi5/pbG26K+5Ms9xrb7HP/tNK+B7Ljg7/T
qK7xQrgBiXG3zrTkCFcpaMVCehmlVcSamFJDLJRo8W5sh0pefWJ0eSvzlmYU
GhKTURPH5CbmqElZImhx0WJvbJudWNX+S2GmDI2eUM2mCtmaadZYyhxubODT
9ECydUSTFK5PBoHCowsYVUeE9PP1tHyBj1iJstV4FD97Rtxl5onACra2lA4s
KsX9USYKQQzTTjQrT6Q18InlD7W6j9ERQB8MePNyBiyN6Kjn2YUWuR4HA1SF
yCysal9efO533wspUTHqz9f6IxiI+iGjFdqwbfDlJwEawWDvwCkWFFH4JZWC
1CbSJFlGkNuRZDWQMHzKPGBM0V/hkGSd7oR6/ub6T7MEf2xV++J7VKmY9muT
iTUgbAH4iBEREKGzpJk2s2iZn4ubr/gir9dn0oMligIy2hgFrhV46vRsTtjr
RoWPPuAZwSZeiPTLyDUWBljtrs8RA+3i+NX0AuzKOaf39jc0BmmwYr3JOBZL
S/HQ9IkWtyKzcZC32t3ze2RDtClUIvK6JdmgBBMqsDe/4uBMmBq/IQ6X+zT/
Km/jFu0sPoCo8l0L4EcDoMCMKB2a+CLtK6XhVjeIo/k8Tdofn3kdE35yv9HC
oNNmTCjmDJYEHQhy+X8Mq1SIQN5rQ8YCW/BODqZkDrK47P3694X+0Hh297et
v0xKFYE98WHRPHjpjLyVSoH/j7fgwUMC6eRakO9VyiITgWswiUT10S5aj5yU
D8wz6vlBbsN9PoDBR+7mnQcMRjTgQEOef4r6hslo5l36BsrMZwW/9vrL7GYa
hzI9Wq24f4oKQ2EjXw8wIHaKPq2wYodYcXmN3oHnMaZ259hX50QDUke0wLcy
LS0ak8zQAMF7IMqxPahTODaxo05D48lOUKhsk6aWrjwLjuMzgTZRirMPo34n
VSHTyRGEIOZlsV3/+IST1twENLr0UygWtRutCNLNyJawuVRVq2k2BQZET5SE
bIx/IwwyS8hL4P09to7H7dkK/QMgSq0Ic0WE5mZ+ZouA8NNqCmivK5EAavZH
NHip3a8aqsesKiHP40Og6DnogRKMWeXaoz1t7HuarLoZhHAIM09d066WDgUT
As27hSGFWvk5LjoibV9aDqbV9tVixQrxmOfR951IjwdLYhjrZJEdEVpJZRsW
HQSoG82kLhysAICmukytAuboi+IXVx6xe+nnr49GUJTPpZtddqTzJnC+EXhb
fhQHn7RVyZAhC+QalgPWwwJcpu6a/JTN9moV4BlmAnGHIntfyuUltgPACluq
QIycS7zd2br465C+FJRxAcr1ejN1VtFE+cS8XSSm8JWUS555HhOQOSp8rCZb

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Zc9KmeYltYUgpo0RPlQ0CEPX9+29UJx8hnvszRjZLLuNk4HJ9IKtc/cmu/ueasr7j0VF4908JtI66F/kF0AYqURi+Mi5Y95qNulunHg6lziZk9GRf0HfggsFNE+GKF5YqD+LXhJ8yr7krCxjUtXchhStMOs/fO4csrZP7XioJeFYPcODXbGzq2Tg6stNQ6pMKRJmw+sV/bfJVtEFvWvB46/T3GMjfF/mgFbmQs+o0q4wQtcBfGPV4hpKiClES0KoSeEv9Yy0ye7ahEVdmmrRE9jYWwpw8ko7gxoVIFLZsWJnyYGFu2ESMmu3y22iyGn2dmHqhWPtaL7a0ljbwyU1tffO8Yf+GQ5yB5XCGz5MMaHF05mxqKpCdKbfCom1RT7jQ/hnUkfFNZt8Tjt0693j+F8riB++9Dmck0BIwetvpLsdt9vVEFyupnzDviHrA+G4Lh8LJT7fA+QIak7Z4tuj/uFyopJLs1WOH4Nes3v5xnRQEjjoXqVFOy02rBRIZ44cT9DLc70RDfcpn+eSdcfMpTb30GBB/yBUg7ao0XV/kV6EAFckkFhSRgKRu3HNOTQZNF9ff9qEiplMRNjZyqCYQ65YhCdF++TTr2l9FlhXC4EfdFjNNvRO7jl/K/aJgz9Npy4uDE4VnNtxJSjEFMtvTlJnospU3G/05wkcWnkFfu29YPurXxOqI5K0CkeS9tPjLxx0z4P145kUE0P2Hb900zBs7K0zHU/uE8ru9+4GiMle6tVhNEGURfQw+8Vmn3cnl7WVg86lmQKJbo9u7kBq5otBC5k24hOXleNDatxi5AvR1RSfuVqQZDjUPKx7PVds+vT1tVV5BXciprnRryk+isU+/QuIZWu8haHxxh4mNPMH6m65FBgy6UrfPPpbCmahvgB8huEv/jD0jdcDlJOh7e4L3wiApZVaIA//mPaaj0c+p+8oEySQA1uqyghbiCJhZwgMls1qQVwY0mKTacqGwd4BW+2kdyWT055K6A0GqsxYgKlobcwOjAN65xpiLB1G"
`endif