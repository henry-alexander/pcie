// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
D8tlcRLcAae/r9raTaUlYFg5kBMaqcNbqabUsTYeTs19sMC26rDvyrKvem+Y
wGI8V2x0wkWNG0yRBB+6DcOr6H1oFY/KHSsnJy3EdkGYIZfIQEfwdkqZytsc
itdY8iMDHQ2OXBydGYj9NtXc9pnzLTMEddkJ6BhqtSZSmIoxuUSr6rirgxez
gOhdi3sygF0vC5MNZFO7xSOs0lYaQZZM1vCfy04hRO10Kv4Bd59VpIu5eIPm
lFgFF7i49MiZY3sHfKPV7YyPcS9cckSKkSms2d19F28D0g2pVAdIgCWB/8PM
F31344dZVmqaK0H3XmLX4dDSW9OsvQqZoaPhL2GqxA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mk9NFAn7yDXmwfv0qSz2dtA8ixspOg6N5hUOXbb4rJjWIi6FcG0ZLr5MAIrv
0l8tg7Lm51SwNtrsQz6M6+Ym7aXeB+C+cgcayGOUq8MEj8jvRkOlKZovAt8I
0DWYsr5NEhIkonaxxW1wto4lotdosqTSd56IISndVgyGCV75e3enuVzzafzZ
D03BggQqzJVpkTPVDVQZoiFLxQb9/Em/lLEkf90sS5UcG+pq+T7qArwdz/Ip
Dx4S9H5XyUtDeEqodj3CisD2UGaOAHsXA/lrCzi5yolDF/LWE9Nb/K9tW8GK
eStDK2Pzam+C8R3I3QS2Winw0teoS4F2jK38CsEaBQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p42J+W8HZN07uRwdT7dMDIUW5XhgBLRAq45KYOOFmNui38vt/Ec4gPVQJvTy
y0VO9134Fgjyi6RJ9YHzKcvAb0Nhj9if+Ihi0cuIcndgyg8yYMytkYJw5vau
4+bsO3Ef/KvvoxpFh3dwKvenAfDF/DBWnUOaUEGuDUeEJycPZD0hYOISZQX4
4rV0Lc1tyIWlU5SDo8gGDU+5a3hsQn44ehTUihZbXFxuqV/LN3Ddfs7HJFgj
5quizKR85g+K/FjT88yy0uKtrRJMBE9Uvfklub8JcnXpw/mBMK1MdRSfZ003
yPoqvMyJpA3dHujij9SJHJjhEdzl9NQsPmbdVx+RWQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
K5C+oampT3AlehnDjl5DMDCgENKWVSvLr2tlkUenMvOpUzh0rYWFUMokFkaV
K7GXxYhREdrTKT6Yp1oMFm8rGmFcOTLkUzYWCHRMUKwXjWQlMD49EBNhxA7y
nUmZ638MCpRu8O9kdLPljfNrIkOifPb2qgP78K0zWG+llu0ngCc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
KzjwUzISWZ9n1h1XA0QlJI4kyXQud2U2wwszg1sui4m8T4r3eb4dPMYXh3Ty
yW45ereUwC9qsYH+0/vrpuvlwLPKSwOkbNTCS3UO9pUYAD59YEgIvNoKSIx1
ESWeSQqlOC5NzYJxX2q+OuGXCqQqvf06yxYICYMkWTnIezdcHcjFiMfXynNN
x+WRU4qUJbFavxIhKcklbYTEeTnPneVnHtfceub5S06tpXGzVg3MG/3AQK3m
aQHgOZH7JRcS91d4FT2Jtb7E8TkgZyt+gOM6/9hkAciSnuTHje7poFoTHVLV
GBARgtpN0BIsCCHfWVT6/8kNleQy6/39hmjQJpLAQCVKiXzwrFr9kxabo9hJ
p48BGqc6cqRa6Dft9pQOGSeshCkz2InRLalwrozDOL+EjR7/OsGMAEGDzC0+
5ENDcZUl263v+MvN0lSqSCSP2zh32n+ew94j1K4OW7izIAn7a2WorY36frkV
cbrFHijfHS86yhaP9t3g8EA7h6AEDAM+


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
SURwgjtMNfsVbKe5BtyOFdm62Ce5S5nQAonNdP+Y/AYqLSwxdS055jrtCFJP
8wKvAvx/YMbrQjbNGhUcorGgHlM10uE93pZwyF9aDkfFdk1ozUHYmAJ2shwA
O/oo0QI1jEhVg0jf679QKaDHqbUC1flNzZyKuyfZxwePmZj3+AQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
dQ7cKa42ZUeDOzvwzlYMut1ObWVVeT0IscJz3OLp7dn5ausHCuZSbRctPKR2
vBTjr1oEm2Veh3OkhxNefDADSAGtUn/QVNCDEerfgqoPkU3JsVaZIbJBylsD
m6Ge93y/9cL0h7gq3od1T8Q3KulihlWaj3Nle9SNSkFFQDrHdp4=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 29280)
`pragma protect data_block
bwTcWZIkAvoZRCM70/KSArv/E8N4NYfgOFM/nTYgXA7h+XgCAUdngHLbf7Tk
SKSgcQHW/iEoTSWa3MlSlrzogYyKcKpb1JtWizNPabh4sKwzFOo3jt9BaQy8
bDkvNcR/6Alfrlh7wkjqOep5F/FAAeSY4hHt9sC0a8cYch2aADsUz+da8PyK
Nlsx/qy+AuthxUIHnsqmqY3jE5Q4JUInUOqFMGvEOmbocyPqb/wYPbDKBd3u
2HvtDj6kZOjAWTX92Mc9i4+PQBK4OEqkHmwNl15qFknozbkctrWIXC7vqv7d
dX1o2UJsCby9XQ6/NHe03JzNib81as+rD/ZhbercyUTEzXIcHHfXE8lOV+Hx
K8INiAshglTS4iISCQIFTSk1Vg5ovZfvKtdqmgWZJVjT/fLgOqxUdk4SYHRQ
ONCr9YRx+OeyWflLQI4f6gdAkRTrW5t+XfF27+1v7r4KglO/eQjcvuNNvVDq
fDZ4fOVOeL4r/IEcjJA8tlQrDG2G2ZTHyXf4HJ9Uxg2aWVEdvf2cS3a7dvtZ
oxGB1+/YtIjIO3XpDLxa1DUVdSNSx2r9TSTST7btZ2yf/4qEgR1SQnKJ+ZBp
1C4GpH+b9oNBjI3v5pZWXsFQDfDC7t9Mwg4kWuODz+dg3gDDXuVsUSDhdUYG
ya0ccMDuLaY4AwDU25c1AMhaFARUZLE8gdhoumpt4+gGtJMUWIFjSfShwbwL
HWX4SaDaPKbE5jAIYAakUNZh8UZJC2EiNfzcNYtrUo2bZRkC2jyR9xsRRVlP
cDtYV6lFA0CjtbvB9tslUVZ+HfLte1J9NsVllzgVLMc6epn+2Kk+NoNlBAfM
JO2xil9U0Xe6JJXDLZw3pam6mKMfXb8GGafJn43Xw6gkdoMOnQQPXAYbCHbM
bq6QCHTpAqHimkQerQFkIK9ynyDL5FwxdyVv7k5bt1a9QEb8bhoR6oHNzJIf
SifGCRlCZh+EKJO0HvG7iireUaZNMz1Z5xb6FvYZvEjo8Fpfa3A1VaOU/9Fb
GdeBF50J8FNdnaOZsqVP2VLvKB5MWGDjuqF7SIDO5dBU4WYqYq+88GuJH4O/
iI45DbPM06EzQdaJbt5w8VlnFjmk/NFMSKKD+HmWlib+2DJdhTNJQGwDYRHx
12Eb+dfi1pAQJ/a0OHZZvELqk+ykw6dt9wyGFtuvOxpItwYXWkdQwtAXTfnO
vxWDSy/zWPP2erff9P977B0uwv8iev4GP3Pas7lCVUp/FItH2XIHqq+SnAmz
WrRbhLhkRGyZQp4iAXst8W9S+GkXU1xNXPxuC6UDKTyKUlCxbkozQsiZeZMS
2YZBzzvkmMyJRIxm1Nj/2epQiRIvYPGkHbASet4F5WjO6tLnMMwd+lhRmfM4
K89Xq2R0gI9mpyCkhnYO6tIaj7d327DG5Cquux2/4gO1uqUWek4tXcDejQQD
tTmEC6YJsUHPgBezy5CCZsNn+rH0ATve9wlb0+37kuTh7qmTe5JcsmHIQ/6M
QBP/DmCW/BuvcGuB0jY8S2clUXwn+D7dhWAiyvSq98f3jBZ7rTHk4obOIjOY
MT+9or199Std/kLHLlSVzw3mHSPhW4xvpyHpSj4fncFWpv7sHy5SYUg1nwmf
Icw2DadXZlHpGvJ/iTN/Phpr4xsuNHkmjcz2qCKTh9+9lJlt6i9sEp5JS04L
wJCjzCgRLTatseiP+k99UJIzhz7jwCD71hMbHHdRqe70yISNgOVFgHymPTTv
yAoeJqSY+bLctsDJDJPKcGOMvEWybZp7BPb+nrzXhpHuJsKfeZ/3RVwRARpg
y1xvsgtPePNFvF+Rze+oVUVztAtd2C7Qh88MlZ3hmsfGZM1mSbI5ogBSX7Yh
yf8vK+gIy6IjjZc5hI6v8Uc5RsBxcWnLwXGOaiNbeSI2pUzvr6lVN9FEDSQz
ydfRmXnuectR7ALXL9z3U+5fnzmlUINRJTNrY5SyBd7o6h2Tc5KPCxKzf1Ov
dm0+O2lb8rWHhqqTGvcZ54C+QGkMUjwKdpKxWoLLnEY9uomXNyYjTgrfKJOQ
cbdlDRSOb/nit1YJjpboXCRH0smFGOYhCr7P4F5T0JPGFGk+K05rT9Y9NSnP
grjwEHCckB5wxbo/9TDQRbITpFxyIAPagFzulJW9wfCALKocku//vSHEPxYr
r8uFnlo4DEUadU8nqcHPdW83fN4ZoPkNFBtIjLW55HK9MamhJnlsL2VXszkg
ZU8I2MS4Ox4egrBrYs8ZMF4n7svz+LwLU9GNkkTfuB+kSB1lsPMovFgxVojk
kRELt/o8keC9DQH0rned4adViSYzm3sYykWn9YGbo32P0tTpuAC3zUjyCzWp
pj1MO0dodvwwtGjB+NiEniNW1POkWXAoStubfGqdszJW5F4HhTkC1hoQ+cA5
HxGqPVLJNQBbsdreHJJTdVfJsq4g+gjWpbD6zT44VSBRMwnhoSt1fh4Yol1D
Dzd/p4M9/sj9VSvBIzC+N7q+eEGbRkfQKmhmV3836eV5DTV5xeTSXJpPeHpn
ZT00uN2nIpFKg+HcDmnjDQVM8Je0wn5fJw/0b01bDhWWlonnW+ZcYdkdAwxh
qG35FY/nUgn5v4857qGwWejIU5hJ8G1YWxJ2DZKJ5Uubd7oLU1AzLRZSJd/F
iNbMhQ6+DTWFS+CAGRhRhtA9rprbTapF8iAe/UpOLiqwemEM5bGeHuqG2xOr
MPYBr5e5jnGsOTds4PkUBQrEasL5g3li4gAUTiuXkIb4dbyPEYbBHDwtYoSx
lerN0B77Q2vkH1Ecc3IbXqspchqQ3TgZO6UXalJ+OoBeaAkZ5Pmes+LB5h0H
SEq8J2znKto+ayBpIRS+XAMxc46h5/dw5DYvHUKEKaN4kVEgCg9KGB8TPtd+
f/W0t0hoaHHCWbhQw2jnulL1isILMqFgkL5CQ2nOtXk1pMe3CA7UxKfZZOsE
IMAQ+UGzUvWLQX/mDYFufvmaNL8DT2myuEfe2MH2+//KMa8MuFFm0YuNnPeE
9sk1zTooH4uHofJye8R53fEfoW/5pwK3rte/EnLdBSFGvGxUjxjGzChU6T/b
7nzLOtucB5Xg18Bf5G1XGl1+tuVOdM2T7Ml/59TTB9F1Hm+WJt+JEvB8rCkd
j4NPDCw++vdN0WY9CLuvIru9PPbELakyxLsoS+R/dRgLY1q2I1FhK4eZFOp2
4SlQ5zi9I6F4OFl/lf67i790YTorBtgseQezbBD7DLTx+XwX3ejIW05CorJb
VR9cvpsjeVMW0M3tEmKcJ4/WKO59mj2rhiOFRRe+rQzUDWyuOgIawcD5bE+p
ljpok8FTQWtjbapoCy1r8JQITM7Y+bDzx306DjtVdH01IYIuHoX4hIE/aW1n
88nPDb4vTSQZNcrgwZB/Cqw8+mWb2CoWF3toj4SpQH3H84+uCBXiOfNPV2tC
b3qssjbrES0fEa45uzJqH1vnfikZ6fwOLhR9SyJ+aZZBPBN3GRR37209bv+H
qxsXrCZrDpWIaSCgAiw91XdvnIWwtj2OiJ9qhcQ3NejhHeoXMu83TeyjIfXb
shFLKFF1G1/C03yy/TC2ZI4OQsrdVG3eB9N4vhsDMZyJ8i8r8JGoS0M4bzTP
lBE1PBHlotz59+JOSIqk0ZJQRm/DnZxITp8+MrcbdaU6fSRMoA5SEwf6erCv
0tPv0gekno+UKzvkJ63AUi7yD7a+kXNQziH0dPZ3+j3BGQ1YFU3XjHz04AKC
RpEYb6Lg+SCkWEh7rAWSc9nI8uI5EB25HNbpmVc+Dm/QepJS3undP4ga+oVk
DoYD3TONq+DF8iJh2oH6WGka677t4ENxTPIPeK3cu0X0zrIbnjF7AEvO3/Bo
eYWDdW3MY5ysb/UnBYxEQRdgzNwkUNTShh1PbXxyb6LMkIpvvpMqADUro8kx
7kwVG5Mt1td2rvn4QuuegwT9T3TBSJhQaNOqsOLyQyREtrpVpotL4gPi649N
VwSVn742NW4YB5r0LRi9E38Nebe69q7DcMr9MFZHSyIA2roJJIydWQq93+84
Un92yiZZhmFjBBTj7jkEfpsB3TJk2f5bsIkHVEQKOovVAK9cOypZhnleUk9o
OpXH6o2sSihW4t41mFvNX0m3bOs1RrrtR4MqEskf8vN3KUxDGUpcx6Wle5HE
rAgwv6qKocCsmrdpOcIhhJQVieRcM6FkJ+4Ij4jp3BKikUjkEwWygYvGMVRv
BXdSIHWSpVMenWxA58ixp6HwU0QB9QBZqMq+JGrInguh20bi7WP8cjadPxG0
A7PQ3vW3y7wwK2kG0HvAnevaSwMbJI3250mZPTeuIMAvhK7fnSKQSJ64vUvI
cfkL0vv26RRahixXuibQBa/DbHjVOtFV+DkurrLQeVJVvEIpZfFFqaAuiX7p
e2+ABmY1UiKeiluE+kwev3lRclZnom9vxbcBaxBA9rsItesrLhQPdHpUsK72
BEhwxeNdPJ0EMAupT3y/9g2AH3uQjRkgIFcUlulgB6VJwcgV+D3d20DH/+1Q
bSXXCLFWjOblDaVeK1pPUumuSiprG6/lD2fITSEkoXkPV3RMySiBKIWVOrbK
x/9SXg8tiCwW7Whp9gBcP1AbslknBxSd+s2aUOLreE6XzGhVhTQUCG6iA1We
IJJVWYptgPAa+W9zB8d6kBExWOqxb8laFqfTuviZLy4tngSkAtRyC95SNzCW
MnUIdTsDRk46hwwLe/phr8pBVZTUEnZV+v+G/KA0RxvClsmLuoak6zRYoGGb
Rx/5TnCcjxT7ep1J61u+idPnrWuGGF96ezQ7vkOIfd1WKGTsb7knFkN7C0Ul
jn5HnB0slDkXoVdtayLZq9ZZChvtG1ORe2Z2c0CzsYKUpZYHHCWtY8Y6zMGF
E4/Xs/LpqceIOrSaOyBks6EQOnngfbdKAYSy9QHaPUbkXOr+4EQiDNGEkudO
N7wgX+5bsHtxcr5ZiSpqp97GLL/ErEIUmkOcuB026dDnQosdUYONMEhNAciD
XZnM/AXwPv3U3JmiC7ERYbGCNkDSAdLHsgbTw781EjfEMIgmBauclJofrMjK
H8sUSJMS8GBYW0TTCua1HdN2A3bgvxipdjJM7LPovaJskm5bXR6Tykdy5Dye
v1uDmu9sc7I6vSDzxp2RINvbmi3Q17EbswcqTBOlAqrL5W+jBXzVU2PRUTsT
ViCMBSgAfq4lstn8lZBkUT0msc9lOLzsUQ0VckbZ2JMZsNezSCPPkYg4xFlB
WBdcRZ4HI1uaxJLcv7LJq3jmqvqR3Zd9uWp/tNZI+vlCx5YiuWFo9V3FNRTF
0PtoaZQV5BliMbHdGpOzdAw6stirkNUG1GljEwvURwQjn49wwP3MywXYdIFk
ZwSQaS0g87G1eJ77uaOpswg98ujOMRYtpL7hbcwEZlvRi0uSsnesbkvg1pED
eWOnJoxmCCc9qY0mfWtt8hCvsXWaDyWyRMCFaUo5uEdboNet0sA/Vl2wHKnH
aNaEjZaTBkMLKoVo+aH6ZlNDcto+uX+uPJQ2s5qxwUEzezYclDF2OWW9eJTl
eSTfiD7Lg2eHz7YZ4W0PMQ8V2V40f6vFCJ8lCSqEZsOi0hFKjUsKhk+0we6R
GsycaquZkmj2wNLNlYgu4WXeqJgRqtFjZlI3uonUuo2eQhpNsqBf0USc5KKg
QPqZlDHevZs5TJ5+34BMF5nT2Y0e14PiHJhQdJMErx+0OnQqk7Drx1x+CIbX
+Lv43WfELxvdIHDOqevqOT4fZzIKZPrfyye2kvC1r5Dlu1rmzxcyA3YY28Oy
8sFkcNTm+rQ7vKU3D/LNuWPaiKZTCFOwLO9HeJIJ0QPVdhIBeh+CRQ7ppVtb
HOaaDfF2ERvy8GbJVM48ENVkNQi5W8ghiEORgUSVeaYAG/aOPhn+xXp1QzzD
C4gsb/PDvcSVhhQhPKseGkX+6ktS2cd/4DQcAscm/R18hdYyoSe36M3NUJie
s+GLXWmSy3ar3mBt2XYKf6rIJRUFqbCh09L5AiPhwkDTddx3wKT/yPcc/3jU
wKZVNkIh9PRhmmiNLGPh8dv2omkC0LQYUMHE38nMelQDUfBfboBSiMgOco2R
2g8t0DNMgvZCL89FwKH5MddPWsiBd1vhRG6M84V2lNfM1zftShCzyVWdAuxT
3lV+1+11e8YGJESaUcA7IaA+splS/SUf4HpRBwwmZ4G/YT4tLDp4V3I9aFtC
jbxIABCW7/RAA+npQrSV+s5qMx81CbE32EzAdmWNsG9TKx6dEMK/Kz6zAV3b
lid29ibKEztmL65zGfYU0drpWhjBJA5TmPYqmz8sGk4yOFxOgkuZvxITckqH
DLnEFC3P61KkIYnbybP8+TT7ZmkmMCzTlfT31ec6aHyMqOZADmy7ctmozQn9
yJlJZRw0VA+fgx+QpFWZUvCEimHMSO70hq/uTSvEequd3oYnOOMyzxH0fpNg
JZoLqcMmF8Tz1ruZYZ+zjJ9E/Sy2/+hd+NrdrQ1IWl/v80/jNtEUeO4Cv7q0
e7C2MHnRSNQvSqpRCx3mzaOo+Th+N5Cjg9BBGtJKpbkeKxlNHA/9JYhgKvNr
oon4fZwa89zXdc1Reyaywcs2MevkbADlA140Hdvkx4Kc9MEZ9CuZ3UvW3WN4
rINyJtDARVRx2UJ4cCY+FqW4V30ya3jSmceVbjUgBOXrx+C1xrkVxdTGvMCc
sdkpvE4rdCd2R210g5+rzONO57cDexjAegrRnfwXDClqPS0bsqUGPeyG1rFB
9cfei+8izUlc+G9FR1QNi+ep+q9fWXC4Wb0YJsjfH19ehdwAV8xEsnah+PbO
wsmhgwcuyIs5BKF/AXKpGewkcN2QX0pBu0/dYFY56n4LHTlqFQ7REL4R4OxJ
8FuiZNd0LJXVoqHf9Gorh5P9PevIj2zkE2w6ZsXxgMzIz/0PNFpLfwzxmL37
+2Zuqr4p0refxL3u45RNAfpZ1tMD9+iB0+/RL+ygxLyk38Y7LbpuA+sq8yKC
p+YvhLezb9hC4ZnFbwnVd6EKROXjVlxkH8iHNFUJgt62/FdbWG38orn16kT6
EzD95qp9t92zSq9Zpf6F4OxMhvgXHHDxT9XIfthrY2grOIedIWv88mh3g6uN
MSYEFsz4QQOZfxNbGGnnQnA7p0uP+/72BE2SwG3ODT0DEcApwg3vpN/0uTG3
Ctoy2Swqr2zcQT5d8/yRPGexonYbDo0mJo62HZINaDBlebrvFoGRCzIy+wpy
t5WaiWDJ5CicvysAQ2Nn77kNlqpYqlWnpYb0xeyz30T16IuxRGp7aB42PRcc
kyQJOMkDfbYIYWJEUVLmPZh/hj5/54tzrfMUYF8MR4hXKYgvbIsEG4nAmC07
KthX6uKbF7oQ1Og+4sbIMR/DeIkwRu1oDpaZCSdbxKXy1fvnWs/WEoI9BFZq
spskyvf3dxjdF8DhrfFcB5CuCGxkJJ1zcbkzzlMHz6q+PtTk8O8ZaoJ79GsB
smXizhKuFWUmh4iIw1UdXdkVjhfQm2dYUPskqZ007LhpyMErSCgCKpqmebLa
AUiCs3oChckqLpmPFj16ZTpRAQ+8ho1I59v/q0QaMgB9v/lxl6RLDKWN4zYu
yA5ntHDWb6gslc9feCN6morUa6xosqmk10+ec3w4YlMutzdeFPgeaXhsh7m4
EjfjuiMK6AZ0sHuF5W/BCneel0xYcsNWSd3fwJVA86/DVCnLVxkirJ0w2+Yt
rIT4poSf2kX3T8YEQeGnLAY0lnh1BHHBOmxLYnCjztP9LMX8vazXRA4fq9JH
oGvzHdn/X2FLl0gPDwr0dW1GN/WZcNvH9V5aJ+IvGwhCKU5Hi/TnpoyPHVYF
5uAtQDixv7d0KuNApVoXEMvoHBcxyEM9q2FHkoziDNyfBFuXg4CAzxUeNObZ
KnQYWx7vSLLinThVDa2eQN67ZZRFILnztE4AbAew2XlDd9TAIjAFVUwG7HB2
Y5Bd0Hn4YnU/vVcN8TWLRkp981c+NYf34ZMcAu6Q3GCjyDDqcUjJKXhDTL61
VofetrXwToE8YcoNsZ7H4fHp+yy3jE2If7SRAt24pGkFAOHtmALd+7Xdnja7
Sc0oe33vvO8NN6aeCBfIczI8f2oyE+hYNdRXMsQWnE+66mquXPgvUHWd1en5
i/A0NiA102V3YcrxWHhS26W6QAVueiRY9HCH/4qXlRipDE23MgHZc0lpdY8l
e3Qeuy2Bdba7cu3H72lhWf+k1y1dSPJIdBuK1U1H20iDrnpoHec0fdGbvKMi
htl9FHXRvFAZNuAzKpYowYz2B7jZRaTcyizy1eNBPNHZBuq5bp4XulTM1zX9
eBaZcopjsV/tpK5+z/afElsWa9qos80p6gR00p8CA07bManxznqH9EWqHe6H
JF6yCEUvYywLpveYoL36BVBF9xQiAXT7xpW9hyDv/aWzhGbhszkEog+t/3Yi
Eq57MZJP2VTwfWK6bS65xHGuGGVZU97dBf/MNPqYvvVXWz2ucvf1q6box09k
DXakzPaOpU0CMHZDG3wodMG4jKV+MDv93bNXHWbR+rO+W/keoTuaYVf2n7cZ
TPNosuVhFPqAN4xGDjXMtpDqOgCGtc0f2poLVmlhhXiZ4J56WLSk3lemjeqd
sjX9yz2+uOPhsKXx8H1iJFtuooFvdo4g/vPH0Fg97G9aiE8LUiBDjynHpsT8
aQqF81BTwlKdd8627bet56wdgzt6WsiQWCemOrrWeggX5gwZDiGWSPGWPUt4
EpfqW+N9jrtmL2WUB7VW2wvBAZj0l1YNoknsX5VoGXUj+JHusr4LN3r7TfKJ
U1uO8Ig0bRvuC/xQxcYmYMf+SYCkp3GcxTYKRYGvHkh3EyL/UrTPUdxzysLM
CQzm7JTNcorHqVAU6tRiSM5tmSXdv1/EXMN3VxWQ+4A8hyKCbqpF0jfLT1XC
AMFQni4Z0YVjOFZWVxThbE2AxnQaxbYHdjg+ufLre6whKVPSeWDaq1n1HRd7
WrP5m9PSNELR56MC7hX52udCJ2yxiZmSUwXcuR520O8xbo8ziYYWY3fpdjDn
cEANEHHIfqZfZ/UM2Q/tMFt5ivxKLn7U+QK0bFnEjNdMYomuJjnyxGEjI0EQ
zK+a/JSRSnK92zsUF7e4EMGI6jrQ3cStnr7BltCDIoSOoj3fyJKz6oW4upvD
R5Nls6exAVP5EoEAdY3OgGvxxUN3p5GCrAz6MfOTp0zDOotDTYC27QPDZ+kW
CeOK98Y/ZkUPjlML5SwMs/EQ5eg2ZK7LNT2n78WmeHYGXw3qMY56i13JpWxe
7do0vy/qx3rAJmB26lT4ZJknbIsYO4C6gl+z9bNXHjw26pLxf2pNnD6eTXwc
65aXWr1YJZlMIOegMmi6L83VMQwJZbwakciifTVPoThkiQuyZIieDgJ9tkS9
XtszeGtNU+zCCGBby/ZV1y2DsiflLNj3prLWSU4ROnYii+bgHBO5Bb4XrYDm
jxw4oObDSynk7wizPvGDidp3/0c9/tp2QuIiDNuO0nq+H+mG89wctj2R3eGN
OoNaT98fGAtEX+bvbd64w+8c5Ov8kC1f43nQj4nxx6hqHDd3lMPXSpsnmTIm
2B/swORy9mGp7zVPdWcEY0kXl0atRxlV4XUIjZYXRJqJ/QOXmFT0EdrEx/BR
6GmNzvyeEIe72VmFOxfrUVu3vS09EHLRj6JFvMFgiLAUC7tk1N9bo46wlxuH
aoKACgqRscKEpS75pRt9jPxNgOQl2gtJRaFabfiNWRA1FC9FiIBPHccQnmBg
V9AUe1xTBHrPL52NCftScw1I98KArFU8urRmRCfqsLyAHyqGw8G7i0Thij5V
T4nzlzjPsCkrwcEQkb3jimjHltaZoSL72IvhU3M1XtOVwlTWcMTLXDyNHP4H
8dBzd6i6SI3kCeWEgS1ehWXBzh44f4THRKKrGlgwKrOQAxnX5VIAJqlhxQUb
FLmpmd0HnqiHja5i0Y0ZAe2mJGghTIFVCOoae+cHghZnFxtYCSIbRVlDQM9F
5PHiyIVB8NQqqA5iyOCBIOzPaA3MYD43RZprLVFdUTZ63Sp/VYycT0Mb8mwy
71vAp2Qf00srGEi3aqF1+SYpkRn+sGVTMhTRjHfH07N0CHh9ulrpcKJY/v8P
vHtzoduP3eo+6PudaH+nNbM2mMpDq78ymoB/ciUdzBbeRlOTPxtKhvdeA2KY
ZmIjC+RMf+M6gxm6TP1FmzBRjcPlTcnbPAV4CcPH6HCwuYYY9m4AEEjY+tAa
NsoqivlyG3Z8hj0oeSp0tFqKxLiLJ0EnfX+74xJEG8Z9aPFT00JaUwq45PvS
5YX2I/GU4RFbSSFUUtedrBS1fHDIL1OkiN+P5fSdm1EVgQWIVwqoMfU7jtp7
6kC0am2PfAhLJLS/PvQnY05xQ8e5aBU7k2x97Eh7zIWMb6rEidxov4nwkX18
Nmzsh6BvN+wrU+L9FFSgggMguvbCZ6VQkQWURH/APnD848UphCv/FoyCiOqo
EgYk6KY2xjgjPwJVULHdQsbFEs90/mIcEPCeC1uYRZQmkK/lvtBk8eQIgIxy
uC95qplFQ9LxWgVuLgmhdtL9Wqt+6FoJEx+ARyHVub0M7wZbQr8domSQdpZE
JfDsoD1xqJDetdzYFV3sr/Gku0iFw22dcli9ZeBNe/ROJvVWeCkK7AgR1W9J
+IgDKlRndjLgUmTV3jp0Hlo5Jb8CUe1+VaQ7Kug6jlxSxDwbTNmw27RhF+4y
lkQBF/T6AL8ZZRkVkr/ZIt/ByIMQobu4fPzxJxfpGg33YM98gjYkRxMjxi6B
uSwnez1No4XGDP80zhnyc5yZVJUc7OJmaPr5YNIStIchSqh2B4U6jbQSCB1x
kFJZqIYhEh3TC6sSmMwFi1gCNPKrxZXFOPvWyonZwHxYKoPxhFjsUq3rlpLY
Qn09KulDnwN3TOvuDams3rQP5+ffgsz530/DdG6Jmeu7Bp2hAq6aEL6WkJoC
2mSiHlOX3ZSto33NjGTNCPZO0X8+x3OEFBELygiukyuteztmIh0y/5x9niGw
fv325KZPPjUPaO61xREiUKYRUfv3tISFS5FdtdL1ttlbiAyhUKcOGMe7oUK4
UZdzsi1i0NhFCYDnWzoxRr3AZjRzbSI7zeYU/0YOLx1lhb24uGemkmEgB3B0
KLQNvuue9AGHxTKIazEHykXZE0x0SoNAAnVGWd07ywjUG2Woqe5eptl02hQV
9N3FbgnO3D1ZeoLmEteW93V53o6NwgInQoKQZRLWYHLCf7OdboOUHDEiPKam
pyHaql64PBEY38rDiZzYLQtcFE7fO4dQRCMxSHZrn0OoQsd88Xbmyb0xqvUJ
YSaW7m5FNn2f7ElauF5qVXLvsdTFwHQr2MgE1BjYa33ScVnHyrPUxfaBx8h6
tgiC9dNNQ2dz1HHGRdEBAPW1l+99+Lo7o5TaC0NA3Gqy5Xp1iQ1e1f48ZI2J
tdTrPcdIHO/hgOCPKok5i20bnvGFfjwypnFkAuRUAhkX0TV0Kg+HVbOKOBeM
T3AupE5egkseEl3TCPTMDiRkmDyakhUqE9tFAYreSWULx74YlpzdXwR3zyz4
0uSCL8XcvTMqhYjc3gilYTwGrBxmEGDJhvQrAQytEDYGci2rD+uKgLBYDkJr
4l3rLwT9++q5eMFEFmeOjfy8hRFpIm5YMf48Gks8WK17rJgTpMfFyzJ7ZVY1
7lLRv2vsOChalDkDvhxVbI5hF0mJgnsPKmWfGJ1gt6bPGnPWHYPGC8YRZt5W
3zfkDQDYe0O6geZTDyN20rK4HwhcGLIstya24DAvU7aym/vDdNcT1jQaymFo
bc4euSwAE7JxqlJYS9GAwBrEIz96n0K+SvlfXqLwxWrWFKUiC5iTVgncfHHO
8/HXcaoZH3Iya9fjNdJMLiq4smkkmbiSmeXAs8SfxehsCIV2YrhbQuqgO9jL
gkvgvvr9jqvCKwo4UqqoiRqyRUEMTkNKyk0nydWUz4Hly+wmGlq6Levgt3mw
R31VxWXmAblvcmNwcnHYv0mEuRpxnmk5FrkiEjcmD/2gUSaCXni3iZgPAyqF
1O/RU8XpeYhor3g3LzCNRPYMq0VGmSHu1wuMl5bLBm0H74qVdtsr3TN1slLO
F58VytDdz0X7AKBMx7TK9vqspxoDV4hzQcvdgsDCkzvf1k4BW0LGtE/r665n
BS7KNuX3KrU6yytPYCzkHI51DatiD4ABDZtFX9sRzdBhQYYC+6mNrGoRF+16
Gi7rbh4hs/FWEBJF9hkuN8K1WKhnq+0iwxF/4JM8x5sIGhk2e+kWXhrx+g9v
PWMF1kjM/4d0EYWFAtp8OhjaqPP647gPRKImXvrOZhRRELIWHNovZ7g9UQ+8
Act2tiYYE6wvno1Iph7G+73nBTyuE7gDsvD9WnKtLzKjcLbXdwUlMXHspXfR
yf191cgZac813b9jY/WXyVBK6Vuq+FavIRhc3/ZMCcf+awSKYTIfQsD4F2b2
WXmmChe3P9oeQCcxhbmD+D/Liu+oAUvjXn7zBybUbo7hYz8xdOzQ+C9LFAEO
n8z263nvHEAq2DCsjtYsbfMNVZH6qVQXD27JE1gWz1dJPmUXnuyU5Abq1Y8f
tUHNQCoAFGMGcS95ms9lRO7igc+e2vKkWcOW+EvGaFpijcIrmSFYwswYgaH9
Bn6zUBnM/GZV3D45ihjf7fbhJjQsLwaCtCAafZciV2abWdmXxK+WzPY8HhX8
/0tBJC0wmbW8yD0Q7nS19B1OoBdHgzPBK4PW6bYNuPcOBWvR9mmfLKk5M2NN
7YSYZwottCeztQqGNhgHLOuc/BVKABljdk47w11MCyKhtVSXrt+yFfbKYAXW
KbQbqZgijUpaKu/2sdMjD21fJTe0c7t0Axgy/7AkGfJfRQUsiLGLsbbiVug0
VVqrW9WyYcScP1OVSa7rrKOsb+njFAB6ZrfXIKb1YF+80O1X79JP8wR1g7xT
0nUGmPTkjVSFA2f1WA1bKIhV48bnD1s3WOsMCi0UnMI739mCACyHYWeUZnK7
Vfcw13F6AJ9L0Fvr01bSIpTTm9z3vsnnSVJMD5awVHBr+Aqv8fIj7UK+ojGs
7/Yf4LZEoVsHZZGvkRHSKuX0ugutTh6ItY5NfGZCxRo1nuIX9cW1Oq/HNUS6
+0OtSTmBH8ejlBKb344Zt/JkkQ8gT0YXfQJtP0/O2mwC9ALs52OAfPojwdbH
ikGE9rqBdtzUlSik76xDqUIzOveHRPZANzd6gGDy7drbnK2kVQiyBrT/CPT8
cx6KDlpixdm0E4yIMu2DkXdOGM1jzd9kpk0JZ3UgceWwcGrqxvq6NGtgYGhU
baJOlO9jzSTmcNxBTF7POnkQ7TL5SHkPkPpyMdz/tvm/oaCBtBThu6c61iU4
tf+QfNQNzIBy3Gr0VyvvZbnkkT831Vc4gIuF3mmHKfuE0c5ttPX141ZXzVq/
DN1IgqewVRvChz6MBVTW97oled0e0NLB+q4BFUaXPSBHRPI+TxyS6LtFPVbu
GrKcZDpn43biRfF1UYrYXkQNQsBSbxlNKLi4zLRhD/LoJ/3gLgMOuNZVDopU
BnCmi1rskw76f3mm3s2zSRezkeGfd7rrNiLrNHiFy344i3Il3Pi5CrUEq0FF
59fKdBBpTiAY83FuyXE+mAcnUOUy8EDBw9JaK63ytVMebX/IOTbW0GU504TP
oeCpGC0PE9x0Lw+PJntUheLJWwLJtStc9Ik5IzmtWRnMBgqiM9Y79U9V9rZ2
wpMG+fCPFxs8tE+txdSaeXGAP0BxxXMw/qdAa92Z2D/zIh300P3lIvel3dw2
AQSJts9oCIvw4AOPaNSOtxJD/4BDbacYYW09Nhia79l0J5ad+gK8cxCdZ8qu
tk71QHb2YgaW9PmKTUar1o55gC/kSpGwVzhpuOGHTKw0iqiNILXMWcwetXno
0RkzXEZ2F9QaAOmXNJNE8VKjqU7fIn9AsG8SKqMgsZJq6uVRwd+Vu5sm9RMu
ku4T6KxxWQqsyZ9wwyfH3Bqbrt3gvSHt+DFkHarhNPeZWPWo+yFwQD0vzwDm
ljUaOkbie6XCpBWKK5RfWMcdZL62RRKN6GrV0/mbKf2Ikb4xm5HjPKFz1BtU
fYbL6aGeqtb36lpgF8CnyOmz4jx/me7CEroxwChCpoBHzyxuHFcGL0dHDBay
VmZe0dhBuUZqqL4VKFsoMFSIwCB380lgYQtIOkDOgXajGXxStlA1FLMJ6TGI
RXbQLPiGsvIfIAY1Woe4hLl0CQkgzpZ8V8/bl6uWxz+f64HxBWqALVi+6kCB
q6PdOJ3pwyOPKCXz3tUs9QSnpVCtuH+CsM1MrMRZCXoPtSXjNHYwn3/1fFjw
hCgSdPzZtH8IS+/6eVvSM+nnWQiy308UME2O1TyYLkMHQ+plUNt3zI93x9jz
UZS4Br04Hqi5dpwC2XfI/yFeAZHwQQm/8citg/jweF+rDMEAsDeiIA/CAbS/
TrpqF1jlaVXr06l8GDZl+8rPpvqV60oPfjhA+8QlmaTU2xA/k8GaMyfaue0B
Ow15eTrfPPctyqxPiuHzw+0m+rdG+kde8JvzccMgTuZto6UvX6ZR7yhTUqjI
G/4L5dcaEV73HQVooVL3fccQNHrFmarUdnZLKdJa+se8FoJNcz1vMZdHD/QJ
xAu25hCih91vrrDwDyUukty6N+qoSR43y8Gbgo3zFlT2JffwQpno2JNMiQpX
31egmLpCo1SH26cCVA9sEwq3EybQDiVGNRYFKf1MoiO0NE3m+EwdG1pKZVJk
D4tE/4byr84TRrf8HGQrTpAQUyhs1EG/JzGJjxQNra1vMPaOaz4JNJRpZiyy
I2BJ8ex9htAx7H+CkPQue2UgLKhZzsi3Omb2LFitKjHhuWEPuy4lgL73y+AX
hFImuf/S4zaUtXhDyungI03H72WC0Ecz+mwbah6GpId6yP3RM7aBeSp9XmEP
ObCvpkvrmFaRT31HLAQjbYvdJVIZm/bd8QezZXYjdIYFVuWA19Ho7qpQZLbz
h+o/NqzUUmIV3/UyhIj7d4m9bZHvs6AjR9sOrpZbepLVsVenpe7hDLkBHQ5u
v3tqNfeLKqQxqdRfPRO2V8CDle/vyrAGmYnQh8K5Y9FN31btvVs2SK265woX
UBWYtbJBMnVe7hUDsjWgSj9K1DQJzqUsyDN/DF87+MQy8+yRX1xcrynMXCyv
vsnJylF8cK/zLSsz+qrVX4Ln4NHGD0qSCAwp/WMl6NTqihoL9/tza9ZzortN
qs4fBYu9EP8wVhP9NTl0e/q4tUnANTyVDuFUC8e12irVmWM3P1BNQKALxEng
swh+fOaK/Mm16lKpVsrO3iIz030x2zfFvTI3VJHTEjKhX5F0YdC9y9Azl7LX
/J1aNv1yqqBQJsk6LioWmzeomW+4VhkcMgB9qYxfBTpwGswPlPPajMJbq5Hu
Zi6e/QqmA9y0khHww6Nqyn//KnrqF5UnWKv4b/aYwlyA/WJMRJ1SiTo2plaw
gfkjCVxxEK/zFsBVrSPqI924E5cckMX02sUms7UP209ji6+grEXfS4AuAtmg
6q9B4MrQJWfZgkQ3X6fLDJZsaEYIZ/n7/XZmgetMU/GZazuA23sNTvJDx5Vg
PaObt9z4u6fnJNzhb21//Czfh59hlDKBDNkAMx0E4XkW+2OFlrp8GG3BtsoJ
gtmkVuyMz/glF3BvRfOr5uxBDdkTmjMZDuGib6DdTFgTep8qxpTnffx7p/X3
uPxgKnl+0tpH7UP3zKCQ4Gs4moiqzDhn6aaLk5xR/Rj1hJuDQTzRBcAPtz93
isnLBoztC3fllykDo+isknUZLBVLu9DqKtNjNY2gTowhdEALsok3dkwF5WYR
r6bsysky9v833cVV1ZNQ8sD8ZglHfvyvjS3ERNNRjS/4xxZ5EEm9HJZl2uUq
W9GLFjYtMan5yj/edPf/bzJnRWu/3NfErDFjqqpwZ1Ly7AlTYjZZjJjRYSHl
gTo2/KdzbNTaWZUe92QeSaY91XJ8bD/muQPuTSTSz7B02CeqXqlZqyDvK2Nx
H/YJcOTow4jTT2NEDKFDwOC05qPmsW3xBIiDBCxzgpvklJBIu6o/fdoT9bTj
RvvA+D0Vl9fHUUij/+EZi4VvtSRmZRHQwKR0cH6JrTXEgfT+0Y3DXHQpG+VA
j6/fpkBixmKJPtQy6FYCcjrkYyD1V1A9JfPgr0rWMPA/ZxNmmdac73bIZMhy
jlicSy3r7CTZOmZ1z0LVirTxqrCSuYH1ra5vmnuptO5SVu6PYBDgIa8flmcC
AdEg2Z4FsMA1w9h4nDxevRvwfgIWTgFJmJxXJWcV/T72DFjToVh7l3gMA59w
5ucA+2IFyY3ouyObmAoOm0EoxTFdi2mlaruXvbJdYdSKTu3wYvhRPwJyBsYc
+HJ52io8C3m9L2RNElaDr+xlpKI7c9FWaurtPup7DS3SCdOkQvQsCwFiDjYS
naJgc2EQEiJAtQ/Ta/XmO6/HzydpMIBqolycO1KTs6e974KMttplyPig5iOA
TloPnfnyIZnAaaJeRqfx86jdW5eazGzLDbvUo1BiP3dbSXIbdaF6RTka5LXm
RLCUZRmB+qneoTr6L68sTQNrz7+SBVfGmUsI4EyEPoXgsDWv6OHC7pMQHYG9
3G06lHocXyrsd1PVrf02udf0JyJsw5w+H/uJpw/FMcoykjJBWk7c6jr0ogYN
eGRqh2S+sc/FC7KUS111iiszvGe8sjuO2lU2caL1aBXXjFcmrMi/NKGciyXz
aPUKnzehXV3QrDih5xTk1xTJivNWKZAHYO6MPvM30q4Qk5/K47DJkC2RCMr4
UmJpx5tz8zanXx6Eu0WfhpbBgT2bL1iKzLVexXNw9Y06NPupwF9+av/9Xba+
+e6ZTn9+a2jOX4GsAOXU+roYhpdpv6ePD2/RQVcB6qyQ/C9/Xesu95CIfi/w
zrJ3f7O6hdgkcFBRYxRLJB8/3FptL0b/rXUEICOH5kL0XpBt37bawxQs0sqA
06xYiUuA4UAjTzaEHs+Ul+pvpBPC8c+mR7418ch2YZ0Kn8Lfvd9Nrqrx6oQ3
+QLZvZ/2iuYrXiglRsnTMaqnW27Twf/F7ZhD4BRlorpljuuU/Jg7g8JfLUVi
3jMBvTKVYCQAf2kzx2ex0tvlhfWFM6HYb6vOTvKmnr0BvJEPGowYfpy2fpfM
tJQTkarF7DxnkH56gxr0P5mCitfSZD+89FfpBUVJuRFZsa3yFgkpEdJJRPwr
01rnM+lV2sWKHX3WtFKBPGy4L8a2xXh9KiFGM5CHSjdE9pppXxJcn19KMGID
OJS1fS2ZdlEgRkQp3ado3SbGzYBO+hUdUIESvAsJZqXUTo/1hGD3rdSTjFdL
9+lMiq2fHDuHxFzlr0CjQJ4yRbqW96WDubRT4l+c/Qb9c3OjEOh8buqPvr+9
Dx201ZJ4PZ+yibtyloN5h0O7RPl70Rq4xopBOJaD4x2JR36pudPs0CfZz0Jb
5hkBTbzcZJbM5ftr4oeRtHmYNFlSbRUKClMvnvkmT8yoEe6iZeShz7v9d5oz
JeNPdW7phPV3JVxrpsdGM/LVgFc80Fhy4sKeGaqQx3EQF0RG0eHvPFgIcsGZ
IKgBz/hcuuP8l8pSeExZaNq/0Jb6Ga0mm3nHqGICKBl/s/bA4WIaFO9mifDq
4LjtR4s6/0hohmUulpvcjTpv7rEOkMBkrscj2sAjiwyye/qRRCNH9qbaltrz
v8pv8Zj6UhZiK580Goz4VYED530mzWS0GwVa9FHWURNiDukFql1B+wB+MnY2
YpXW+hHMFrniCjjqonNZcUDWH4SpZlRh4QhfI5aZrf1Yw4Mi6KxzbmmC8KPM
6+8WXN5Xr2Dn+YuFwUq58kTorRWpv13kcqtna3Czq02pDhdKuZQFYmLto8pv
Yzldqd4ehiMBteUblSqzDpsRfe4hiHe0kLOnDKq+taONonlSlBdaAgRvt7Wt
qgqEERa6TBhaJJ3jPVKh0iFKrFyE5dKhO5QiPjwjIfu45j9Fto9mSBGeqORh
kMhOz5ED3aSYDW7GjZ50dGhI/FbYnyPDAy/GDOYYiDY/EvF5dSxUGB36JEgR
B0w5bDRzzh9kV9nNDfN0zzsm0CbvqeuU7QSkMk1lEls3C6GQj7cVmxY1PPi7
Npo04DwX7ew6ZfVkurooqN9q8bURsvmHao5CJvArhJzCBkkwD+v1o4x6Iqgz
fV1ElMowZ20eK0388y9RT8PkCJJ/eIj8b3NGFb8bwQoBkcLrluSfVvCsc4LD
7yjKci1DivM8KHfw3DC150qIXOE5W2YEymgIrMf/sfysr2h3y5wOx4qwMugU
mGdQobhVgEGKBxl+h+zgDvSAf8Xv7L0uQdfmfmRF7540FjlDCdYB+lFsHZyQ
7LEvvDhTt6YaLK3nT/EC4x3odSwff6yJF12wbZ7MfS0ot+PK8a+GJeCmgt5J
hOHuMSF5GWh5LP7qOrnEytLbjtEwq6ifJizvBNJXARHDkl8eYCOUa1DE5jeZ
iRigChtIX5EmZUnc2PYz41zEy4b5cjqeoO9XDmw0ybyDtqA30bvsNJ3F7VpW
NK7CUdW5kFcvf7ldkXaGNiBRumQHnOQChtdvYSzsVa6Jhu5GrrBCL+/ZX24V
d6wUzb7g/UWymiPHHXzcNKyFqu6ZVvPmXXXajHQIubUqkhXuIvQgtiLBssob
fMrpiO6WcK2gTIaMEssP6zHBWreCxpayfSL1CoiIoOWrNmNCtugcfMge+gNm
NvEO6nRW/OyrrWLrZ19R2keLMI9cLGJZw3i58M9L8VfeotWNDySYiduewBlk
lrn7oddZT5FbIPDwoeeDN9hxu78w1Fql3tJpn0zh1akpPGPFymh4ssfYcYv4
swKo27PNQVS0otjFZbXsioAGp/a2GOQdh2v4vSQeAISaU7sDwQAeqayEfDCg
LhgpObo4MfFgaVMPVj0TknmNJCapyV35Kk2B1K/tYAIVi9/pQJ4boAlwPG8q
aGw+G0AdlJPIpqaQXlocRmG/+MT7xUXRQEzpgFAuHVDfGjJnQn59HI4QIM+U
mG7vxpDMKSCAUIdSNnngcbAsXK1ug1m/y6xCkioRnEzLmJS5IOVK6asoWp/K
fChLhVtEtcSOr1kwpbn95+tjbfUz+zpDRkTXPcw+286sEttm4mSSHYFkfA5B
g6ne0lis+Ab25+o+360ZqWi49drzv/Z9Kv+9ChwxaXhYTds5YFwMGIh914pJ
lXbcH43zulBhLqOp5QKhRruabsm5bMTWCv+k+K9bZ87mNNIuxwY14zlk9ziI
ipgR7pvaXLodejWM/yykIdZ4gc3Y0H1D9YGWweoQ2k5rdkwx9lwArOcDgSWU
TtmXi3Fe5Yn/FxHdv0+0a45CbHiL8CpVLCllZPJN3MScT1l5iEQqPMbxLZWJ
fYwkr5TpMsI282pSDxdk6WFjAHA8rjdZmsE2iKMvTqFcVmt6G2T9X6/LswGO
4ZeFd3kV5cP4RVJJg/7TC12aSd/g4rzcxMMushMB3EIV3yfnN06mOWYs/U67
E6t01kwZmPeJ4P/wI1gzug2EtDnPQ1koQaXLcySaDzTttTPIEko5J0A81SNR
EldGbbc/T0ctlW8WdGaT+haZ95C2BDawnVTIV/+B6050mwrHCYoqpEWhQTwn
lsb9hqKm8zcSS1wl5lAqNqAl1SUW4NvgBfDql1cyTYABPZXXuXwxBc6xRVIT
Nq4toeQMtADXXXb8sJzdEV6BpjTgtM+fMZjSn7zf0KaM41n3hV7ChbIyyM9c
t8MrzH54tUrV27ivhlseQRB5AA+20yYoFGf8IZVltv6C5affpmppunOiwDJO
CuI7WqZS/Db5R6EDvAlaMJKm4VksGE3q7Sr5wgreyyKud7YVZ61SRFfUu9/+
sOTJpLQViCK8ybZOfffbHiPKdvcrl7LCWvtWvvVDyHGXS8uLDVAIuTLdtP3P
NzVGKGNNRRPUp/Et98mssUbqGsCtBhj++1Xyrp70+Am25tHWOWimuj0ctGd7
X8/1Ftv4k8ixoafoGVebTrTKDGCu0nE07ZjTOHRsVS2yiWj3xDaPevgdtgSl
ZoVCxdViDDzF/F4mlIFF6/nVVFwyCnbM7siF8YZ16KxlXnbYZWEyr6ueMX0/
qv7MzlIEc0/alaiQqWGmBvqsuyQbqlGl790ClgG2LxOrL6TbkEl+dTVNqL52
Ceute7LsOoJaNmG2G9/Wit7TjUihkdkkfDEGAJpfpVJpyaTFL+d9cjNCRAM4
3hLP74qMogeHwjzr4IqED+LwscfjsCJPbbH/MPGlAAL4U0M/UnMG5SWBOwTh
ssx+Y2nswIkbA/j5hZhSMXfUoj7u/WPF11L6OoHjD8KyKroF5X/QCYhtLtgj
73IJoM1u3I3DHKEz+ttdGIfNX5c+6kq4irNXJHQkBzoDUdfsvkvLKrUxdD7k
K6qysaz/KLh27YUB9m40nNBMpNBUPFWT+yxpoa9ed6aWrwT0++lqK7kg2Ovd
2yBUaGCgpFRN3keyI5yqCuM+mpsIzbeBwnLWUHjlch1/zOo8j3WKfR9axc8r
YjE8iLzkJUoDFvV+48rvJKvOyNv9soRQlmY+krRJZtyZHH++Mr80zmUlp46D
2MadqOXTarO+e2IEQysSvHZmti1raX07l+3vpIEKqesaplP8wgw3JpNjExlg
k1xUtCdAAkvWImctv2VlMPMVB5jWUx5wO+ywbjoOEeT3oJ7maTNUzb1BgIJ8
QnvkXSPHWhT/mFAcZa4SgqlDPLGpGBMf2cqS1DuFPKaeH0OLMId8wtj7oFEC
F3Oab7lVmeRQE+rsjUhMBwYOj/morkFfr+8mTkTPekYHaakAKzsV63f4Zugn
7rkeFUw0Y5wjDI7xj9tBcqQ21NOMH6yzyYAIoVt12IVLxkXcS3eofR3oBiQA
QzTix0M/vnUlmUFWrgMXcjzaSJOIuZAsm8HVwUVakP08+5CqIXvjWYRpIL0H
EMMgPWzlKEuiDpSKtMywLzn1hVg79WX/zb/pGAubh9/43vesdkGhciDpKbrm
HPjOMqluWeF+tA68hOhMh41scf20odEbRYf5FJsxpguS9PHm9k8v5kvgHv+T
aBTqUMScFVcyGD4jPb2tQ22WlWi6hCzGFjKePJ2fBsiAYhZDCLb91k/R8Sss
7NrGF+0XytcaT5uJ4lZJX1KbDRXhdJOM1meb0wFmuEcMAXGpztFtWm9Pvrtx
7IMNp/YIv2tdDd1EoXmzVdJ7Et9nOhjHVzhQyubl20mjfk+J5JbUO9hBGNVN
8OVSM7T/PMQQGLgGXUSnyXuIvjAAuuU+jRv4a8Ow/05ISIhV4WuuYeUX0A5V
BxvasmqcgoDz60SvGXl828bQc5Ti2i4HFAJEiXJ2AZjvVu55PjMe2jKWPVXk
fjn0gyspKsFNa8EcymFujuq2JhUq7pqrZIHnbmzfQF2KOmdLq9EY7hoRceF5
G0Z9gbLZver+8kXtysYA/c/mqFe3Cy6EvTMu6FhTS7szT5+/ulH5b/UwET2P
jxXOALQpJKtMAAVZq5facGXP35udJqLa3pLcEvcpolKdWK+YDfwdHjpW6p7b
usjO4wAeXR9bDASuhObh1M81AOt8JyOFSxTWecX2hMgdqffKiGxcIc/cFclO
75wbP1ZmRZvTRkEICYHJluM8xxjVLuILPL1eL41oMgsickwBzbo6AKL541lI
cax6827Mtnxo+g1eJ0U2hMLyDcz9N5IBcTRvOE+9xvTiBOAA8RWLUMcsOE2Q
9CvkuM7DVIgy+uFYOeL53fEOfT+cG7bfhV6otsx58G+Pum8eMJ6Nspym72po
YyZQgfOqOJBDmlk7YpMoIbtB39sXOonlY67Po5UJfwIiFYFY/s3xK35NT0+x
DC6eAAzDYc3Tx15llpvyJ6dW4QGGAJCPdZTKJZoKZT2DjZReWd6bu918TXSa
G9S60jYutjSPQ4RzQq7v77JFKKlAprv837wp3PSE8S9TNSriMOMoPbR6lshC
QKyowb5sSlUZK4xIkn4+9x2cDYCWfGmrYEZdPiy1vlNEPEurltlujI9C+BhN
aaRqMdoKsXKkAhD2im8X/Vijhq0eacsy+xL7PLE57RKkaDhRT0oEQ2mUXw5O
O/Yb0Ww28X+jc9GtT0zyoDq3k+NqJSh4xeMFnAZpI+nIctUkQ2P0bd2rkt5M
HKGPvnlBl/q+piQAccIxV/25CEsiRYcWJoOHvOB3m6IsXKmIjH9rs3VfKaJn
Ri+clboCAiFFIbrsi/WEFLMw2uxb15zHQqJb5ssqbIPhKrabquecMQDsfoA/
lUf1lsS9MLKp1pyyskPsO9n9YtXTJO3NDG+HUExDGIehHvD97o5StnvU6ZV0
rMAPgd0SY3HyIxiKsC8e9DRxE+j1EJZdeWsR9sKfzeDyVgi3zGxSuL6wieBV
oHnc3aEMEAAeZ/0dVnWPcpxnR9VR0C/Za0qabufRNqjHSPSK4YbjYlumMjep
aFhBUKjQDxqZ26axjaykmK6Q93vDSdaKkCM72BjhRom1MO7Ciej6XxQJWhVN
heXKv0TiDf6BkMr40yk6DcgMPtdcWRNUGrcCqbaOvcdBMWKRP3ND7xfrRXb0
TnKxAzcuBy37Wfz+S7uNHIULAfu4ssP4OQzhmNQbwWgPbLnaaPhXpfWGN6Vw
pcwUcr6SBJsf0kcmN+c7hq8h9vd1AKAF1+KyLKAp/ym1vX6sc7BlKKRXXZlU
5rllB3bCLtC5h06a6ZDcz+mp9k96GBtk/JV/2FVotakFL9pdlKGHpEkC1gIk
IV/AGJ1bMvPKiiUBTH+pOZ/U/uUTt/hQUgQ3hoB4yN3x636mrI43CaulDiU+
8yMJoJTu5k16mKubwgd+bpuuvr4I3MiYAddNGl3b0q9y4qo6FWVspmAmWp/I
mqbMFFJZkfNs/4gta5jNOmzlC6HhvaAb/J0p7cpojcNhJz5eCG8TKFHstSWv
EJ3Fl+SEg6AvesAF6Rp/ggGryKt0Er+dVWh6XJW1WFuxVdYyymnN/gsme4lX
OL995IXAbd5SXRFLODHaSkYl+arHnQvFuhZADaOYzNEoHT+eI+Tvakx1K8CM
P6TU/gVNyjf43jjjaORZolrrcCeb1yczgd6/zrLltr6sczPKOXZI619mSFla
mbEwyWWbm4PgYx/eQq+5GfOr40OyiSywBGpgg+0z8naVFwmDegVe2MYA8W0e
9058TPW/ciKwI/v+lzDuEoJ1EnuOKEiX7b3sfqm/7XIai8kUTvUz+okfibfW
YsBZ7Hdr1475ufGAT5Gny3S4Js4rbVegcBe7hvT+mvJHP147buXq1Kap/coo
bAa7GUlmeaLnf3Xj7miwweZupHQsHHNZAXj7xqIHY5DJvo7jL6VdOn0DQb3Y
T7tXkW02AWhCb6irl7aitodJdVBIJWc8SoNe+fRRwoX+ghGVa/JDAGMISzGl
bMsp1TjdKs3VGSzSyF1mDG4tDVC55mjXkYV4SdFV9t9YGnp1WDgPkRQ7V3/9
hMi1oqDavi1Mydo60YnXVE51imM470pUGePJwfco0pGXcmckA9mUFgp2Kvsi
huZaF3cSD8ECbpJ7iCcDELsFUxJ7IS17yEd5r8/JNAfz1W0a56HLHgDcIzzw
wX1sVjsKnwej4atwsIitTKAphWjShP+nJrP7i876QEe8N5bLti2H0aR9waAJ
M6yDFAapv5aVKhhM2IDucsfevr01R07l6ojTK3Vo1UFTWeGSX6sDLi+7V6R/
MKWxUecCclldhlA7cKZdkVoFasP2tqVM1KsWK+B8+ZXfuzMu/XI48qUjT/e3
yWtZ27857a73dQhkGu5BsQPcE/568mBYjdtycC7hYzgCCWIElI9ab4uNIKCU
EH5KMRyquEtJK3Xghu4u0pU/jF1fUz+C0LIfk3D5V4zexYIUWIk/8AgwjRNR
89x/lZW7qmh75IiHyi/xV4IGBFbZyi70WGmjITCZQvhYw70yoyBTys8S+1L2
ZOmTBfv+fH66G+PrvFtfYTtVI+/rpYB9lrsENAHHyv5EOj9XD33oUIE20+mZ
iicE7PF/2KllUMbut2Up5tjxKCmWgEUVX4LX181A41LOnKZ+eyx7HDZzUe+1
SVqb0ImhIjBWZxic4yIUBQARpwGSqrK21Ifsk3l6e+npEVhO67xDFas1/9Ep
Q8AZhbHX2Aq8vmuwEdAZCku6pOFmS27/2/DSBYcgnSY4536GWIJSwL/upWTV
GKnxIrWxs5U/ZSNbDP9qwZZ9ymls/dWJuzEAB5GliSiG0K/hzcoRSayM1HhL
kd5v89YOT60UqhoLPFzltcQBxo7OHzbOhsLobkVUg33ilm7ETTuhOGDae4tg
WfbYVy7ZxWul9XvHJVWL2oRQPcIh6a/0Jl0xIyFp+l9UqcQ7hBkj306T7fGM
HgZBdyc7rOEjiD5xOmzZ2myb/hF0yOxRHA8Kv8RTEvLJkszizUMUv8oieSs3
8xWYgu8iLUUwlWdgyhdaYTmmCppTZQT0//eQo+iLQ6p71oTmX3EmBHp7GTfV
3HK98N2RW2YOW+nIC9qlGXsD6YuACkdOdyXnHaGI4dUT+KDZDRjnvmoqerlC
xtcGfGqXoQYjZdYj9C8nJ6yjbrJSRh6I8WgyIDHOlZi1D5s25KvwEmz++v1R
cEPV5AKxPsfdV0hEdssgqhAnsZd0IKp9OmgWqYGl33ncsOVGjb8wWJe572eo
8gPZ7Xz14OifHZP1HsTPrbhc2CttH9OvW6tHVTgXKh1DP2JyQZlG8zoBUz0N
7t2aAg1zm/q0LM9gBxDQtGnpxIREgFV2wN0dVQsuLWsLkXxXR9IcAPjIDQj+
LfqX/ALd1cyFzuAcshPE7FjWjZVK97nE04rgdeVnh8fbO8muflXuGC4zw0Db
bNQUck9xoeMlIFcM8ej7/Kchm6eZ+n4dz5CpyetBDWbD8C/fHUQyHHavEuX9
vK+2M3vorZe0WjGFe+ZMfauEbTZ/dgLSWGIycseDXazxgTX4hJz1GgIO8Mwp
HIdpGf2cHD/ynZDxvYqRa3ho7OUFzoYfxxTwODQzJOFuKVnay7bjs4pq98wz
1i+srNA/dyMCqgiYIYOw6LWAkfiXKeE/cP/BSH4os/ouhEOZxfnXeWKGpri3
m0VcAMJGcO2W+KHwewBeYRvbTiHb+nvc8Cju2wNeCQZz7xCTv1Y95xAh+5RF
BcwRvHbuil/x7zwCC/RQgOQqSrwaay08B4zNMHSZaOlpTd1jXe2hYhE778he
ZrAL/WrixUePagcGchxhC6XtnLMX7enRIzj/2t/Hy/ft8DjElP6lL3I/NDse
5WQ0FgUr1K4iariFJVfwT53lQkSYPXET6TBdoIL31l6pGZEPjFm8GpKidATk
TuIz1AXONkJTozPX9uMxcxmD4XGktmPGLuULvCpA0w0svnD91m7EtsaFoKnr
mq/E6OhR+yfRj6PP8qn8+/iMSd9cxSOAxs1mmQP7fk9fIdcXFutzpB4HYiCY
FOI21L6np4hp5wMo0xOHs4lmnkDEsPsAbQE6hmEfDTF9MORrMrhoGN9pGgwC
2rX7PPx4WtPFP7dGcv34xDuuNTx+j416rHt2SnLhlXWhcf1wB3wpDdcR5t6n
C9bMIxAxgp1O45L8otNWRe0YpKQGsD2Ix4KIEaVn6YlvO2gNzbhBnLIvBGfo
jVDrSb7vXXoUu9rdNrgbQbAoknCzw0c1+LeruBpQHCELxsbvBkhy9TJEsVBA
wK/OGPRxrwRKqoqlk1kqZmQsDZ/7kPALbC+GCouovHmZuY5b2OnASnxt3jK7
W1/ugZZzXt7+yyKvk2BIWbK3gltTXr7Y08WNBwc5nCbHkjcT4yd9mE7Zx1m3
YnAFFwyctAKC+cGeCJlnLEtf84K/Fa97p3k+k7E6eyn3ADnhAn/itS2zKlGb
8tQ8VM7TaAYZx9XvPTh81G5jVmMvyXTYD/f4LXB+03ODhTCr1bzvJf9EwTNi
S8d9MPJkvuj78FM3pNPPRFov7KHwk/jhlfEJrRPsVlClTS5WGhB23RaazlCL
5X5PhLoLO9+1jDS3QeXh5IWv1ZrT4u3dvrU6JLNlrNMHmXmQFsxoo+nifBWY
cQiqgLomlsxVmrDSfMO9cJ7KK/d5HQ/mXUqauPHgReTocA9+pOJSUutLt+Z0
qtxUsH3OqFP77p6xm3h8bkxDXDl6sfVcvS6nJftgQjVO/aEMCJQ5BFVawdqB
bjJd7/l26HwoS9lNVZyG5+PwmffqUfLCd9WDWHSXfUOXW0HaTgXsmuPgHY9G
mRlhgPBoT2FptOliZv+y8Otxztv5/Mnk9kdf4Nl34nVMGg5KOiS8YWlwN/Gq
NAAMTqNIPUMwCqqx8rDUchs6rlJcVbGf8LyhOmrZLGtotiGzTIgWJrOEdetE
jEb1GWwbpPPBYUhOnlmN/8jtZLWejdHerQboKyozAWlh+f4q/EhxOk6Zc8ND
IOV5rjeXn6dA1/ocGOn7PS/TqoGC1UP/VOYjd6zj2HdhPwHEZYPmn+itnoJf
5N31+GD7nyECHx3IoLDVWCa8gJk0biwunSGGfWH//rnkvl2GKtWIkQRyBGtT
vkjDeqftPjNoJnkjHlk6OAS25n/LAzixDAdlrMeu0pA6UoY48pbn/F6dnMZ9
1RBdFKT7ETv7HcLtrh0iVRBzh73y5BP/fpvOwZCfQYOFviRndP0gv9LgwJuW
Y4shoX6CJaUPsBOQBdGIOwyoUEKzkFBsRmvh4BkN4Lbj/mGxCe1MRq1E9IAK
5q5MzK0oOTYkykyq4IQfJZ5ClGmmaXdaWOnoa9HC9aAo+e25YNCZNYet5QYc
d9/bvgeZL6ngBiyPiaEcTbMal02sw/tBaMckKg+zCA3u814L9ZbH3rEeTKcu
940+iEJc/vKI2UhXLE3UxNISs7f+ijLBkr96Qf1nv/Rs32f9cvyN09SlSPBv
pXkdL/E2/QLjPtuCewm+5TOl5xEzPIUWeYMhi+kHzdrmoc3yGgRINir74qEc
UWCv6FbGdDBsnp3qJWknsfOYYZJRAFoTQ0/yCoFoN4IaOGJNJetyHhbPRE5d
peAbXKomPF4ijqbuFJ2Lddr8ueE/ybdIgEwblRPIoTLrrpv9KHjXOEDkO+Ys
+lIDuIGtJ/N8kGH9YlxXE+a8luxzzCpOjqT9brrOUvnGlKKJkZGq6JB82Dzx
l0k3BVy1s6wxc1eqm771m3eQB6sScFFE21sOI7z3NCVQ5uZYzMqdWXZBbjmc
/yJaV6VoDv8R1Kr4r5VbYTOsPk5B/+LU1kGa/8mueraFiKvwadmWYktz2IOF
r0ME/ESTs13Gn/3wyIm5UmH6ILl50CVB+5oL7qsgGZoHDQp4s29gRUXQAZPi
wJfOFVw+3VVvpvJgB2X+SQT/HKkradPLwF39SH3cJX+m6AwiD87B6eeBty7/
/Uta8w9FbrfRui3W+0+qbZwWdrQiRqvKdjf+R9+h6wDiHtDg/AzaUrj+mDTt
wUsu7+rNiksim4UhfW+XiOBe9wArpBiIyLwlXzAQCRD67tchxtG0HYJWDeuq
0ShgQj+AWLHLQgqMX/lCODXx8RRgqZ+5Pn8cFgKcIRwe17zaDhD8ayI6xfz7
j5p8G0VNRkVJP1FBsZrbUmRAlxmxd7YF1rxurNVavW79UwMC5FYt5ZxUrEF1
V3yhra7UMANAaApEi/a6ZvJ80X0EQfRT1FOYv3qEsBiTxELho764tIvJOqUI
Aj/fRkPtKrKtSh/IAPwlBTArev4TJQ2vHcCIUwOoAdzbsVXgMqQPdHkmUqMK
FL09M6tNypyI/Et4gCGLBEC6mJFHoMhXu7XsO6UnICFtTIMbPMupfHGMDnVq
3YFDvoO+7Y9V9Qv902jmHilPQ4KavTkgIJVx5ZhZbX1AfcuMDukEFetHUSQT
ggWE5FVmtcycK+nZADcglmPckir5ymA6ZIhOluCBNO+vq43NTe+xs8rIcVfj
qmGcjxXdCTcQAKx793p9duYHz+T2Si3Dt4VJCeX5aLWlnvCVZF6sJwF2DkV9
0q0d6oNzPknTwrSVMGikPFk+Wrq6tyjcy+t9u7Qd+jL2f8Yi1c1iiVbSEM5I
ddz4zWX2O3dqhoid7fDGPQa9illOA51QSg4EEAKS3q9PV3XBFhhIXXM8WVJY
+vHo5qKOgYDZ8OQMp0w0691R8jTvpZZI+5CSsuNPZsIFtDmAH+CTsmiBVLAV
Ceg1C7LmZCA9gdfuK+TVm+eeuAYV6KiCGhysyygQ2Pmux/EnUASJ+hLzbgFN
mX1J0lcP87B2t/mrhoyveuIyXNoHAexn/1DCNHYzpmWfQldVI/xe/89ES6u4
M5UVfk3HhKxJb0H6ZbmjQgTzkJ8NEokO1CgaLwj/U+aj/ZU2i6hrEnTMTDDQ
wf4Lsjp2mBsopJKQPgXu+dTVE1cwK3ent3t4h9+Z+IrdveOlIFUKj5w05boC
a4aGWB7mrtYHnja/qzyP+9atrwJ2HWBd/mGgpAdLSx6axUm5FOLVGK67i1h9
hUvVsRuW42ZuwjaayFDAccLVgPcCuMoPQcariQSF+Jbgy3Btjr6lYW1kQwg2
0P9yLr+1jUwaBLPHPvyBOkDhfPpPZIRLWs/Ag4HjfGJegm6eY/ky/4gMwgS/
o6J9Lqj4ba40QxRac399DnmVHCUnD+a2gTTKkGnhuB4rMwvh6v4WB2YFtmlF
fB4Q09d1gDMQxP+KIG4TfNHzR3m5CReB2q1VhE29QncFLL0uzKsJoHPwjgJC
YcFLu8kkbQGZZptHIv3UZpbdiVLjBVZRqy9hu3Bxs5T4oAEFUSIe7ThQTIk8
+XZSA6H+AKSWelOUZrnP05p+FRJT+V/1X4I8XNH7NvJuCp3S+lHV8+JObEhR
tfr6Ad2mlwREq0a+49JcaQftQ49pK/PmLP7131GETPE7OxdL6M3O4hT8GBHa
doQS3fwq6m81itP4zw51z4R0Txf8cfbkuQ2YUD1KPMqmUumY5IhQNk61GOET
RTK+aYAgLbCvrpROEu0C2pWRwBT37OaiatWUDrBQKPe3I7sELT9uQDTXdwnH
Nk3h/Mr/iKfjoDnarJ5TRQ707Q4vXx2BIBcSPxy0i4b2COxj4GeP5armHxOA
Sn6fWGH+bgmomS5vEGUIhOIl+c0im/UWWShq/gXVs9j8c8SRcC6k4OarVc7D
DHu48Zwp041Pvb0TIJWUIXBmSkdqXYtFUHzb2lKADaGp9Bx6Y+ng3USS/8bT
kUayrX3rIpXDm3jJnHXlEoQDB1lKTEfqWnFnTszpyl7kxeQ+GdwIUOMzKdhs
CCV3h7MF+Nlnd61mQbuIS29gb/WGAKwi+aKBTiU1ZV9Py/s3a/OOtT7ZaqxN
rAlLYdp9xLRBI4uuDZ6hfFWqGpEYRGVGY0EYdpAOjy6cQ3KlBj7i9GR/NCuc
Fsd4EmGW1wIOmPOXDmdvEzqMrAjbCH9uRQMkJ1eoOuJqv6cQCVjcHIMKFNBH
uI0KadnDB9USdTCeJYQ8MfcLw+7alpRonpEOJZvHFrFM3M8VXWj/ujoVmWTW
GRde3mifQtxzqVl461VNG4Hjy/YRWniuXDRbQ0Zvw2FVLrNL4OHjWMFGdt+R
3hVWYblGIqCa2PZkNSx2Oo0cOetdEYGOYThaWso6k1N0+0Dfha8+oJqUP/3J
FklgeI9Tcrp0zty9tl/i5ewb8EwiyzTUg/ewRC1nYUfKsXh+N4WLN5GvChl7
tYdZ4OuQZDb5pAb7unotV/zoGKSFgXm3PIUHm6rJRsybXKw2gaW0S+mJ4GKY
57K8W2AoWefZHX4EWxeEHxLl5bV91chReBsRVwm7tS2k+PWdrIlljj3kiz7t
6UrW+By8ydbSrSFkNCjMelg8G9ZBXeG8zLvhoyLFgzuOdpHQHVeMdAQL4pQu
kKT1Qd4RomyVoX30fM3iGoeneU4yg1yS+igHr60Kfex9EzfnPEKY81v2ZWQg
nefQVsmLu7HgPuQC7eyIg9zX425Y460jQTynNy5acH+hoJEM5U0vBujUWAzV
mfN6wsTTLGIzMLHOIiwE8lFKeoSzyDj028YEtCUNdiALHq9HCDGQp2cv/cvy
N2ISbXXnGkuyuidVGNRfWEH5CmeR/j2lc8eTwTNSbgRbmHKWvUkoDziKVuZv
hUCQvxLi6b1o+o/7W9N2QLHCn1072kzW88hEQ3qjzBR36Jma1k7Oj/rayWk6
ZkHc4xL9qDqE1GJMum1a2+g4wk4YBaRP+twbt9Psu+TeI1uo5UlcRBrr1Tso
RRFTbHYqPy3arHJj7s4UtS5q89GJ5nCtyiHEPrWSRYJLDGBNBim8afYPcWCD
p0Bsm/w9MonP4ee2ttp9u9I0ZuULYiSJK/62fWHnRCEdNltCBpK5iDHBF/rg
zG3rO8SzPRLimVJuuafOFSVNdGDPutZdxwKR24+G0HwWvxKZvtqIBMOc1pfJ
l8Asbm5AHqYr0rq7SwBos5FN749/Oq/SspsBvoXL4d3TZGZyCP+pu2JaCK7F
R+287q0OprXuSsF5C8QA7CHdD++D8OP1Vb2PsSeFyq8DYrSPf3E7/XpFLp3G
B230N3JzPNoGEzwn/j9txsDrZKf2YTD4D4+v8Y0Q2teiSZwGpB6h7k3oYYUf
EVHIV+h5PTwia8IxXV4mNWsw/BvyGyghcYtKGuXtk1C5/MVi+5ZDzg2ljynC
8x0cIyp0PvXBRriJGfP0lNITaGzbsPhKu19MLgeGu58uaRgqhViecIGsWQ1x
wgbixLvUJYeOrSgj/Cm21hrDUyBB55apiaZ+tJ2bI7o79DRMdAiyNgo3hFox
5Udg3T1FK8TtwTvaAfjhBsue4TS1Mvk9sG0vHnf0Q7cJWywdu4XRX2ijSU4z
XWMhDrmFLyANQMSaf/qKh2LSezUUidpXeJII1ImOEdGtZNYjOCpBLxpFvF8+
s1viFvK5rvCEJkHii3JMU99ogmu+GWqEB0OUCAMq2Fi0db2OgzmAkWZMaLQ9
rpbGH+wC/k3t4fr8wFK6RWgVqBU558joPg12qzuXDycJ665X63+YRDLyb6JF
90XrTqv7dGLdgfG7cASpJUU0U7guQ0Im8Elb2bPieOlrmLtiS9e6PsqmsCG4
7SgqIVZlj9FLb5pPjG1ELUCbDLTtSjbkDKLufWSCo+LVLPRUqhk2jwkTgl21
6PIlet4f9rr3xIJX9tTaHrl5rcJPa+OV5bMEr1Tjr7DlYRjhxm8xaTfdsLBo
zbOrSKVC80wiQTKDI4ZQE0jGKClnj9d+aj+A2r92Dgc7oZqG+8FkAkTRVGSo
C4UFi8ZIQ5hzfgZCb/beAIx6+74GLU6G4pGBHg0wLmGBBBP6Gi69eLKGqGah
0forHuzCv5ln9oGdyrcCXPpPmIy1vAhav3mnmp5yY68M7s9MF4KFreEJH/hY
LXD99Ci/tvNKr9BWnyxXeSYyye9jUCMOZSPL9OWTgtR+sA4S8Bwn76eQlcaf
+qLc3Q+3Vy72qndLLgFFb8LzrjfZwtwMVDDxDgo4MWHOy1sFFUwl8b4Wxhzv
JpxNknhdK7WcFNQQ+x2ztdNyblkIUmL4BvHzvgBXSQAJ663VXdUtoaHKIbZy
defMvOwRyBCDTq0kAseinXSSM+A0uT3dwjAY+grcoIiEFU+9uG+0yWzuTEzd
4yWEMJudLJlkfgRlRgQZAeMMSD95l23ivIFJOyWU4VHfAnMD94Z04bO3CrVu
9uPVzpyqYeXpQ2pyxUhEGAfiISWr2JraAUpQ8KBuyp04aWWPuH0bJBWqffDx
BoLjzr18+paJsFjnK/mMrjB1DUTm2xdmWT8fRJirpee2xzC46+9S1TyTXpBL
Gvu98oHg99ilP2N5lLu3nsgLYlmE3oDWllf+GO3yxQkS4uE8TRYCaHOkeG26
vpEatMNzQRZqaVrIqsXmTU37xUnhDH7rYBNexDyzCBJ5epOGkdxE/KqdeMCr
5kMTpKR3q2faoe5k0nplnLDeP91ANUvdBbE6y4IHZHpp5WlCrKJMVuDd3PgR
99k/g6MGbvFZze6TnYfGr/2eos68wvUW+GCT0Z67y67Y4Ff3v1J6d0r4YsMZ
Hdwvc6mPbeBFs6HnuVfEs5Dl/d+Dq1i4lcs91qelMePd5Aj7PYnC/Ypze13s
F9lRtAt+KEy4+RPNDRuE4qRaEdvwsE3hG3yBw0p/LltB8kzGPvkU34SrIAoR
dOU+w/iobN5s0H8LepNR3KKpqlWptIbEBWHoBEBtz262Xnbd/o2MUEHyHMML
0Juz1PlLYBfUlqozQrQyS6ReFH/fZQltjz4VFoF9P5o22Xmxp8wSCTd/DGbe
s3Kz4vnAA7lJxSlHKcCuZ5ECPrZO88DlINwNyxl20kgC9oxCwg72KS+CpCZx
uaWrXu0rvxv0MU8nIma77MMnwEy3V/8wpvj8BHe37ALSMepT/ZCuoKBgbI+x
yW5XQ0BLCS6XSeZQfExNsIsE3qDN//LXymRtO5ZfYEAyn4hy2O3b+MBP0QgV
LkGcet3LIqyVB0YFpbjfyVUESyI14I4dFfbgp5DFbrW4s09C98Mehbkxw4Vc
SAGPc5w9dbgt+Yxtk+/S9aR6hoXO5tB/pzhjRkL0aXLEFLwIFoyk3sUHKqxZ
9pQUUPfK8z0g3+W2Lse67BbxtTawJHXd35ukfC2Xa7szAYdcl1gj3F3MB90+
m447OKPpSdzpLShGjnq/UhDsKzoJJ94fhSMb/CHBCBi7rpRph3Kk5f847h5A
xTsxRtUND7eLuynG7lLOF6Tq7oMlPfjgl5vP2j4cg6KzoQ9J9JivUlbUK41W
s0oDT0zq/yAqSPEbiiH3pIYVeccnQSppmFQDI/KYKyrbhH23As9ODxQEpNMJ
X8D7Dj5td+PRQr/xE+ZH2XGOdMoZLmFBXNPV3oT8aIe87L9dYwNfNHKFU2bJ
vRV9POEEIvepO074lko6Ma2Ba3L6wDdoihIw1llkyqjI0mHCQZkU4ZHv3HMc
AeDhT9gqGvJY/R2IiRc3mM+Zk8nvJBD6D9SQM7oqfJi3k8oWqqgqYEVNs1TL
4FBQ0g/QdgmqdcQv6CBfPXVupW6iUSj/KSgOuKIp76xDzzQLW73Dx9Fos1k7
waxe07xgcjsaCDUO0tTNQhJAKYXWWY555sBYODS7qoYpnSY4H4bY8Y3FfQAN
UNHjuI5bYNXBrGip2ulHGdG8itKiE4PBo8t4+SvVVroAwB9Fk5MQpc9+YXiM
jM/u4fbXB8z1ds8VEnyscgK1EpC6b/J8kQTE7EnvY5ju/VpR0ORvTNhiiDdE
YwaxyeObFjYd1f+z6Rd6JxfsAPcAgxxE7ktAPjjrklJOrBUwvoJoLApTtpm1
y/RW25WUMy5+RdOXasmIzTUB2ifiW74GAR1Yf2NoBrnWEFZj/F934V8AVhRq
AGZ3BEt/tP4NxMF1asnmghhGFDo36Ia2OFeSYhUFVEJjUuNXB98vYp4e3ByQ
L9xcxkcFqhhxtmkcsskdOMR1lHLKbDK7o5mH6BtlLhJaSBXoi0gH9FGmrBx0
jBXZo8PAWI7mjDs43w9gDd+E2XmLNEX06SotCcM6uVO/kCKEkb55T+cCywLf
S+EvVYwqVdWNCul3ArvJr+brv4fx6lTcPhYXcBn+g4SkvjUjcLvqEl0QeUpf
4BtDu00fwGC+Gndn1tUw+nMBcbbxouucnsZQSKhIzvoqdTLhcPKFQluLiNz9
QFIkeAzBuatWDFAQwZHzf0aZrpn5STEPKztp+yf/WkeFgkqcijUqTLvvd2mS
zh3MuqTO2g3KHlSPWIlZr/9cOszhoU3aO273FgiLSx+ckdNArzQdrUAK/cN3
uCr1QbDKSdx0EATOtI+idG1TDvCI+8sagL5iRlN5Qk/azcfwIzE4/v8+PM+1
cWiN54Okri5d/gCbBBivenM3Lj7fQlT7y1zfuZR0b5GcwDAuGGFRJ0wJPh4t
Hyfv701lV/mpa+PJlSbsm3fwezsa5fpjc1nY8JDiGYs0Y/p5Twh8jc7SjG1i
yDRTBhTk0QYWQ89PMu0UsXt3Fzt4Ieg8Bcu1vpe0gMGCORgRm4N+L0Q8EvnR
pkZWc9ac9sOLZhiBar/agANGrFCFjWDsgRxPjHIndxqyUt9VK82dtzmf+rHV
nHnKNqYTXT0hgd07ofu95POSub4XRNuJGsN736zdlSBIykyqr+e+htPk+VwF
vfxTHQv6eGCFSTceGc22Gn323S3mZJBs0kywBHjTktmvSQm2c/+RjO8kQZyN
KQmKwIbk6X5eH4Z6ICttbpc9OMnyXNgGSmt5xCSBshbJXvi8KeRzR0QnIH46
GHu3wymwGpmhblkz5mN6EJ+PLo8LOEefgqpxBbbP8g7lNACGKb+QgE3hX1y+
7vy/0A0ICfP0ciSNhB4+ycMrt/4mh4YT5i3kTurnxHag4AI5X/wGN55aYg1/
x9xOcmYzd3J2ejUG9AowuJ6AGprZo24KP05kN7mhnud7gDz5QEZ4JKDZsOCQ
n7qzzH/hBN7wAHnGQRQIj/gfpwb+CAS99cXDJKqCvM3bTtEm/0Yt3I0/nqg/
qx3OC9/G7yJdlQ+s9fN6ZRZD/uKx6fMS7as2DhEcj5UbS2ShsbcHp7dLahJu
bvUJgEA65Mz4UA7Y9R5p4QqxtLbcJardyuDTNpg0Ln8FmiOtCxXiCbgGrBkY
NyJ6T2UrPeI7a38BRgFe1dIU8k0YgIYgGpOVufJ6TrMdjsIUoJBCs0o7wXST
o/PTge2aosFbJAhEa4AqhJnPcD7Uh8OP6Mam9hqKnEgeCRGEIz9eutJ6eq8x
RDB5FzA8f/poXY6RqGgEYEsfoLqqyWvfWv1nndnPl9p01+wGhV8/G7r4mhBM
NRbnXlcAmybY33TCoVR9xc6d0bGCK+wGPxNMw2eaJ3o0kotw8z5oFejnkvsT
vzttJ7tGEo57jV7YYLA4+gH/jWUKilKI3dT8CpEnEC7LgEZ8/6hPbhH3DmTe
YzJN9qvhAtsYVJvaicKtyLwbniWaj9TX2C+6VCK1/kI0uQ/7bz6BVa7SM+gX
uVSIec6SbzFJHgH3cGgsp8Q2Vi7JPJxHnb8z/Yy9JUgGqLz1RvdW97zFYbmd
8zXciWummTcmCvwaIz96TT9WdSE892/rqMC4oqAeO0R4TmnRHsAhIIab4/N5
A+Uy107Ad+LGVlaTUXpUAPoaaj2S1875UvqWYJlgMAHoDdGhmcIwb/1mAi+c
4vnyvEiZ3FXqzZxbSh3hBPsG3LGTzhZpqTefwelohQBqD77C6pIZToSfG0kP
XZCWkGeTo8bhu35kSyaOa2NHOf/ybQW2KdF083fiKxoNWt4tWq7nTMm1MqRO
Z8TNmwEZ4GWIZQ4RdUVTZECyHjSDMaKfYh8T0NkPcZOBLyHiL0eVIVGtxIYN
jZhQX2ItCFQwcYKN0sdSzYNEVDDVkDURnJGst7VYMMbZ4iLYVMFNkFHFJkdf
auDYlx4YRll4hJOp6fgkHujGZtFiLaiu537JqARByVRV6DYpfZzi6X3mQnSu
vl5AljtpkR626JCRqfsluO3fUbPOnOUflmbOonrc6H8OOz/07idaMraaSlc+
B6j6EHhKYfQJFf0kG6QfD681g9WQ5WwpCrqNTRo3EovqQFKhLwHi3dUvR6dq
8Oi60AI+tUOpBh9wsvBOhq2X1X9pKJnsttgOwx/jQDIxv/WG4HF7hm5LoTqK
31Bjyi4T60sHje3El484DaXt9n9lHPzmxt59trwWP1G0HW8z41MWue0Tuzkz
fWR5VN2lQLhdJeGyqszRJNcBeGLugmdecKAtkIEJ9v2sQ7DU5V2Vx37S0qhq
PGwEeHjcEQnUz5FlGDQZz/JjGWJiSmQtS/vNBxhZprtgqfq7V4lKHcvOcYZC
7KCgDYAkt/2UjeHQrx8FO1/ZueuRQeQq3/glvzJ3AWyrOVIN2S7n2lht5vz/
NUEJP9+b5as+Y13KyidObujO2l3wyqKSSbwVEe3gq8WsW9tX+nIuu0Iu6xmj
waSU6hHPMYgzDcs90OJDkXBGW0MG9NhPhkvR9u3p/QKR4OMuh4A91s6AKKMQ
auDo+mnJWVwU8hY5akcHYo4IsgEWhyDFdVhrsXURlPR7GBb9W+dFR56Dce+P
J1pA2tYoKHEErcXxmGpKwypuaEGWxNKnYeLNLBL+vAZm9gvQERZoQ18HuKDk
lKyDR+7LprQ71D1Hx4xe8B7UzXypYEbNwo0va/GEZQAZ3bOZR10oTV3qfvzG
6406WpqNoDI728iXB/rdUFaHXUJmAHd+FLtNXm1AJEd+LkQkZMBjTYP9zG9l
w0oKEiMq1RUS8E5iUo3gsc5G2hxb/FqZv4r3ooeXMrzHIt7Jn0ON1EJDNiHm
lF9PYrpqy/T2N5qkmP4YQSKQUs+0hF+epmPJae76vRtt59dAO/CTqDJn9okj
y8bOJSye4voD8U6N+bPaAZ8pn9Htnm5le5tGV33QYV6jlWpsnHeJocFqibUM
P4uPMKqLyB70MqH6xTAVHuVYOQ4rLwKFh1gmPVPCXjuhSnMzWW0e3PCegNr0
Q9FItvcBB/yVP2zQ3gYwJ+XVTDTtCdiw+1XA2jcuG8WVLMGZ+WJZ53me7C9q
Nju4GKQ6TvF6fqMY60mqiYeVuUyp2a01IIiRssdBbCD+0XqbaHahrrVYn7cf
U+aS/eyZJp5vEsyfYsaksi7wHTHoQoxXp1BuIcq6nNZkvPb48TbbCprGKHc+
xoKuV6pgCdSjE7Cia6OqGsmUlL6R09XHlzvPIb3X6skAyEGIadIs5Wv0yIWX
8CPWZR228QpnbTnDzFagwUyNJEhkdBaLwdany/wpbfYLHF5tm6YRsA23Dqov
DDxibotqohIOdoLeUkAt3duoNxIJsL2GTV70lmmJ7BQ98xAM6ZpK5wYUuZ8m
o/xqkEAznrUyiyEkqTI306KKDrifv+mSUhupK2QiIsH1UDaq8Z1pD9Zp/fuT
c5nf+PWtcBv6QtV5RSj/gTmNfbFOJQurNZdyYPqX4dqkpTasE34tlwKRrMDm
a0IjeXqDa+5bP+8CWR5e9QeN4Ne+s1n+rg2okiMWQ4J8hiyN/KcJ0XMtbjmj
UWYA1njwUye0VGnnxTCmGEdoORtnU5NNlYiwlFnLqNLIdEwOeDynNlAcywew
mcl0GndcDRrxuWWG58DKvCpNMBSNo9/FqSpXmGlRzgZUjd6Bc/EMa+c6jWSs
Aoe8tDEVFp6KwSqKytdFoPFvgsayKNt5ejhlnwDgVhkAYH/pKErmJGusuSaS
VqB5iy6NzVxkbugYp0CUt7X2Y1THkzfkuJMHhs/BRJeebh8Sw5CVus5rc13x
JsyVFbCwntgL9KCPopY2LGmNltKtSyj+dRXq6zZwMN3mPc3sHyQtFI6QpcMV
g83jvJPrZXkf2TcRAU+wsl5cRDYPlTCMa+JqMllKjWeBMNn6cnsXEzzjphRo
3FN+qvAmPdFZyz8FiiIhxY0GlPzU0tLMZ+8dOY42yF/W89gA3uuGjgw78Q/R
iOf/Ru8IXOQbw8YVq4ZXWEf4o+pa+migxrH2zOtiB9V8ywomUXVdaO9/4MUO
cqw0MBeCuOcmJnxtQ7Tkxe++8S3fYdFSJFQOLFTJJjL30lFICxsoJhb+xoUq
yATsuY+wXVr2/YgIJXhThDtI7Kmah7fijSf/PMrN9VzQpg8SbpaOJn5hS2fx
aGgPz/BlptsA9IT3eEBsrML0FMrQk2rmnOtbKHlmIcFMKVZWJWO/1/aNCdJK
ar9eh+Crp81XblVLxpb+2b7hLBPeDEyjI1UZ/3w7bW2mruTRkblOOfIMa7YZ
Blwr0EzSr8OZfjSGpaDEw9Xc+5TYd2Umh1AXW28iRwLZq2lfkVPVhCx/ZYsO
pZXk/T4EnkflK7Dc35p4gHsEUAYg07PHVH8hzUJKMF67HqcGar+71JPn8sXJ
O4QkEDu3YFasHtss80GMIfC8k64EI4w8D0MSvcS3V/+G3HWAMbglLuIK1cyk
+BbNiruurKLB5jlUzENJf7idzkhPl+gnS1JIgC8jn3u4BpqYhhX7Qe9TJoZu
CXvVCLMXNmuUuIKf0RJcvaNGORCOyzWOZUow47YFVWMz90c9aEBMEWewnhpw
hH+F4mp7tWpT6GTP4WIviZP+Vr3GWC8Kfd/5YTodOpy22Arrk/TPsV5Hm8Qe
jCg1rXJ8v4lV1U5z1GxfGRSRVuVRN52RT3jzE45J4zCGNM1a9nhdu25W+cF3
ahrRWnOaxHfCg7L1HdAhHg5lEf0ulwd5s/S9HIa+gNKOm9e7/ua06kNVQUqk
0uygW3twPVsmzu4QYbiAQ05nReY9V6vPaLEi4DfThQnSaSU7hW4bEB288jcS
n+2UjXA2jL2VHrjoNbvKwYWMUZmc4v8tdp6v3/ZYCniTuNBh1Hs4Uuqu2Ikm
xOWtKwozX6JsXjg5vGGyTXBP7KEpyE1gq32vVijptiRYdYbMXuKtud5NHayg
QXm9t0EG1OgsrLS9Fo1rGbl+Ia/JUPDqjkbAGe4YaEEnDX/kilYQ1O5/u3rw
sBp4f07KiUXwY7lMC8T4h55TQ+r9X6MSyrr9/7/ceFNl35MZOfsYRrFS0kJ0
OV4zxiAn4DfLANzyN3mqcl6j/KI03DyQWxj3bYCvM9xLwQ1vr8IK1yFNzlXP
fDGflrVquc890GvosFn/wobbao8jeHbTIVovP4pLSfuyK9muAfXRCb16ZLrQ
4nQnBBqbo6yhtx81NdSiMKqoK4bimyZpQtGK/USexhzQf8rGj7URuPDrN3oO
YB1R485ljihlMzamzaxfND3yC5ggaEFOoPfXRwGSWv4AdKcOgacYuTXgLEDr
R/0nRPczlHFm9TOYuo9tE7eykvWSr6FUHjZNUOJzdrXB3vU5TGONsUBmQdcq
LRbvLn76sYc70CRqHbQDb7Eu5u3JgBI1gWj+a1etrSZQWQrnZZ1YziMSLLMX
isUddHv4zMj2gasT9+MNugspmNf2X8efY416AmYR2VeHWcmxBzyBCUz8rBBO
8Ub2EIEfMJIpYf1gXTCiSm+gAY1/iP62regIVk/Lh2F5W2hNGAIZd25zu/9a
0+rnWIgPwIjDeLvRAPlLqEadD+F+dATYY4M8B1JNbzeAIiFp6DrB4pWF12nv
kJ7NiyU3w+2V+8E7e/Bdc0rxKK8O0NqVeoCWHL8lMaCSzjIJJIk5jAjNm9vU
CGRqtoyc4/OzWhMlE0vlpYU3WWzvMKT3SAw8UiMz

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3E/nlnEvXwTOnOKCtMjVX2BagCc0Tz+4jHRdI4rGDYXsh6VbHOl+XX5pt4GR1IXlgHzAzMwTId9LYL/5cxrVdbYDHpz4Llb2yTR+JIVNSLH0An0WvrE55r0vWQZoo5V47qWszHCJVn+/a5Mui4cCGAW7dUp5Fabi9KJMMnSYAukeqm1vMkd8VGwR4wL3kVgKI6Sp0loII9sv0HPNpS40XcBm3oEWPj1QX+ASjLcY+9kSU9qCY2+x+/dZojiIhpKq07a4RNkZGLGiIdhoVHxM64pCrWEvGf79R9kHigg+/gglw7QyJNmXaRQxj3FXJSsBjffOd31xkyS7nilJhXkvn/KHjeJ+gi6PiM30iKKtfaK6dQdKQmpqns5KjjQaY9mO0dZKay9+3eWy6JPuwG5pTONdZ5Lqzhbs9fEbUQdO0T9IUdoh1eZjdZSc6ErX6tmwXQMyFMDZgyps9oRBGU6HC7BIwqdE1mDww1KYQxerBf/1z4Lvay4VOjTSpq1PG8yPXaqAdZ3b42lyJny6OyuGvk+KRXEKwrHK9mactMn/g1O59DsLfh0AsTpwxhNFuuglgaGOH7QkO8nbmF7hK9HzxbMr9p5MRHy+fvSVu8MYmoqEJcj2xzqkU0dy5AKq/U4G39VIGJ5uztP+F98eIoriPqcaHYy3A5OZ+Rd5EMkJPOBeDt013XOsuEIWbh2buvv+0n6bT8TJ/zxnP/2iT+4a09rLQhYcWNLNlgnb+Xne9ZYKUcfx+rFTkCkZUkfOU14qIW3PV2gkW8ELEQAn+mdUVab"
`endif