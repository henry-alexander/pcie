// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
Gl1UwwqRLWNmEHW4gZrPbpbvC78W+iGbmQYeXoDuFuPkQTHYXqAnj0llcFiS
afVki1ugvVbLyalGjK6b18gVYBYxi2fHUh7XK6kkEfPNwoRZkrFTAfOZk/O/
U3u+mmCV2ycqyqN6n6EJzCZxcVzk6dRpDyH2rC3RZITwE3tEwX5o6tQaIpin
8mCCUXvcFZ5Tc8Yl/mEGIreMt3fQZGOZ1PBUo4nGCglDYmIcW6Ixb4yLtoGR
voE6GjWO64chsPk+n2a+1I0R/+pA76Pj6i8DuN/C2JLyxVtimi7DKuQ7Wwfk
Z7VJXJp0SOtYMExjSWc/kYN2NH+CiCl64n0KldVSkQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
IQnlD7b8d55sMJuodhr/9Wh/wD3ZbIjaZQPCn5R6AHoIeRbuB3Zfvml40zo1
n+iwCspSK46cDrm+v4BF/1kHAwAhWmt4CkhW9CXrZmSsu3t+zqGlbc/qwVgu
OgDCSCvAuSasSpLBha2wOnxnrxI7YbkF40fxO+oKXb8P61j0btrU4+yBL6DW
/8NLqZkjfuKVkjTIxqxQttptIz6NG/J5zma+V8zU8mwOzK1QJ8hBiyeNEPJ3
qZevUYfcXlg8g9JTBToCNmXKB2qi14mHluhwqA7UEqmGUZtwf7qMIr/R9nSm
qkibVf707GShsWpKr878C5RL19BrT3/QAXCnrR8Agg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E7aKybBDgj6jeIDzSMFFApWDpxmDsb0ro/VSPk4pAI6pCkh4TXx1Y1D8pi56
yyFdbaHMFyaCG2B6uZj74HS9GyCbLb6UZdq5QAWc8r3Toy7VvIrSW/ytNJf3
N04PyairlC3rrJ3LAf4BnsLXaRUZqLFslJapXbNjLxm8k3VxBdtXNtft3AK4
bR3hQRrKEfBhTI/NptLH71OrlfwVDqDENpGH6EbeY938p3fn3H1OhcFsWQNp
u4V6TlTtyICKVclJcsWitT8/V6lKbKKJJ+aujVnhxIoTqdPaBeoe6Q+Fe3fy
kCkYFLsecUCSqRkPqOUiqqzmEkBD50egcEMn8XsYAQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
je3DYS2Jsk7/JqqRt847Nj6z09lNmWl5H+8IPBhU2WE2OD1ALIKekdsi7arV
NLDY0mRRfmbjHSF3LktdLk9+FMnd6kCa3IAFAhMcy4s/6BsY5yrzQDN/8gqo
PXSFhydgz+Sjdyu1Or/kjQZZPbNYM396SkiZxo9hXXM4+RQ5qkc=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Z6GD1MGkhXCXCdmkB55hEa9MTE4FzilnK3kf99sNxA8CyzkvfcZVplfiYJIH
2/4L6wZ1g45+moowzAOmspofQ7W2eRshgB8pIwSm7Cyc9uG7Xg5imM0Wq27p
pl6FJN2H/Ee/CVhVoso7RxPyrnWHKmuCjgcY9Gz6s7YrDords3Mig2D25tIv
5rYvz8lR4/01tdbVYvw0tzS0ryKDTpZyVvIQ1uXNrZ0x2LBNkVkBkfHmlk/7
1sgBBR8AGvBZlxTfBubmbiO51fIfFqoH9s/pgdKNtMw3wM/rrwsmz1qqboqr
CiZJAmizeXFcsUVTaJKWMJaP7EEjTEeziqS2ooZECFebq+KfAPLNzVaSEpCN
ZnhG3H/0fzMMQM/WI9gR11rnuYLEmysy8/TP1Oj5eqLUNeuKMylCM00dW0tX
YObjHLziODN3TmXA18AZZmPhnzqOCnyDIcXe7gUd2oVjE5f8Wvhu+Z1341vB
1VF6NbEE8EaFCITJwM3i+RVx8k7sMG94


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
I5s6QKYnwLVFL7SPaPpt7gD0artVWbfLySkcadAQ0D0qMkznOWaL/7GE4oLi
3mtb3aFvTNUPrBkMlWP1HHidKYJxAZ9etqiVuFNXdHbqMXpDCeeBgWEfd/oB
3+uot74QECjxSSaCO6FdoaWNBZvqBGUDo9YRl1sZRz0oKTLjzcU=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
eG6Hr21erkol7+bGEl7sDTZp4fE9mVN61+EvgyyvJHrk4zGQpWzeEOSigM/c
l5IAzG8ACyRdsXHp142C/ZcuTsZdjaoAPpWhnWGgR8wG5R7E6p/l0VSrct5J
i25v9n5fBuj3JEai/WOSX85CuDESB0QTIy8H1ewIb9pJa/+0ddY=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 22880)
`pragma protect data_block
VbRvNkoe+Ma4eKUiLNqvmXoac0szqm1b3QCTU2DLIYE0rWIxByU8Vn0+BpGu
3Wi+nafn1Eh7Zct54Jrltry9i4IXURm757bttJba+OWM5fxkgd1y2ILj5buS
Y8lqx9gXbE6uzjXOr67Cx9ktTYztGvk7gXD1eqPvNBXz9heoHmBZXOh7ICUm
VOR+ME4WxOV4FyHDX0SrG7iJkdQDajqlbbVQlXiMI68Umqfx7NrrDJ7cHWeF
t2JIHE2anUDRlScpnmRWw9GhtFRmsdK4OiZh5tAyWy4C+DhqMemJ/isz5gcS
EfZTCSyCqCxcO24e8iP7LmReBYAt2yaOSg/pqbM98NksKJyOKuBdTI0PcQR4
g8NJluLqjNbWGXWxGxkB6zjyncGNic276kxQSQcNSZ1Cw3ajWEDnShKV139W
3UTleZDF06KEqix+Cvbx/SQ+E0ELNPBTFUCpBEf3d/0Yv5pjwFEIyglrWkb/
YodoL88tEgnMBJXOsyAADGQdWbo+e0OHEFe8UFJF1dgI1vqaQT2pHz7cWMXa
ndo9V4Rpo361AbNIa1dyUkHhpVdyiSvuprr4Q1UwG2VbLtb80FuMtw7V5F5i
pDiKCEO9s5Y6s/i2mO88NpmvRft2gxrNP9BKLyox9N5PhMcmaDldqyjExzjG
99qZlLe3GkRJ8wuIDezz1oiWHCBe7kCp58HICClH3EN6lajCZxZaIeW1Lvk/
px/qBRZehpNXcaJ5+edjYXcMn0ReEnbxz+O6cCwfizdz1UmLlfxqEXqjPBwg
sqsBFnqgRjyV5vZ9U2IOq79n8Lf+Cjqas+9ratk+h0UWXj6SJi9mVwbtQmNj
H5agpwLWVfZkhKUO4G/u5YxcMNXAA4X83d+lmlc8zJwkQpct5KE2Wh11NSrq
jCR9G5wscsK6+jxj1YDD1daG2hJ7/RGa0dOamvl1M/dSoL968v7b/n0cUhbu
TResZq2/bz+0g+615fY5muaAWx1HdlaXou0Ttv/orDO/Sx/uHRATw1imqZh/
44d2rl1vWRYFxtRac1LLDSWY6fCQROHFgKp/8o9/DkyvKVvqPQTXpnYFo9VT
gti93St+zCVUziobEb2uEYOQz8HLNuTdsljXgJqJOWYXmnScTM3iM52Pt9sJ
Nl/CflBVMSISrDshtcxoMqWdy8GR6vLVj6s3PBT+MrC9/4M5b8iacyWFnBw0
sGOIs2GhEWJqBNFp7M6vbCnTFnjhYVJmIjBm/7PASOuGQMfovz2II57DGh/c
nXsvO7DE3vIi5dV9/Sa4coc4jhYrMj6PWjvct9ae4hcf2Z2hl7m5LE2EQ48C
zu5agkU96Tdxw0Ss0qs2A/x6DHyYjcDvp+68lYXyI0PYJmlrrHwquERq37c4
eM21qwdOMzsEJ/Mfc6sMmwrceDvSpZgniF/YuraGtWjNFPg5zRU2XxyTnWx8
ooDYKduyJP9rpBE/WVR2qsZlVTNJz2qH2N5Bt0fIiD+lbLN2QbDSiVkiZ9oX
ET4XzUoiM6Ue3FXzOSSvPVwFtypAFrAyYTBtyRVJL8jhF8s4K42sajq4OuL0
FHEXTBFa7tkLMExcsyel7tK2QN14PnmVe0oWEpbRqwUyJDax+p3EOcm4dbDm
yBY+rZqmCNov98pHLRaPkDErpy5bmPYD7nLCAE2w+XHBLEsa3p5dtE+wQ4w2
Te8gEV+z1+4LZUG+19uB5SRBB7xFK/rJmUx6rYV91teczK7psZafGY8abSGy
s0SIwjRjj9FxRvpOGjc+memPZWgJ+ACD3s3p1S5LoBhfSFMrU8rj8RsOIl8+
cTfzINRJsgdxX18MDibpwywkx7bwJPZmPn4+Wx/J8N3lZ38bXbDStNp50rLy
m9l6fipcjzOhEQouQAptXvOOanSKWC/ryXwN6KDmsxrQgQ/l5+rLY9v/De+N
41rG7O+guZ2NPj6qYnFgndFzgOARqRj/5A3GmOylCQ6lXHqBH5F0FTfPgd+W
UPXpEXVDqzyzbkg98N4/IurbE2yKTeIDFA5j6iVTRnfubH2PZIACcITpeFYa
DyPFDPRn1TOLnQOQahPEMy3NRLQrHrvxFbq6IfxwTID/ndpNP0vMiB3nMOkc
iw/ghtGmi4wjVmwxN3x+q3PK9cu9A4cz/GyvdRoOLs8l3fo3EwYs3wEBVpMB
tFOKtTiUCDCbdiAn+X4rYHlDvfyFFFnPhHpSDz60sNbY67R+JEH4gE9KEQiM
5R4Cyc4U3g2UbcKSeIC/kOJBh3SC6pxOE3ODnf/exgEph/PTHIOT3bmEvItW
1PUwM+OwlSPQd4O94/scbVP2ly6O02j6uN5uM8I3J20e6mZS1rbZIcgaTR9y
ebfdhmmIovNwIzLmULYm1nfXc47nREHe6TdXUc1pWAaNTgiDBSnVp/1ZPRNA
r4Vb1MSbQTjpUfAmsvEfYA0EN0mbiRntgnmCkNbu4yrjMD7jCv8x8NfbQGEU
eaLfPkAFFFBmx2ALHMGBs8yF9Ubw5FFiG/MQfIvSlYbDiplkRug7pOEEbFto
50sRbPaZKfKDYQPizoN7VP58j/R2JH+LoCaLGOAltTDRtOJqZzl0JN1QGiFR
4XYve5Zc8Ry7TwXplTM84IkcrrAB6tCEuB1U/EICoPqSu4xGW/qfeku1TBR1
TqdryUQnOTUA0m/4q2Q6snDJ5CdT7Y/HD+p+soZpUQivtihplmzLEZCDoZcj
6yPWBbAvyZmu4RhnqlHeNhDYdyZI5NU1/nThTRNZ0qPsC8aqAs8NjDOWc4o+
Eok2AAT4hdpak2Sww+Kz2SZkTs0G5+305SLVk+0QIn/zEZJ9rXXBqR5UZAjo
TAilvGjxxYrfmFkGeTMB0KROrIpSYTSe0Fw0E5fRh8LDeZ/4uYGQZwvgrCHd
CmAnUEuOb4J+bsMh0+xcG7fkRwFR7DraVN+ns1shxeiYFdmxvguloQO4lkSN
+cmLlsrSCO3FbLNzRVQZ2MbVzAVcYFkqxJDU9Ysj28SDjz+JyRHJOvLRyHwH
kPUNv5paQ7OWHhDCXS6uXyto7xuVUYuCRlkpf3yRXvmldyNTglUlEopbgneR
hn+p4VIvWVenCIz21BHYZS+deLG7CNnKmXXeaT1NzWjCEQ4Z5Nni7O2mzWQU
ZnG39xJ07+9ynrihWNISY2uIyK54q84IVohm6Xjg6kItFYnnIh9uyfykm7q2
lQE3cYvPwK4PgPWsWKCS46HP/lgNNMXCXMaH//HIOyrgf/WtFZEDlSjJZPbW
g28yhzJvZQMcBkzYXzl+exLi43B14KlWR84c8B/KvI5/cgCHGSEvow3cYQLP
aLU+GUCYQIwdWle3dRL7408tozl/eLbsjkatBWyOm1EjUr9qB96ngpaesy3C
B1v936QwAwNam7Q/ruvHyETVQy4sYy/5CRp7x9pdmMBZbbCErypAuWbRvKEp
rj3iF21HKfA/+liV+b0kaWhzGzb6zU5QEawGI9v0FotZiYoo0FBhUrggk4W3
L8mWHClgD2Gygv1CUcHoAPp3YukEosElaCaO96J4H4tNE7u9cX2u1jXqZZFP
XE4YMLjrjCB6xE/mbbWdQfGD/ZOu9h7zzAHr/cDURVDoa6I4M93/KAXhthlS
p0RUumZhBSpbjzoMc+4jCtwBT4OcTFrkOD9IzcNnHpbLTUg9/hhLuENGmQNJ
jeieNoPRO6lk5J3xrALYy1FuAgnm6gPCf1VpS7aPIR842Ieyx619WmmJd6+g
9DpOeyyR3pQrQyXrN60QzRnAovV2EJWSY6jU8U4gzUSRFIyDdIM1isD+AMk3
R7nd4uqJvJqN8FU/1/zhRVW88S3EIVA2uk6nWWvg+4OY2W5SCTslQOrvqcYH
BxqF3fOXMUJlMc4LT24ZA1BDcNWzg8VKMzcJ/W3uVT0IW4ud2Ut3GVVIsVjX
vqdh0SMNRLoUmTehFcvyzsVeTLmQSyDIlcLZVxzmo4493pKsld/iQiDPe9xH
Ij1rGkBwoWOvpZVHSpl3U1mREpHfD3EVtSS5pHuDG3Ma/qFFVt9+NrLeLsSF
VtNPc82OpiVfJgrTIas5c3FTRbpZLlKOiEosWxd4hMzji3yxvIFv8gPBfdXB
SNMlueXi8p/lwqY4TaGBPjL65657YRvQ3npe8laNWeeu8OLlEO1SyP0k/NdQ
vcIklk6CyhuY5hm7kHK6iB9qubZYUJa6t+EzTjAf17KYx7XTu0pAfgtSuP3n
OKFMP3++8tBHsfJkoe6rxEBJCsZDkLQgazzZRZR0y+JKC9JyRhzH2qN9UlOL
fuPGwf+CDFYKOvd8WHEE/iLx44eL/uq8UMIB39n0H0YZ5iBl3MDOIfqEHGrT
IdPeif7E3oG3DTroWD2y0rxrSgjjdu1IpdK9gAjbwdTnbl2oV+EMJs1XrDb8
KE4dCcf+kQhoz03+/eOA/QxareTpKuBn/s3tdrjp/zrrYLpj8yv236CdesTd
lqUZ/lkqhvycpKbfvAM+2Gf3swdEBFfDS6FWRNzDxS8FcvdG87K+gkCfqxWt
/jnzhiCZD4Vy6owhRpE872JeLfGt5e3zRL0Ayyr7q9nmyaMEX2vE9ypUkSpI
TD0NcW5gGGKjrfeJ7ammfoBM8VvsYcAN+jt25kyUVQohs5o/fP85q5SSedvk
LOxgJG4AlAa1ixih3CE8jdUV/jtS6D358gI/AXodAfWEqG6GkttGlk+t3TpV
lYIgQje2r1h6RjNQkxaOGGt5vRGK3wjumQ/fa08QUv2O3OVi5PsZq+p/YKwo
cAB0iv8w7o347KUL+i44PvkXbbdb8v0dVfBYDt3zvhmscD+gwO2dUWFSAp0z
HdbT4081eWmBXdKLDoEREUg1U3q57BKaueZdEL6XRQHMj2d5xB475ASQ+SCT
YAiFRJImDnk/6Oczgjby6Z7LEK6WdZX9TLUcz8ymV0FQjYO7wZrHc5hklxfn
EkXFzv7fdHkS2QY20/6HwcLKVIS/u+fXaM0ZLA0lX2YqqsonRZhSRmwrDoU7
42qMjvoiwdRnW+vEiUIFd6jjzzND0MwKNKaoMzoamDV90fm6t3bIfihjVC6v
mxMGSV3hQJcEOtXfuTbJtpjiHz+ylfOjFBnRkqX8vdqCtV9iWIZUisAGvIkN
0AOfeej6Hr1Ff5jWCtLkM9c0dkSO/+uenyaIWWzBigwjr+8KV4I3Cr2BcVGK
yDZbpB8y3n3ppIgbmE9AXLI5x8QwOEvHdviPSwlDoSkrZPiX1PoCuQuPrCIH
U7KcB//Se80tYb09bBPSYzZ3OZXco3cHUQJqO9GPU+BO1LrKe4mSnKK2RdYJ
mmo7bt74KKZTyV/ymep1HIt27Ihj1cFPVCJXGjquDa1R0GLjDOqGM40wyvis
3HV3+qg5VSbaZoVmV0dOEWBBoR6h1cOBJ2uOgWBxK9MqopUV6EobVUtEXh3v
UVBCTtH7hk+4hLk3hudYRAhDZODvYX8LqFgpeig+Egrtv6L21gq2KrNOij8p
He79nIQhgGDRY/RRIBINVXmhsaltamUMenC94LQDObz7jRrZ+tQaBVIUOGe4
R0/XJmb1wP/EYIOHl9OogfqW+PLTOo3+H6SY5Jqt7AaWtdUOitMcgFapHIF1
MPSWfxhsuiot6iiaXE5dRwYvSoFogbHYbZl6zGvLZvy2QYvzPqWYONMVkQIH
Mp3RuO0B3Xgxq+H25rC831cSuvjtARCYR3iGQnolJoo0ij+3vQMUdzPP4cQk
CvE3TRtdLdj1xOMTmih617ENYdQSdB4fG8Xtab2lYXuOEPq9zd5kQnXftPIZ
2bpRCUNKLIAW4IGszFJ8B0M9/8oumLkbgNGh3XLVao3qZlbM0K0SPPqOI85q
gQWgDnxEVC8KoVfCN5dilNK+xoh/j9M8zW5Au1ND10b44YZZh1BqNOhCGCAt
iutm3y6PDAHkawk2BPNTrCQk0NL5BpRiAPAKX2CguMMIwyFy36rKSPlbeCfC
0SeckQqXqDfYK7HQkYqocgP7XJUE+CL2ikZx1wKQiydc5VTGk11p/Db+88Gr
RHehLnh+oWtazIOKVHdnIkD5bGCSuuJAy5NmUgj1FpLHnSnJRELxuwgc0WTK
tSaX3qavOOXsGK6uw3jYkIkW5tAc0aAvSgDG+uvJVtI4yIPwSRgMJnJbA9Z5
bwfVLsTKX5ExmhkDA/NbKi727vFEuP/GCymjiMpvEXkE3hvgQ1XgZaro1GuI
BE3k5abXE4IOqb8uCeHWRwmcVgnzvET2QncbkvMqZbWM8yimspaPKbPI9fR7
cJ61ZN+/eQQIZ95aD7ic/t48L0Qh8UkmaUVigd6Mnm6YJNC0DuFC486oB/5l
rQY8YsSR4cMFx9ilG8Su544lUskZtMrecw9EOrFwxoIlzYmBbuJRprNQ+dre
HQ3BzPV49W2MhjFhRHNhgn0x9lT72YRyqcpA80lMQROxGtY9x/9fpC002fSW
4nFNDEbabDech1Wi5Ts19VSJeZljY+OwKZ25VrO0qGeocU7JlyFGcdPdGfUv
3AaKmVTQ2qqIdycEEmd9tG6h1cD8jlOyttfSts8XPFynCj3dW1o4UgWUe9DF
wcHOI6cR+oQGzbhb12HT4IUXiTlu+MQlcXau590JuTvkMMRh7JjOL1nZEEuv
3ChSei1zvHhSIYReLe08oqCKCqEpo2F2GJpd8XpsZRLzV//V72ab+nZbSd5c
Jd+xbhiH79dEaO4uTjcEZhulx+AW0Q5Rt5Q/32BSuS6pVcBwQLT1Y7EkGCa+
WdAowzKBVtBLByd0zkR78kRi9ThoHOzs4wfeXhoI9sALkKkO+rXBJ/GVRqV3
d8E8Z4V+TRFg+vREugwM8qtPcep94lLQS9WrDK7n04WtfTals/zCS4BAsVTQ
7kgdSyuMpocU3qEzcgP5coQsdLjD+W356hXC34ieQOHQ6CdJKZnq7pE9npR5
kmpJPHNdS8UM2HoKKbi0m6EhkItndAoH1wFgQE7S8irv8ZGVvlTOmdIblCD5
n3Bab8Kwz8B539qIR0Adbr1Gc9IN5MfVFH64NqOiCyKJYBtjF4KrRDYnnOvR
i5imr6Q/X2T4Z8qQnL+l+mROUhb4KTtdQKp55gubTXRBw4kjdd472chpwv0X
x93Gh6UniN/UNzRbt8foE5qQx31M4ZmWeZcf9SUpMTNezmLkuQZ4dLhS7mgo
0OXdSqc9Aste5rQ32warXin4S6bmX5+2nzu4oc3zinCSe9y9FFkpOyXTRXXg
/6+Oc+DNGS1XEC0JuXF7onsHDrqf8RQZsU2NdVCclDTY1Z+nxWjl4W0C3cWC
f3eiH7Q0H8yK+qWhfnvIS1Mqu3bnx1A2WkHSb/il7ru616vnRqp08081s86T
eU6fmIPBJioCIHfrIYlieMKYs2vTS1Ui1arMYmn++eXCRPR9Oe1wD/In0wRl
CYFUoiafQimyELFBP0sqJ+b9Wnd96ePKmJMTxULWL52Q2OUs5UeUbcNQ1dXp
STZGDHwMFId+IQ85xgdYoWxlHWzbwW7kyPlt708cvElJtbubJ+bHmu0AA05x
u5WVV2jhDv3dN28ZtlG9msn192kF+WgyYfAByrdjPK8OYVvKBbf5NlTq4AeO
M5CEunaH+9khGf4vCDfHXQiifUNZUsv52B4O4F7+wAeOgAjm0kxuwE4LKk+C
jAXYn136SpawmBsmFyMSL8uoUE6X2Wg/2+WZeCRCnjwocgVABS3LCggIXLYn
UHhBFb96IAUs/EE11csvwJJdollV2+LGeqKXFhB2nlV5aqYIsOEjG3Vpjll+
WC5LvfKoCKTXM4b5t276Vy70W2ndlxna9liHacuPEWZgPXPenH+Cf2VxzfXB
Zm1H6LlxbjIkLCnlyrjQ4j0l6xtjjZ4gssYgLx3xRm8YhAuhjSoiOH3EndOk
RlhxpYkt7rPx2OVT+vhr0FP1YC6HISsm9iYTdWfAqKRA1Hg3tHYb66G2IzZk
1yTg/xS/xZee6lIJ7fQTm/c0uzY1LU/NpbF6SGjtp1R8ReJY+U7AIZlI1BHL
o+uhsw7mqCy0Ztyp2pAwRCr8Bg3OymNdul3ilksonWsMg6yt23oPA+9VpSho
zPPb/kxXJ66Y97C5atanzv1vgBIuLq05E2AKyBLQTsoyFDU75wiBPZuYHMRs
Mic8xVc+2mIPO2HciaZEi16ohJZWOLmo8qzfgB4WgcUSS0mrojVw1KylcP5u
zHJw8n6gYHBGPlXxofzuzPukC9J5LazRhWwIQD+HIYxZVk81PurXRgCNIQVt
lJGTg2xijB1AuYfWEp0ArR0AWM3cpo5diu1PjxhMLV8/zBuTmYH6kl7FdG3E
LLE+fOIMeYDXb6+YGUKLUnYhkf9UjTW1lINgsc4AzQlY5iBR/aR353kpy71K
jBIDfdaNtlc2hibzgXXXwKjaQvgly9clWOUO33bpGyC7Ufn8j9aOSgSBN6fW
URncb1gO/1/OsStvjTR5325OXMwBSn6sh87rTARQO57HLzjC+eEVskU1kKvM
7pwk7QRRrJ2daKX2TiukJvsNB536twGfMRcr2F9R86dY5LZ4860Dwi/KxjKl
gJGJiG3ycmnPX3L+eoEZ6KvDrjXuy1IKMdjF348YhdlS8tvlSdFYRDiPEzYq
XAd2lb5OKTbkBfOq+cMSThGTQ6WF7qFEzfQTmmZ3w1WG+k+T4TXuAz2GabyB
Okj/UePaOGfT1spFFtSL1fJUkl/i6Mxb6q7YriktR4OVSWHThxbcdUsU3hEL
Q1MzSnYJ58qqsX4m2Mw+kJ6EK0VnZiH3i4PAGX3w8t5LcZqy0FRa8sIk9SMW
aE4b7/5VIXx4JN68wNw2k05nm8evM41LlHuk4/xkqN+wbmGtvtm0gSTG10Sq
iYMLhIWiTP1sH3EV/2JAiMmO4SJRUeaIe4m1yY3eAGksAS4cSJGthXEJuvCw
54BaDzPhNSZQWopC7iuKlHsCjfMeTNpiZK0t6Dn0NnlmEmXIuHA+DiJYq8W/
NeKB/DKYXH4V0kQowulB1o5BJ/0XX8ym4w6kViDOn9kAegOBsMHKk6AF49Sf
EBGxbd6qWWkHgnqn3bXtUere864wIlzNjYtP1ver6z9tVbPac+jtPbe3dgMq
VevVJdW1hSE5XKIIrCBLQYpQtjUQGvVGSHxT+81c5V4DqejySrnF5MRofkbB
Y7ujQRTTrQ6F/XPWNEy332y9/gizduXuSKk5PWlp5GNwVQ9Ut+Oqd/P0Ovbb
NYG5nrF64jDM2u7VtU5lkJGKmJktFH7tkSy2MgWTUN+0QZCYxrGm0ddCjyUq
rqzG3lYgr8KLIcAkAigMKIY3ARj58Dd3MXst1kC18pNWAdtLNr7iz1s2nGwB
Ebr8RC3EIwOBwPtpbY+aBzSptj8zt/w4PCZ3OwsNU5PnaugPS5hNilapG2hN
HyLs+/AXuPEoPRQLs+p02hdGASt9A+/u4ACzzu2hANUpcrRp72mdtMGCwk7D
e+BwyRCT4PDNM0JYSuypZHs/HXogpAaOQ+CC4p9+AK/E9YRc2Ge+HW5j6R9j
r2R8wEJluSGMybDdZfSlKpQ+u8EBuTanqrbPrpUX2lQUchMlzUBhxnhEz8cZ
qkazTPNyukIgFqr9ncq6/SIt0RAkLwRwLeNlt+4vx7cBiF/Beg121ghXfz10
dmnDj5SLlHvpMNBTxUaMPr5Cf+jr0UcUc5lS+vC2h99IvHCf/9D73+0eeuTV
CzRrvKymMmJIVb2ujPSvA6MofUhgNi860CAbouZaiNVb87qTQgU81bO1mWnE
wsB+tcC3/O7kx1SAYBLNYAC3JyGV4sAV/DrVcDRyKg/u+FbhbETjKjIPQNzH
Mhns0saMCcHENEL7nZFddcorX6d9lScCcOywywTlFgfIMkCouSakx62pb9lC
SE1Vi8HDf6kImIOyS2aRXZHKOK8ALofVYI0v4/8NWJrwvHY4Kn36/iqh+QHU
X8097TnskDakJ8QIEt4rWq6WLxYD7H4qCqNBx+AqDWANotf1oan+BntNJZ2D
cKCHYpmYS1Nmzt30zbf26bEDAxLNOKazX92va/zw76RN+V8uGS/p8sngh7ts
g38dqftwoz4N+eluE2D8Sdy0JOKKc5JUrvJkx101zmjV6tAuaadDqPZ4kr4k
U9OHnxG3KNU970h5P/a7uPbNx1C0Vcl5P9muREs53EVOtBrw2ylg0+C7es3G
wNcQ+bIZYLg4YjW1pl+RVpHURYziArLDIbQs6Irz9xoVpcTNIyFVypMme7aR
soIezNQhCLD2X4p5dcxQQcN1mg7ZR4JO4K6EkJ5tCdLFmWae43l+kNa2dk51
29QX76P4ZhBUtzojafp/0Izydkq58dFo+S4SAQ7NbuYnn8KwkO8HmIe8r29v
qNnlEZMIwxOHkXu9AQS1kasx9jg0L2k2znwMyKMzId+7jyuf4WArfEqu4QU8
+27sKw2p8z+TcwUvWLAUPyhi64PbqEGDd/7Bjx4Vp3IHK4bMBKkipBGctBJA
5gZH9HvKvqPYAdZN2ZnehlD7DotTzhZ7O2ZCH0awHlb9sZZbVD/gqYLA03mJ
rAd5WM4qdepLqrbG8P7UdXL6a1pzRRel8z9SggpYjUWXwbUciQFn44cadNtO
S3jHK4/cbz5yo61QLoNdd6SBIO/ERGawbI9/Bp+DkZGsaMQ8n5TK9vmYz5jK
gR60i9ljhUzIdDg86pNtPJtDfAR79cATLqfSd6Q2Nt46+S44z8oIst3xWlsw
16bhLUsV6pkWNEXQF4DVS9L0eCptA+JgGPXOdYP5+HBtxaOjqbBAjjQhU1M5
VG4RXle9oA6OfOYGTBWBm1CtuG/W0wzhlOtu4ZNOBqrSrNYdXidEyVEMSDol
0nMVvavUl12S+UCWZ4T/Vfb1RycaLS3cI1b1GrTt9vyv5num+odAGcSlGseL
2qjEG5w3b9z6HovHCxxKrhW3BLNkuBjWO7+uRZxkFaEOdj9yyfb0oLKfTXzt
s5c4dKjzzG97XDqBxSoPup7R3tpj+azYUhFKU/jDU6rKwA27KB0JRYmfBqLK
updatrhI+nNxARubLvxx3yKwaD9XmYtfuWPRImPTZDDQQT33RWPvV5e5KARo
/LGsmpMYC1wYMOfwJpBYCTN6ZM0GsEKpqQG5f9osRDpuXGb0tEKbMZsfh9MN
IfUYCNGirsRv7o9ztBToArxYNc27UfZJ0tMw+XRhanE5m5BUua0th89k1aO/
SO0ZMnGFvDZv+3K4+djBDDFM99EqgQ4aeggA6YqQgi5VQwleri/kV+La758v
yDmE7gkGFwExY+YKbzOh1bg488jHasvGudBMVemwqOHC8PLcHBQih7e4tt/5
phZaH7AzxOC5rpllcLVzK3Pp3GPWnB2BAe3tO6ywERT6YB9oSAq5WeHjd7Ly
U9OxPt9Vzj6DK6Teqb/NPVuSyTAeFIcVULORrJP7dalRMUPgLoC9uRq2rsDW
HIEVd7/0diCliUTU9foOMNjvLHpIVoetuSHscmwkGIuDV+IAw6JsOMexn/qw
HdNhDeqh+XLV0+nrZE7ab1NseKpY3mahuYf5czpYx6BQ63x6cpoFWrRQWweh
xY5dfLZo2YEOqpjFn+T4+rMprKdXBsR1AVStWFpPK7Eqxd6iDmh/HgCUIBt3
aRpbrAK7PxKUqQyAVPMyDLQtniMuLD3ODfma/2QN1CfsQHeXvp3cMffcDY4p
TIK0HT7PuTE5wDMp9KlSWUBpCOEhW4tH9DyKrkk9+LwclKBpv6GJKbSLjTFM
2YlGBPBuDdd4Uh5lLTBFTHz733pQV0nMq3N+Wr7hXsnoOM5AJYF6SAQSCxy1
Qj3kJm2HbGf1Z3cqCARQOiFUDxA+q0GI53nZxF5pp0MohLvsn1fZbPOvk/gf
ad0wRS0szEnmGW6nkxJd6LNLWPQu6unpkzYsAY6sePfOXDXGDb5T7S2/kQ3C
JOGlnRjqBUXtzAfpTEt+AWu0Ye3bt2rCiKykwUZxcb5xS+lvvpgk5xRtqwq3
WZfR2lgojmE+LSruPFuDSmxX9ekbdJaMF0U83is9oPM1RGqIHUe7RGzQFioO
We9KfpQaKGkKOu1dNfYDbtHMI8W/7qdPn7p1OkDy8Ie2FKMklCeF+R4Djd7N
fjanWLLDej011/wSV0eEWBCbaKTDNycJOGBT7KeGc+cT65lhqawSqVPVQDPs
fgeo3f9q+7X2L45qqmmA04LwAAaUeFZ3IQdxWyz8bQqHm0g9lZHErPfJDXpX
U0oqVzfLYoQWAvgVTP2CCZN1eE7FlbDSczmKkmfTSkJapl+asO1eJGoQjaxO
ly3UgURwubruvR7v+sFZtK4AiTTcdmR9Bo5bRAFrr+GZQ6bn0a1ujuStwlx+
zVvOkaYURXZuCUvya9RTKjKZeNh+aJw5wE/QYvBrvQkyK1nEKrkHAqUlKM5k
SrfPT40JTmpdmx2PsgL1f9qad937G3HV6NgCOX7/s0VEzUsVF4gwDegCmrTJ
W5b/JxNofwGkvFOyLB44hE0jMmTOO+meCgnaLBdIcw1gIjwlOQ/Op2/SLP9V
nRpgBGLKKxS0watYi8KGoXjhDtqYX3xZBA3S0fm4Z5nOsYCmiRzCrxk03g8l
E6XhlAkLlGEWIzgg8qkBnYLisRyLxdXUHlbNLSgZ1uRL+9F4Ap28L/6xwzrf
ThcSXDXzyO2DH2yRc6pU95mGkxTh1sQauq4aj4wGbq5XlQ5NUbAHoHdKGA1d
yFS4fLCl7NikroQFHVDTcBD9mS8qc/uO6aoHWhij8TMBnrNTn6B2RP5XTTli
RIBvVlpWkvNvh8nc80B4OFFJTvANvWyC/M36guN4jQUVAylfoUsctw6x/iMV
btv4R6mhfTuEAz6MjhR6Q/RHhZOp2hZk0pe0bEWoZM3pxI9nLzc2b0jczict
V3ZFwXNI4zmtJgsvpy2fBELZnTHAwmJtShEU3M55+eedjHCoQ4vjAmjrZp1h
spyT8GL015uTWHKoOWiNdN/TJjNInPUKQ8j7j+5sKrIl/qCF3GJ87saMrwZy
2IYO53hYJABJ0l4b3KSMwi66eC+lTTOBzxlqtbDdvMQeGUnGMl45vqYIg/Es
GQGf84bX7dzfOctGQughTG01ZIQmlqYJSYpJRPcQombJJqyXQSyGB1OktY+9
T+8enR1s6FvMGPEBqFa5X5C4eA5GUWyOcIOgKyC4qNljP7BAC4RS6aE8wgfb
Qj9SqQK1+m4aWUMid0NRTez0TgbEZOp4JDCmUTNvrT6RGUvN2PwA4FRR7iMy
9bPhzk7l5ANduDh9zp8X/ZkraZxpesYPcX7+KNG5ZxLmnhkckGGucHEz7mve
h9tu5sd3901FDEE+sYCeGkr2ULICYCcAZalnB3OhLILr42Y+RyhJR7SLPOGv
KUSE7Skq+1eGh9RwgaL78kkc0uwxDIMviFh5ZuyEHbkrHvwhFmNDRJASo8Kf
wlPgjM7I2QK0N4p5a8Ewdtqi+wcdr1Pb0V7dFcASBNj8U3MdTnUkSvNWdGKK
xz2V8nDsHhI8hfVVoYSZ6lNwLuQD69uYq/yyKtLub3M66HH5AqDE4i8afhle
TXqbn+aYmnPCi3Rm2cO03D6BKaa3g1hZklxXlh91dqfMs0DKKTnwgS+4XD5+
0lQ3BkMErX1Te1Gp3CdBtU610zkfFAotPBc9WnFe7eC/OK1eWnzdKH+JqZLY
INEYSGeQPtbE2xffsojBeGSkxfkTtMBpm+iIonWTNSJPxp2JTFnjXgdJykOK
nJ70+gGVTSmTFbnc8Ttq4E5mdom39Kha9T0qmWaqQJJWcdoHdsPgc7mkyvJM
X4U1mnXwWOsVxxkx4nxJLdHrdd31S+oYUecaqGUTabLHZPs/G1pDF7oMq51E
G7PweofFgj6/sHrkgAbQwvXdQFonGLQjh2GB63u/z4p3HMk02DcDA8xNTIPj
KaLje+UcnZw6N7wpdF3PWyXrw9BWi+LI0NfmHafklnF9eojU4myzLtHEarVn
0IXfIkgO30jxRyTWChNlftRgJIXqgi4rqgztlS4wr9vFyM2JfqVkdH7pMQ8B
W56uY6Hr/ZFir69rsp/ZhN3T6BRLCHgNagmRgi69w/feben0x1bi+Q/03FaI
MyFQAS8taNwfJiIF/6CnIWsFzuL+T7DsdZRBTjBWnekp0Ls9L4gZ/DbfCH0a
cMVvFIESabsa6vnxa1sjkH7UYclxX63O4h0Vj/lQ9eHHHiILxXeb+VZVldGW
Q1tjorf2EJHerdawacQmDbAjRqnE4e02jkH94y0OBYp9X72bN7vuU7avq9fY
yb/xADsOnaHUSuEUTGEml9HyyIDzd4dTX9tbeG3SzaBtXAY8FCMS3yctiJP+
/PpSdx2882KlxGt1en7w1rKyZAXyHsyxEVuDLAY//ZfUWMjGDLFdXOsRqREH
nS/pMnq72jc+GO0V+/9XPbk4Mzt+qyhAj0fl54aESAwvbRaAEd3G+2wleNTE
4So41VLV0bFwpMbVROcR//QPuEIThTruCj2eUniQfrCQs5X2CrxzjUObVKsB
3usKb11bfcIXOlHGUFbtTX3aXtzoLwMvnPXBAHsWkWrsUyE4afFQSKm37Clt
5c2fMcZ/kPExXyBFTgXikIL9YK1L2JVENgl8F9bVvML+UJW65EK3e7R1bkzB
roDcFKx6ci86nOT18iMGBDfziIn12VCKl7t89rKlbuJ8XatyVa4/9QYAOZJT
ZtSaTl/PEzInISfRAx0T5s5dIWXVIG1AvhiiLnoT/8kuGuucDhXWT1YisIdn
vCh3MN1FhC69cz2DQ3jXbI+kKH/l0XiBMZyuaVHzxQMrFE21tf5ViUQ4BJQP
2xGCZKph8u+9yyfD3/qskkz/NoOkAqDHQnOEEzrKVq/bXo5PVzldH2xA36on
45u/dLgbHUhEsVK1kQOtRiRfj6kDmEts4ahtLbl3xR7OtMkIuj5saaO2uA6P
23DpEQrYYeTU5qLLrBCSBqM/xq36JQctdEEg8334aAFA1N9T3jpoxqtfH5HC
G9P/UloBoJXCvqAR8jgmlH2H4A/nMyyliAmkumgxap1eap2r/A0c5x3dajct
s2EeGML4MnhnHNm3kIRbR3vcTgzmPaQm3zhZmx9bdwqGBafU/sDJGH/jkm29
9EmLrmHqkInVnnM6WUWiwu7GJClyix63V7BztU9TLkmlh4WgtSaPjlOP3uU9
qk3zGlM7h3tw7Q/F15hb270E2oLKlhUgI0gxnfQK3ATsVju6DX1TMrclXoTe
cl3PxXxxtw7u7vxfvLaccLAENqyjEJ6/Jqvbo8Gzj0ivCFMZWBXa2m2Imtlm
94dr9yZPJ+OahVbsRCJPZ3AsPvTsI2t4VtV5PHfH/dEnxWdCZEKwrSYZG7KL
9bEbXMkmCSV04mQBErNwC8J7CeCU1+Vt/6OgZ4ytERmprdpq5xtbg+K9DuVg
dXZhdKaou8njeeHBhJnx/tl1QIj1NkuEDQpWh2dtCRPKUqfTaxmZOzx6BtUx
Opd7V+vRJdFz9fkAQ5fIluYS6jbiYBp/VoZJ7CZdUpZdpBJ8W1qJ8Gm6iqGi
BoTpFo7UQrtPcrAVEDQBetC4bgAxs7xdsaW5jOGa+xc1tAh8SQRQ0adqAbcN
j6m4Qd7DnwTaHeJoMEB/ILDZ+PLl3bnx5WQqPAb3QHk8cK3E0eR0sLZaNvy1
ThRI4HpQBCagplbuJlX4xBDf1BKosdm+p5vF4lBtPU9o5hdLb2h9XgFS7V6b
wyMwwMj9LScgUjDNhl6n5B/7XDgeytu6jk0uMVPArX6YWHpETHF9j1ZIJ3HV
HXkfcCoGk+EJCDvDT/nFSkk4otJB8u0fWHt6ICWUfDZidiDFYtzmGtieze9I
bp1YSyBKY5E7KkmX/33x/cf3GAUCbYL3/UEeNbEbQkjuvgiQcp/yu0BXf+vX
GYwre1/VuCHyE9AAhgSlJ2r1KI+Cr9X9KrhInIRzRFiT4oMXrpI8gctZ9b5U
YdwVDAcIySuB3KGSM4vmDiQhMSQu491A5qQO8ChZIGRUvA+lcZq4jmd2foJk
DL2wDaGuoBmxHVjKM++TauWAubmJ4nYM5mobu9HVNT6OfbBkF7sUCL8bn11x
tUABKS/sLOH4Uv9XrXCD2l3Kpc+AfknrmYhxj9vuzHKUK8acFN9CeSxxPrVz
imMwLkewIlMWpvUJa5toH1muU622U5WLuTvQwrvO0EoZUibMyCRjYWkqcsGu
uD0aoPGtFTVdA7AX09/4PhKvJuFK1ri74LSJiY5xr9Wep4mY1wYHsdVxTE6g
5CvJwIVupSRedcleLRkoKbvMMS6wVWczvKUkN93yez81Ywk3J7+lLW3roOB/
jrqQC2dvA5qEcwNtBjKjLLGHdu20BBDvmjz8Xt9S+zJAB9nscumCDaiiQq4O
7sbDkLHqVcGfBrrygImC5OmT/GDQ7CEsdb0XIDdttgzPXpsK6ZU4VOwjPEki
cn3x0Xop+TVf+uo5N48urjm2DiHN6RxvHprLPlpdondLrFli/YOABXDaOadC
Fr7pFeagIPikiRVHxZiBs8TwW0ZebUV00d7Y0PUH6O+Hrv9hh/gH6EMyUwtU
usn/q3Lg4kQaSzAdrh3qjgZRVuia7R6Tw2MWcUJYniQ1FljjFJboX+uLp+yC
LYpzq0SUEAjHSqA0JMnCjiC98rHSMMdboX9vWYKx86Dx1nZufYe1rqyPSPNB
UiEKYT7mfr5EEKAs61qiYrsl9o2ggywFm7lTECG+qNRlE8kKvkQoOtQtmonH
rt+jWIr4WCGZNXAGI9miLAUB6g9ks/Slo6OX88Ti5NbaM5kmtumiibkEVCiT
wiuFlskRG/pXRmhufybyNdVgf0kGLJiJb/A+mAqW2Zd3AqaI6bOoDJmTnToy
6oCgkXVYYgy+mBjaCylzkCmXoLocLbPfYiwdzcagAlXXxDH6B/WoLjP+UOqO
FgObYz5xKUBmGzTyW0RSB8/c3Lm/Mk6qEKlvF9Pp3yTPvQ7MvJ4eQ01R0NXi
Kxhdxu0ihWx0KojYDDx/1ZlfFGzUf6dyVr0AEPtPDC3Al7n524Znwek7W/5r
TTjZyVdv+tG+OurCYTunEX5VA9jqNu6fI5cu0ymLPeH/xFdG6UrePZlSOqNv
DGrcw9fT4EbIWHbYpZG3q0/5mdg8lNwmsFzSg2+t5LD3WA4pl9dhWLAEkYBr
VY/f3XWtl2qIvi6Q32oILlKBQqqBNr6uUv5O20+OlhJWAOfT84kGzzPqQdSg
f+SMFs56s42de271cYLu1ttAb0Q++ZB9ODkLgohI90Wr1Ud6DfKFVTkup86/
3t47rxJwp6v/1eln3m8zbKTTiL4/n8kDddRl0SO3W0ubQz57bWbvz5iffQVv
ewMdvPQFc9MgYudxc0QKEVvA49J/BBQPnFYrOKOrWjR6qU3oX/TpCVfgjWeX
qch9o+NHfWRTIsc+D3l2DmKJkDorml2IJwCR6Qj6d0ZSPfoZK+ANW4XJL/2d
xmh0qufojuk/jFNxQUJ2/AUaeeVf7ECZX8ZQbljmnfjGnYlc9bU1X+Kj37xX
Wm6L62pY3ENX6kLmQSlcIuXqXo4Hj5+LGEIfYx67Jyr0f5VZWEEULC7kMsFW
ULWSygLxIrkSUsYl4cbIuYy9nyXJNSNAg2X6HI/kxCuDPCLxk5Fw2mc4cUrI
T7kcjzuZObZ9ZioC6D6ayxL6QlVF+pHUKgkF9KB1nnBCXS8b0hKP4Ig2mKaL
vuUYVKhTTydzZMf3H30WeEnRJWWR1ZRZF1Q9Skxihp09WAGkmX39T+jO4LhR
d+D2pmOLJYVc3y4Lh5GhlG53HULm6mvQaSSUlqHk6P9z/J5dz5ilT/giNuBN
k4A0YT8JYJo8K9TFejnsmP+ZdRdWsGlVg+euhjxFF6dOR1fLwfeGL8FflbUT
Gw1fGlC/zJeaAuItqyTK80Y0BJuSBjn8K5GsYfr3kRS0udf8NcrMUYf9+zYk
cvYqRoYY2bXqGJBHZiluStXjSrPz/YO6j4AvEhLnJWGBrBJZVw5ZPETtqFAs
rT+LVXgArIPvOsa1G9rNG6Ans5HpjLZixAEynI8ujvO7IzY9pH90AGm2L7Yz
KkaaB2NBcNd0aE5YL6o3g9jZY7xx32BngrwJC/Nt5W6GQyq10AepvCj/Ii3i
NtvwVig/GEaF94o8AWQ0l0S1BiT4nLdN3dpoKtVyq1Jwsvt3GmbAHS0zuEHp
fMcOm57gqCiiZkMrvMFwgqBdhPgZkkb0FhnYDZTySTgtevQz75G9GFyhUES9
op+DmrmGF7bcEVV1Ms8d7orPXLuuxX/uLiSQ3mLrJE4uSDhggRVtJz4PX5ry
57WHdl0QOGthpo3OvFHSntv0koItLVOfCBMhaHMegva0OqpEpP8xFXUlkT9v
vHmVy2G3MpAtC8ZdDjrUJ4xZx0i3ATErorqnZ2ElkK0I1EFf+L479g82ogt8
D9a8YdvdRNOLIVNy34W9WpWP5Gw8K0GAkfM0uts3b82peDoLi6Q4GvLL/fbB
a2uWTf7vgfcdLW3i2TAhQVnOfiDKwNNJ6PHN6Z8LZlFVeuDb2EHUCTC5r1+w
dHcuRVweOKX55sh8HcoQEA2+tCi/GQeCYbdyhUtZ3+ofe/Jr6GC2hJT/EXWU
AVHJ+moN+4rRRN3WRCWQ/pD/tlIOFAIpk2XiLwfqUG5/v0m0IpL6SH5xBU2U
GoLy78m1n4nA1MTXK7LVpHRsGFKFtYffqXJuedz+9KaMYLR3TCw84lgHHEGp
9e/sVUYbNpoEClYZukTcqdCxTGV5x6HsGDxKvbee6QU+W+xCnD4x19mkjsbX
FPSJQAdUNtorjq9Yo9/pN8lZq8gh8917iSfxHpump9wOIirE05BsPIpE3DCb
mIHHkTD4U92wwNVn7dgyu9L6/YFmlVyknilHkRL4yynNBbcjyNu/GCGLBhEc
e4a/TCiYrnhKJwSCwmALl9SbH1gvSlFKtp/5JlF1/hP6od9qx4yk/3RDyXaV
0dtusGiKIxfNCo75QSrW1EKpYd1nXRnKLNqiZlkLECJmO6HuF9jSGiTOQfQG
J4+1bJkWv+XlQc1RG5rK/3vx3yNfsu7viqRyosz34AXoPY4l7JVUObVVCePR
nuUOyKGWww0aRHivFTKSccaRpwCAUrUgGzW/uQL9C5cqJri5gkbcGxTafrrh
48nt04tCE4HD9QiUdnvDqprxeWoWmfApc0Y2IXjt4z9xEdYpaoZUkol7ARbv
NzaXpnD499S605yja5xs9nbXuJvWGBENTcEINmyIkehqHxjf1oHoKEtisxsc
6lZZoq4Mn3+IK//crcJMfgPGhWhofDJrK2n7FVdrWGH+TZwG69/R9O4cIXML
V0eXTejhYcRndOYCya71yGyTcDD92TOc/NDPFSYMw5iYuWmfpTH4lk6r0b6k
qRCHxza/tGxU+DtnkAQyKKCSnHLOitiND4pdkdClnpugVpjLgM8JM2OGBwhV
EuBNKsxmyKkp0Nrr56me8cUMmW91Jp5aPQ/qpiLqlJAlGIVWmSIJDnUJXu6J
QZO8iKerk5nTVEBvIUeg6Gz8ulKMr2j8WaikPba1+zsDKbEq9pQ5USQnmPyT
syH6d6lT8AaFHicVvfZG6DJeINrObCF2bKEhJBHErEiPavfUd6TOIA+obUW/
tQzvpF8pTVpmgKdMGQQpeSl2QptQdo/uMggRBKT/FKbHC3wsSIW3T2gqK0nm
9FecnpimNz0gGDKe9PK9nYAv6RRE6+JoiK8WIm6pqhp/OxiCZs9LJQoo4aUv
ataKuQqDAnrKaghhiHqMOkpByMTgnlMKKKTsPKvNS6E9TPt0UQnwCDeAltkO
wPVxEkLLS5G2X7tV6OB7c1HEohsenHhYoEKE+eFhzuyvfuPO2UJLysCE6u+F
wukE/gQHK5Qb5Zh7Ki5bUI8fm7rsnarjGpDcyscd0pk63jfVqAuogLhIXDdW
vksP2hVDK/PI23Z1TBQVVZNnst6zXY2MF4i9YyiWZ6OBQdTkmFZ1tOgDLKwq
Cb87MY4psw0KG7uhpPPL6jJavgkBoU8VJn2mUOhcD9JFnQqgS61c98+EVkeZ
AAANJYejyMgsv+NMaV+AD4rd2a85DjSgnUkeGrZjEFRrqbs+TZc7MW0d0u7a
lBOZPRYdz3JNGKk7kLFixvjUBm1SepWJb8TXpVGzD7M1Hep+74q1fc43E78V
na03i3dEEVpfUn/RlRY+Z27AEuXALh0uBuImv7+G3U0cQjqOiwTuvCIGdbhL
RHz2tDaKzGwHSGZYzV4J/ULaDbp6R1HxdG6W5o8ShDJmq/BPvyx98cAlyBk9
DkeZgiTEiVyavJZ6o9uOMX8jfvPBCTiNIPk5/KQ1ZFex4SIftyZhLu1x0SLW
2BtGvSIycOt1XkbVeCDeUBr0rWr08jcVicb+P9W/gBCCxtbMl+YniE19fjXv
MCBLvnwDD+tWyIRPSo9tCjG6sZWu92g2hXAK+TuCUPECphzn98GfblKasaBL
GAgZbJzB/vXiX8/Knk3ytQ/L65JHemtORaAWORKag8OuYyxbDRLAuZEAncGo
G36flRLQAh6lHA7WnWgg4KzfO2k7r9vo9565Gt+a9CjUiBZF5/m1DQyKHGLl
ZtrCbVva3rkhZxcb5jJBq0BixBLhfcp8AvEtYfHvhbdyXMmDh7a0LUANHqbM
lNWQd9xairpN0e72ry/i8aVx2KEpi1X/ihvrlvsvsyUnwVOM3jfEulWNvSIj
XpW1ByH3wUWoadoPk2AsdDOQd4aRtLHdjC3LS2j2yIiaYMex6hh8be4cdbpy
brp22MeohhSacDKby6jzXeStcIS269O8QmZeeyKw2Qz4B0c4NtupK2+1fmxl
6Lm6nah/DYp/Rw6kKWAQd1kCvP6fM6vxeNNmxU4cH6z/rfNPdXswuNAApVyl
11ZBNPyfG/RObNFl/iSo6lY9ugkhmF9/MiorJyDUJY03NBTf0kEQW5s53LDb
Pgzhw/ZPwgahcs++ScL+y+sC3iWGAWePwCDKcmnwzP4j5kNSig1p0K6VXCbZ
UHgvM8PSLbdX6IjtbPRbjdR7+H2vKieSCgRRjrzfQif8HxQVZMeegvFBGbSE
jmDjnCZcJKbGu/bK+J/zfyXCbiMwLvIyp65Y1NMF+kb1j4gXbp3ZBQ7ALv9x
57LPKzMf4D7ZsFfMoY7DJB+LnKOr2934bRvR8FHJLJAezeCsHQyw9yLCriEI
mpp5meA+H4fmPxzlpm+XCu7kaHDz+Y8rs9/Z88hP8MxG1TOHRGqhNNfV5xDc
P4CPR55xwA22h1Gi24iPeCfu1W2sLDtZb8y0lsCW0J7OGAa7bdh6mRzg6D88
7+eicrMIpwvY+OQ2wALigRSTkR+0oWY+SwlR83ZWiVRfLX0sI+egSG+QLghg
VTozKVbYzvR2JLTMuhtiW1Xa2FMs3pWf3N5405kGAh0Y0MF6Pg6nvyP1a3IM
D8470642MPS65ncSr6t7Uy8cShQRpe6LiI/BxxCrYHtHOWykuo/gQ1nvuoZf
K9V7pIlYUmibvybnETQA3rXC0YtLK/6oEYiySUzdXQXgUhrwm8GQINFqrqZ/
oJ78OIaw9zFHbFSPbNzLrNwvtyvSD7W8CJBt0SCYbTnR9jjI1egBEFFi9vaq
dk2GSvahSzrNx/sp6pBN7jM05eJzv1YMCxmcbGNoc26ZSiiogxdBpyQPmxl5
ZbnKIILqm+0fQdMfQL2514/XiPskIyyw8eoceNnlwgqG6BW3VJMEXJ7+SPF7
8QeruoEHx+dltt6Pxx2iXusnHFVaBo+OJVpegvGvc20cBG4fbVagEsxJqWbV
YbnjG/8GXr3UL0aUqugOaj3lEA95jX0q2iWl1y2ueeZMZHjc80bQNIkdPk++
w+pmXEe0qRgEEiPehUeH9mWKhXZhZnj+7cvTbXupa89Esk/KVGqfdmUeY2uZ
Ksn2514jkA9N1g01ltW3XbJDaccDRPfEaW04TFxfCWt20HdjTpHrDqLgZXp6
jXh0z2ORkRIvscqx/dhcoQgk4zuf31+8yqbD+IIN9kn1Adkc1Kr8PolbhcxW
+NWrc0B28AHuGmK8iblkAAIv/ZUpreJDP+K37rgBdtoIRs2kr0+qLt+xzaf/
zkJ3nBOGajjxmAvLipCW4ai08I4rJhB0rqVqUZhoneQgFNB2AobyUzeQTCIW
HhhJSyR/pGoDjJvu+tW3hWkbqU/i7X8080GDAmU+8xJwYH8J3faAndlHrcb+
4t9POlcmC5ATQWdaQ3AetTTrQGBzUfhxamqmDc9Jkh4QscTzVfpTevHP9/Si
hSLWGdFgnzz7RvK805fdXJh7mYm1TbvxvMxM5qyf2R60IF1YojflLgz3KtsV
2nCa51TT+/sAiQcds2UrnmdVTBGv1hbAaLejS1iF9zMv18mxFLbtsbFt8aSe
Pka+DWAraJj5J5VDLV/6D7x+U9QcjwZyWI73xrpD5HtaGUlhQT8YYo9tOfoF
1RMs7WxIdWvqKY2LAttghJTDaHCazweVo8P8S9lqdaZeZHKKsPZW4hyv4r26
aQXLAKcjKZ8cNtKV0RKOw0+wK+h1nXhHbV6Mb2Uy/77sI4+27sZYiygIyaHE
9JgiFTr3w8Ba20QubQ0PbgijKIvDS9e7f5hjj0j8slsBvZRsBsGt+OmnR3zP
zp1q+MyKKaOT1wQ2SsECHLZ1AbOlc8jlNvjQ4zD4SWlfMQkbNsFkFB8fsfPR
Z5hOWHoRuysnSq3GuYHInDy+yCKJHKMnGszuU7HphPyCzrJ8MFCcZdJTBsX/
5fIqIKcQgTzmI6EQ6IoLwcXo9UlrWO+86mr5YB6uFHKCF3VBT5m/r6fNDtJg
8NSTYXBVypT9xQ5JXzHxqojOPHScYG/jdutQF2cRpq+CI3dErL2SrMs1rcIA
PJAsRlzgBKOa0U96Yq9bB3NtDTp09pOGknbHD2QEH8uOCYuGvT/7N72Bl3iQ
FI6ULmhTULxwiW2pEuZJ2/FdfwPOSNUbBOoS8yH1tWY9viI3GnRgQfYavMTL
j5ZnsoedFr39i3nn0HCdJIy9AZMXbenLAC8YjAU3l9HVY9oGyEIJ2jRKO4cX
qJJp9WrFrGjPqcwrm9EqnEOHOHaxip5Nvb9YKyikWrp/nP61Hq9sGe6RAH0v
CTiwVFhnBuXt7ipcW/jbI80jV6x3OwcsX8fTxPZoXuPmL3+EzRHfUipXTffE
MhfxlkHcY69wqalUDV2yx0DfkZC4yaj3gaTan+xTEJYMc2vUNCtMlPXKZFo9
51rrRMCQ6EmpU9P7arboAL8zVFTV9imIRTBQPhbiD6dzHa3UgWFsuglPnaFC
9swGf6j/rPY4x6hgBSu6L1gEmQgqqWyuEUiqbKcesXL50i5zTz/B8WlAKDTP
auqxD3KszcNPHjsSE+c+yS1nbrJW/8Fv4GWSwyicugRF5d2Ys5BZ7JO83tMC
jiq8Dl/7GhrFtGUvlID+u5jjzjHIkBE4o+3W1XEc5JSpIVqgWJdseK9ew5Ff
z1snsR28/1wBWl78SbED4dFe+7lvgbaPWgash6v1ZOo/yiElVkA8cfxDP1SV
/HYK41aPV3tvjjqnj6h+lcSLLp69zEufmPn2q1QemxwbvnJ9SPDyaZn1vuZx
CYZbMvE4C+7SC/IFtMy8Ut93Omzo/F1O/oBoBu1DG0DD22srrOimbPELrdTJ
ia6raNsL9fX5yVuZGpCDc9Dmy5cZwmrdxVX0foc/mXZAYxo+I+2vXGfjAgLz
rswFCS1UFvlIM4scIuQNNCGx9gERsPrOY3EQj22vqRfVxyX7zcw5fz7tXKnH
/MQj1NWCQWBCA2p4xhv171ylI9zTstPwk7d/nQpQPgT9frFxiIuKJixmWVQw
TH83IYO3ZwGu4scy9JjzMwuHi6L49DuHuUPRicOtjO5QNYYBlKaR3rUoMe1g
tQWy2R+JcZ0DPs1hnJm9BalZOfCKGvOHWx+1KRVv+N4JzVDLkZV1dDtTmN0e
Xp3UgDElF/KnvfTvWEB+0LLQ1G34m0nn6s+1PBXPR4vPuq5X8Oi31JrV8Iy2
x8tPUEcJnAvXNwTP5xgC0ZQAyPJs/0lHhEuQc2iynOHeP8I4YwbBIuFyCxIS
LvlchUZpIigo27LkxtTO3g38q3ZPMLusezjwlVHfuewV+3DolKgnw9Lh90yv
RWNWlYsy9UIZeYbPbI0eq/ktZNf30HPto+IzPTGrOx5JZofuMze9tMdAGxG9
D3SwZjJ/pajYBs+8gJ6ixYGrxr4UrSBtp/ooL6LteBUmKJz3TUag1t0rV3qD
XfL7FZFbglLIa7DdpV5bX0IuVo9VangEXxAIiV/kEXWsUDC339QBBVPHY8X5
U0kb8qEncHJZiuAM48jcBHlws0eHLtXkOxpaDGFe5dcZ1Xj7EqjLcp1x3DHz
HYaWCCBM+nSo/nsRLzHdvkH4ujkqbq9ZZ/uzHiI8/0uOQRiPZOhrINhBtF/P
JXtoG32Dkp3gURiKH1/BWosKivti6j5NBP7ABSUKvCSRSDvDuAGYfwoFixqq
6x+lz5nHFJkn+g/oxZATOld+cwZTIxW9sV5BTOT7JswCISnfMmC2Wt6koGKa
SE5H8UO/N2j9RILb/M9BvKRvUIsAGG61Q0nDBNfom8gpnmrnFijRQB9d/pHq
wmNSunlzy5oFD2CjEicsTQAHM5Ph1OePzYk44/OPZEFnPfSLh+iDUvXMH/Yl
8YXPew3gRionsKDOJK4w9QA2LzALA/TMUaH01vZa3JuVbnhOmobtXtMhJvJN
yK3rVZBvh4FMnTvivkXhR2MyYTGnmkHDmV4G823Hc4CywvMaHYY1wzWPiekb
WhCvSiNOaBUURfasDHY5ezPngWJwHK5R+LsuymRQu1S1XCDnUlOJZFKwoVr9
uEOKqgQ65ZyjBbgk4yxZNwe9afqPADliDhkIfbMnbgsqhoe2iM4wtg5z3z6r
6ra4/pAWOtQUTyWNXPE+fUQ0cmMb54pJrxea1AXz31NP/RYw12DaYPE9/5fr
qdaFU0DKdoecGk4zjRWuQwSM65v3v8m4T7JNnA4jd22EQLdfvMxZKcNfAovo
cLpBu34M6fDSwW1pcQDD0szrmR2i+/m1Rs0lSA+8ni4eTq+iemx1DwjOuxf7
Lg9OAEGzzEkk0tandD7XihDkZg67CEohGhL+bnUc6WXbMc/JGtqXECu53fKq
R8pJdQ/mLyJNN7UttSt0k4l6fAqsaHGhdGh58gLdr+bWWDl4zR2SGsgNofIj
TBgyRMpbv1ReZ9wHptw426M9ARtXux0yuLWKlHaE6DFskM3oMvAi0c3NoHlR
fzlxEuhzWeIUD3DqEUO6eYy65r43K7RIWVxvTvxQPfKc2VudUVGY7ypi9SiD
c5u83F8vWvX+nceoD9W17oDn/pXaGZAu+YAkk/Th+LX/Jz78tYZNjjzlcmka
EsOSxmFtWjUFqWKT02ZW+TX4x84kdI8+YPTrgfSMvQerVFSnLl4kA6lrF7+q
yUnIfkTHFzCUNve1quc8W5tdgSfUaNjkQATZbufGTf4RpC/V7+EsXJUm3rkG
Y3vHGeUhbPEyL2PQ/ILGfzVDWzSSymwvhsEh3JnQhXsxdH9NQbiX/ZWtJETh
CV+CVs+8H9XFKIZaw7sNczCL07SmW5egDEiiSYRgKAhL6H2OqFsnU2Xdl8rm
JAgt+sR5DQYduvj/EbVU+yxUgOGa9AHWVdXkdoOQgiGta6IyvHoOoAHjK7jh
53HcfUQ+TAY2G2wtgGB7UskIrXiwnvdtqOy3hF/B2uZfnxdOO1JLMAINSbMR
RW5iBzQey8BeNYtoj2ScMdHjWew1e6bCa11mZ1WPaluMWWQVviBNLA2JKeTD
ArsDMIDg99mTXli1989/OEqUdA43HXzwuZ42VPXnujCZvKLipyUR/j/PJT3S
ZTGn0gYrOSWuAvP1orNC3o1W0DVkBp4msWVzXzbh4Flx3CLMYGitmYLXmLeA
n5fB3l2XeFwoUpOJBcUzHcf7Y3XYKcCE1Il8N3KNMNeiSJob4jdwpJaHYOdk
d9rhwwL/LKrjvi5DUOP/xhFKsm6xAjsjIEgVjJ0ngwyqtKFEx3FqcWPefep1
yWOONOpjUUyhwxs2f4xjDpj8AvtxQrcQUag322kNjoRrR6KMMIasNl7lb2u8
CEspBn6yGk3qqtHA+QxsZKr64EoKgK4MkhADYWqX0xD+yEwmE9x2XSYR79s1
ol7+iUkBddErQ8srAjbIPr1J+Sq4W4fBQMi+k8ZjkC0aAnGQ0C2/R3F5MJFm
OeoSkzueSBdgt+PmnLpn1/w/cYpRqP9uyQwGVlBW3fx2VjClLHiOB9ZZkr4a
fFViQkMgMTb1juZSdosBojKHIZ+oP3afdgMVrsfULD8t9LVcR6g2KoFeOj/A
S1YZvkOe13TqfutC5gpbYOJspBtCxxd0platBwYxu09RfAkVbetMMEm0+neE
MY6wCbktjP1fMkUQOxYi/cnfOW2Qo8dNBSUNdVjWmQu7FtHhAet2wJ28l0AJ
79I/ml4r02OJzon76ZJe7fFjwPIVbPOGdF/Rh8nLDQIO91qSZp1NiWSI9hEO
W3GD6ksCOoMDa2v9B3G4K5xcLaV0OlPXxiyyq4IXUouqsKJMdfjQH/nxoQ1D
SVdIlz+CsyNNAgCFX2v/+5zzfSzbvez0oR/AXpU6Jy3a0RRTdF5QMfaqKc1Q
IcDHy7fGlwFalkB/IsO1hmFY86GfuVqZdMnhDx6kb/z3HEpS7XufYcwEWc/0
UMhOVU/dsJIuu8sGKn3PaOSMtytXzRWZMAU822eXQv28KgM420VrzBysE41s
035F6/oSgS3RZse/Nj9npuZgPeiu5CrtkeIPyHSb3cnBnSrAx71Ru2QNpNtr
IbuyO1HGmsC+HuXI0zbrOk7CospKG+mKWwHsNWzjP10OkcUbasQ/z3hTQk8e
ge1P3l1XLZGKipW6Al7P4TZskRnh8+UjLxZMPy9VHu2KKX5pVfdLaA7MpAEI
pyfXkRhWf8QQZcLVW2gLAb+e+sFtAuLOZo8lpW5RQi61NobD7DYdfHklyYCG
j3QbtQz9nDqW7qnOUmeQR49jqu9HYzM9iwlzD92GD8XPrbUopYEuyYTf//yA
FP/sse33YaX0tTNrpTcEsxFQMW7e2aD7HdinMg3VIyVIlY7F8T+yAbCAahaW
USHnXxWlD2iNrr3B6xZaV3tRJCenIuowwlKy3K8wlSgJhX68t4EhNJhMhYCi
ysa6ru0RIX7v0jWaqviIprL4ONRCfSFiwFTRlOr33l59DmJncRub99blisin
Q0eIhM3qjMdDMuMifVNxvQbUvUE15nzbQNTeUSJoWbvl17NkI6Kebb8libFl
6nNxYg/XoAcmBL9F8YE/xHF/BplHy/Xi7NPDqJygGTiMALXJll21NLWg2cuu
MdREUwU6lheUCzE/tIL4jhiZAed/Bsgq5SeVpGzr3LCVWXiliYnBwvYq/ubp
ruPnfNrzr4eAT5/zMyEvDABzRyAwGVh5GwdHfC4Ll6YAhMOu11uJBV8q0tRq
KDYrGHcbp1wHNAUkb3LLSm/j/Z3xf7AEnhQSl+IF5fr9+YGXeRibxI+T4McJ
NcDYeqCNgwGcm2vY11B6VeprUFNk5tU/8iLk+ELrlvz2VZdCwpeoUtwsW8Xn
H0i7zX0Gc9V5MAGeUHoa5vKlulMot/CQullI9I0DRIKG43x2DCfA2xI6gb/K
ia/LvGqs/lASnge0qhe9Teo+1/GBVZd+yWFqveJrhCXqjlFdyem7wA8ZWoQf
qO3B/HWcFlJBonplXmg2EgDqDuzOPr9JPC77Ev9WdcaVc45rnpTmd8T1uLg7
4xJ9FX4rOscsmn/i1ntmVcgqpSki3EN3dykV6/EzA3gBhLowHDRVq4FCtme7
tPXgEJPsJ2gz7Vwaa7e+hfOPpuWEuLcB9wv/TiCuvjiT0ybSruJsfxBf0H7L
e1Rr6+/ZVAYCnOR4K1ojP/qTlN8eCQ2whPB2Gxf/llP8E6mzqKWgA1cSZCD/
cV45QjRF17Lsv+17VHY9jxdU7XjTVjt/GJSY+VhXNA9RboR9U/gjYJRhgv8u
nPkjy5q4tUkfk+/+dMn2CWGAhuqP7a2KytM4y8Uny7o94BV9AIvhLd0OLFlZ
GI79Q4esId2DPUKRvH2pVSW/lqzQMHaa21NDLTYGybEMTYEN5dkTv2JGLYtf
HKgllwLgKJULEM2YPj59P+3n7fjj767GV8uB1RZ/fzwX3AWYT/Jt1oSAyJ/T
byE73bS52JB0nuwusxlXS8RzEmcnndkqAtsFuUjrJoKuqj+AekYt1kS74j/I
SFDyKgdeptQII9Tb7pcdsIA+S2iqFvTIoYqN1djMj3/XkCv69PdzYMaXjsYN
FYfkDihxwBXgj/yyof7Uo5/S6gMVeDwUCkEmX0i3Puml6noaiGcHuSUnahBU
kwNjDBNvvLX8OddjvKpaQI4e7htpHnRGmNb5UvWvxhMpBSNvSuoaeSl1/F4h
469x57y2kLIYcRwQyvN8rWNFVtlSSHnKbNB268DlhSAbU2eyhseKKSuC6Xnb
PjTiXep1WQhEhSBV8Mh/Q6VyO9DK6yHMlh61RYiyu3JDL1jFsshjsmgPaLlI
73RlfxPLof66DnXOJiH5+ztyj6nuSdB0fx48Cf7M3MrnzH1U6K7xNqDtmVER
VzUPZygC7wq6RnVmHKNdklKLW7ZetC6hq9kp1zP1vRuGBwCIPXXlrXLSFl8j
/dx07lirnMSQKlSg9j7ToZdX5773Jls8YRqG3hIQN6wTRXMKF6wo86hXw0d6
kJw9VpZk8flHgL3SjkwO73tXXIdXb00JmgR+OfD0eWu3gq9BE7upoDD+09PJ
Aj+EyfuHM9HxvSyGjrcXV4KUyECkgne1O2GybthQP4K4ree8ZkIkpdR9++n4
qlwGhRe6DpD9JVk4/oXzXmjRfK0ItJQc5D9CjzDu2kYNLZ55ogy3WE6kRrpL
IQt4szpALF6MOr14VsEejxJRG8Fyueujcdg0YcNJ40kLOZodrzDcR0LxfaES
Ls76d7pkbB3vJ44q9qGjldPZMG05HCP2VPjDA1wN+BtVMyrsxWYXtfICNgUM
HNhiWvFpB3okTB6EiHHAyS/gcyR5I3MHN9pUg71aFboH2vl5OnL1a4aQtvsq
8o1xM4R59RIJXw0d/fLCdlSmG4O1K1KspkvYcaRomYWy2rpnZSiFPWVJpFC+
LPUSL4vEYwXOZEbRU1ZS/a/3/A8FfNuddT/YmOk0YwvaHpqloeAKkBPkzsQd
KCTUq7YOZofn//Szsn6vMiNH1loJCNasrd+MyUt2os0OB4BzBLfkiDgx7Kw8
9tLHE6jtJHUyPLTBn4IauWOSJMRlbOjNExmBvRx87mnk8wjQyvWh5cBMXYMz
FLeGId6Q8eqmd210iTFP+0SlYDdakY2pxqY7KFqAd8LeSbgzmJ4aCnutH9Vu
1snh00LfAMxDKS47RwIWtFaUJ5/V1mHWHHk+RCgR3GQF0tsp6eNXmFhWcEGX
L1+S/kU0T7Pky+3l7t9hz5o2V7ZarbPZObjW0eKDQRLbxMglW/thWBRHploo
nEpEqX2SXC9GQ9v8xWmj8FFzZNERLrr7X+iQe5pcZl33kgzd/FTsDBVk6Mgq
K5NtQdB/4ydDQ6YyYjkqirZBJH29mztgRRCFP06k2h/CtbB4PFa0WUcimbgI
JyLAzIfKiZNWmvr9gPywmIApvn6fwuTbQ4nrrbqX/cO4QvelEiQ6yslgO5CD
s3qA7OCFLvCI0ZbkZURXWbpqwxA2I0ZmfQ3gnSXH6/9YDgjtNxDKSAYCkP2M
apaTy1fzjKrL8dHZuVnKjP0TyienbC8GzZm2VRU5EmeQ1kVLF8x0wiXa3Jf9
Y/0Taqp6xe4UcZ3x2IH/ZxUL36n6BK3/uzGKK4ObcQWy0vyIQmEHugMMb9D3
SRXZTx2StuZgXhsjOmP6n7wImw+PrZr+ms8JC3TdCNg7B6v+4FITPwuoFmt9
I4A//6LAgQlhEufYNtsq+h0g1fWam7h+0THmswEvXj1a1m3W8g7GVgrE4gwp
vJhczxvPBJewcLXPIdnlrVYB6i2lI3fe4QhpIdKgp2qg18B3/xQGTKNHC0sG
Grb1f7Q56ToDzsKTxUOzLJaLdonhiqIQ9hYEJbVVJgnb08MFwbRYbojTYT3O
oROzE27Pvgd4W/aV7jVuWE5EyiuS27jQoRFwiJLWGHwcs+a7BnMC9uLScSbE
bzEGNIM1Hih7A00H1gxykrSNFdlgRkHogm1DajTIFEWehyw4Vu+R/c3u6p4k
vliQP4KQoTumoJnKzhAJ9TWAKYh9OpmxhKFXPtlbyyloKS03UjqLn5n/e8dE
3rpY6/kDw7Teudb6vaHwOhEUvy39r0+vkcVZ2zJR9pRL66B4yOiuCkXhN+sj
taVGGy0OWsw1nE805uPCm8Tby9sQY7bKC1mfslhIG6BqsOc9RGFTs83vZzhA
aaGe/9Xkw/ngsTjcOjKoozg+qNkj6zEmvwi5ztb/1M0ONCXP5upHK5aRhVLD
1qClIY8GDGMyRRMknZAwoelzqK/OH+nGgFizzEpVjo/4aubv2MadlDanlGin
8IxILoU2oIXHo7mOf1EB6mUSlLU=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfSbU46IkJ+AVqlImE1XEPSl/ikvxOGRjYuORHvvBtzGzh/7L5tJkBnLhnpHXu/xBoDweu6tQiWSUuT6Og7bmWtuKoHDI0morYYu6CUZ/oxIcKuswrywTnLukV4n9w4r1QgmwkduUJ1q5+uRqi+Yne0fMMvLaP1sk7cVwJLc1ST9NdqIcbe5JNutdH3W6d1AWBxe6fIxZNemsco814Hxg6GrXcnNMuGYLNZ2j1ZoBqrR16MCOW+nxm8X1t14Nj58AOm01IkUv1JRgzloG/vhnsMGLgQImHgjFTAHcy45l1xe4uN0jHH3t1yBdeF3LxPGEI68aHD2UEw/0AUJqLGs47m/IThuWRK/Ucz0450I1MWn1w75Xt1sezKGrZOpIXdDGS9ND4mRjFMI3FUpkEQOmesbmCISmL+HSMppO4LYR4Thb3VBOtUGgsMDgie4I7geIow7jZQ9KCFPFaqOuC/uDWMkW7yyI29nJ+a+WJIckr+ijXkeH6CN8FupViHPDhYJeB/l8YCFcBC+EuPgBCG3L4N+Wyz/VTwARZRN5/TWQNvQO/dIZV8f5gdZUyacrQPKcqwKrDeH97E/mgA2HIqjBQqy9ECUwFpQr3XpGfZRfs4UFqk7b+Pw2w3jUYF2QXdBn1E/GnzRZLlvKYxorLuFtYSuaPvX3nEESf9bPSPRRlS6D+P8EDiiVvJ8eVZw/EeSkiJBf0Ga2Yu9WuTJOyBeEdouHjSOmm2YGXf5n3GWWeaEGEJSUTkIEOvcroKlRsOwESiqAtNmNe4ozzutMrfMzk7q"
`endif