// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
cyCwBNN80N4ETB0GFCjK1pxgh/wXYYeU6sunWAvW/MAMOfoYLsy6lBgSQCeM
Y7Az8dGSekTh9wVF3He/ULoYBZUXFQUvuyk+egaglF0bujCoYu2GDJUHrL3I
iCl0gzQegpyoyYQ3V7vu3CSX8qOGQ3ztoP9+2EPWBfTh559oyVVpFNEDzft9
VPkKx9CzgYr7K2jqJBbA+kiMP//DmDjLIgGmguyWGWAffq7TG6Pi/dW0xxww
Gjgc8s1a4dth9l/X9+ofPatmG29p8m36/Pm0hp+KrN3g7Yv00brpqva/GIMn
b4jyCkWFHZHusGj3BWsKEByAKtLnMbJQ3MOcpgrBlQ==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EoYld/LBQ/bxIib1cY0faXdylHmwe5dFHCgBFjoDb0/LAFsA71nwDmwO7BTC
KUC6CKfHIS9Z3ORd2WAP295XrZlouKkvMAPy4HgAwQkk4WylnnHzOGMEea4/
4bEd7J0OwTP8d6A08bY2p79bFRZdbbprL6IHHDdTRxJnfP4r+pCE4arQ5AAS
nJZrLnCg9Z/FP8035Bfc+mBrXfeSSpXw1XHs8YCDMt5mdzpWz4EoIMkiq3WF
Adgkx6P5TxN1xOGcvKYNCv+I2tXUguUsdMp8A4bqiAkHTAwe23bWfCyPDzPC
EJnxFBkWSj8NlxJF+E5fC30MPycPylb2SIJfbtqAHw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
E99+58tp617oBJ3k0IZcDLnIF9xEBlFqyfiZ/oQF2X2uRmKWJE1FC9MkAhaJ
04VstuVcFsvxO9TW7MKFAZiaLlL8qZGwE+a3cJp0vkLqvclMtVLfoLXf6On1
zqfwV3Enx3MMvN5hFVODwSKU2byH4iUySA4pR0OukeCbzlHIw5nLD4xRjtpy
pQw1b1ycOw7ol7BpSZj6uCSp07hpXZ48B7zbXyuMs02SsQxkwST7JH49GB9O
WyT5bzh0qcXn/Ve/tZsXpzWaYQk9Rh44DDosBxW7D9Kn2g3uKlYxVQs0chKd
vtz9GpROuX3q0JpWln5clRIFIrSHRNuix7t8pRBpjA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MmHSGbqtZphls+cmMVxranZe2AjzV11DRUZ0prcx0eV/Xm3N1MXqnFW3SC+9
oi3h2cEFi07insr94OKRtD4IzbyLKNVawndcig9GnN1e7XNXY2SxvfWgES/Y
4KKvwjVflTPDTgUnLhGA5qqZhkO9sYqYgLd68GYRLI/o+u2+ZJo=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
Wq2Vtq6aAehN8m9L0KRPF0ES9AUBVaIblfFoC9AhDZf7PbPl1qJPv3lsAQE8
iprXWpv5Yp0YUjKZWDtqT2qfFIr8r5lMIOgLF9n8+WgOrUdG9nPf52KcQ/1j
Njk6BTVJoApgyUjJ7LM3dOr+ejaCe7flcqbcXG6YoDN4cZwGOP9WotXC/lr4
GVP3Jpy8Bl6AlqNrceu6QCRWO020xM4tePnW/xvhQYeluPTnI4kQiFFR1M8k
j8aAF5GxzQE79CcC80vx6ComTemFJNksVXtgorOUjpHR3WbtsOJPpFWHIilX
7/hHk1JLy+YXkFxhMHlsGIzGO6n+mgeNGJznwtxMADdN6CaSwUlBCjdQnMD1
bwOteXQB7u+w2qXJisB+fPEZzbjQVO5yZTJnsIz2zjoz+Vrto0btJCdCB4AZ
3XmsOP6xQQqM5Is/E1KpejRpGIfCvKuO6ajjZTjWsLzsKkNiby2/UZjBJ/0M
MDzQEQG0VPeQQq7UpmUAyEPiafKWH6/N


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
Bp4jWM2YXRT+4ig+WSsZDyS4GGnnphliE0Ah9SEPLOjlolgaUFTEcNxzSpwS
EDfeAI1ywQ4t+5iVoo2fKKnHwjNYfpHc/fbI8KvRrqlpFCUUiwJfQ2DoAEfy
K9YuT4huQlzwMwNqMpRAHY53DOJi7OAK9GCBbMXbucfRw9Q0CGQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pRoV/Wmiklu3l30ydlr7evtmGchXCD1qQm2fN8m4xc5U/PpvhKPCBWOg7DVr
9R+bBY73B2vImHyCXxJiHe3Ls/Wbwb+11Hk1UuUkhmVeWaiVFE+2v+zvoiBt
jmmPQjS415eqWqAwaI6NcuTIfPsnAXSDNyaNBnyu9BCDoCmDqKI=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 82480)
`pragma protect data_block
d8tRN88835ZR5xOMtYIkbJnDlCo70gaEQPdLQB1Nloik76IEL7Da8Lemmy7Q
1+5/1YgK3b5aD/DHHo2k4EvxEYmVNMX9ZqIiMfBo4shCygVxoI7BBTM2wbJy
OmIIGIGHWc5R3ywTd/PY1Qw90oxhTdtE+H0ZY3PkT8D700FOfZxdhmbokgyX
Lo2+AYvZHtPkGgA8CVbhvmTAHZDdLap4tls+IfwFKVB0RhAk4RIceGQimXay
+7dOpkPjKg9QCHe3EHXKj2spHKU9eg8goxM6lN+lLIF6kFoqb+Q9KVoka6tC
UEe4YglbPMQEFzfE95IBSPjTIk7YF1tJR2J0mFTAQoExEAuFpcbmKNr8V1ox
fMdTq5to+xgPcOQLKnfYawRqlfEdLxBMvUUOm7d+xSGSI+jr0ejRxR913j7W
EMhGxx4yzYqmDB7ktpb5HUJHHIiU1nOOenXW5HRR13tON4gE7s6SLt6ebC6Y
Tao1J4cKl3nhVSE6H+XJ8D51IepjCfVwMhrcjmwis2TudZEf9YwW9bj4Yirg
+wDBFkC7iwbXqyKs3ElDlG51++6aoI9g+E9w21QmZowgLQPXAR2EtWotpfIO
uB6EGDZmOfYGSlqF+RsG6UNHetWBm3bDMHW7fNhxGfFf/nFjhi276/veaMa8
cP8ZolLkTnu/GYYJ3IJvwGREcw2dvJJLkZ01gb2IgWQaHYtbhaOKahl2q05t
0qeDwR2FYzJ9KmBmHaWb6CLKWTDSjTGMRF4WI5fS/zAesOG6ymy9svRuLWGg
d0YUmC+2xObAADBwTnr+PzT+sWhu+Bg/MZgwnGoU4PUXHtKjrX5WqV/9L9Nv
/ErDrqgg1k7DC3/P/+gVyfh1QOwzLhYyfwInEFKuejAQyimPS9KuOCp4odCP
10pnN5PVndoVUjBjOzTBtaHB3rHMhu/G0F99vsho0O35DgE1RUhHDuXhgxqv
8A2m/fm2d5qrsoLaj+accjKa3Rna4zMiVCMOMk/QseJk5DEhNE8MKfVYWow3
a8OxFgivDqkNrWv8ySVZHvVsbUjby4wtaWL6Imm/ZzmEe+NwJVMlw+XyTabq
L4MJSFa9kKgNkSjXcNtNGr8yxHTkziXWtX6N5g283UUh1pm4CThTJz3VHaX9
KLuK6LndixM1gxcOptsJ36GHV8aVWMDyGZpYy7QgwxUXcGtEpKZoQ4aAgRUp
jzkNsWDWYYMAli0yfxrkJv+O2slrQq3PUPQf7w1lb1aqm3jvmdV5+D6a6uZH
0H1raxcLVELQOVB+nNsqOyM5khYo9d+mVt7/hhsUsvEwz5nKdWSV+2QMYXhl
B+Va5LgCzKuz3dTC2l7G5Sxs8u/wIbkeePp6XYERfDyCI6MzMdVPqUOQPmux
NFkVrrl9hQc8QnaiJiVJ8+ZX3ko0JIFpgepaJMa7/UacX2kb8iIAPGE0lK28
Kir04cJJZHeMhNgIbX2YgZRBnY6rTHJZyvSkJOXZLv8QPAVOkNvljjxbHRLM
jEs3ZNWF7HezxMfdP55XD0QuMkJdu2RlDG2i4ZcDMjdtcWC5Y0qSm11xC/oi
EttB/W2J+y6XKQhQGYuG7fX57WAW4k4k07WHRk1d1DoLFIqQ65wJIf32eM+d
/WYLeEjw91DUtu5Z4cbKcjrS6Bre3UjWtguYPteya23ePHVQ9ecBpS5T1pgf
vYfyzwoMP1244qRLhQ/fcHSmrSrwNAgcCJ1LklRpolsXpn8/85PitZs2Wm7h
OjLcC7a/VqXIyVsZZ4aAXquMB494IF63luU8i1BMAx1wqJBMl5fAGRVDzOwH
M9tmFAUuEZ6H7etErfICt9xua4C7c7LrZ91vf1XxMtPNuyjSXLWoVlQF1V5P
j0iwVvE26TxX5bG/LvZ4JOS4NOV+xu0x7bf9sPiMy/knjXakGMx884z4E1JJ
yKo/gITjVnbxvrQ1LuGtYi5KxrKW1G6e6f+An2ld2bl54QbNC9GrIvkSmrlo
7UCncoI/rcfEFoz3hPg6f4on13fsCkbb9Nwgg1v8oQxPclTMZBRitZcKrSa8
tsmHS9HTtOAcMN256YhlSdqJ6k2z2pT6gA2JyD93KVQ1xg3Qe1MYWKZmAApH
ns03lWiruQsY7j69v15U0nNQzv7fE4aJUp6uY8XqaeH2jAAShz96sVkP+TOn
iW4w8noLBW2Z2ZLZTpKvvReLwC16AQTRdi9I5Wo7C/vrVS/kwlkTMkjqihUV
08oFeu5mcnw+/Tp3ffq35SbdURPWX0zXrSXDXqzxz473giXZdXrgBC+lGfn+
cSFfwBi95/Xyn9wfed5fK/9Mw0lRn0NULAKHogNgxbCCJS3C+l1i38bWoPud
0vXmfCdKAMcxVjufMijKPonfnO7weORTz1Px+HBCHGrfHgXYdMhA/nbnCCFT
BZM/kfAO7PWFy9Hzw+STMw8+hLXxTfE2vSukMKwgmyGJ5uueBQe7yauM9Hld
u5DkU0tNhmcEAwFxCzEM6Df1eVg5i8OZApfz09p+H7I7cOCNjmVl57PIDxl5
Jl34O3ZgIeW4pClo+mYB9Ni9M9e3Kp+EqlimLA8DML9uWnBXRAbtpJnRbEP3
lyVYCuziUpUd/RiyzZ/eNIIilO1HdXhKrXPxnxS5XgJ+pMN7a/yplAeNKNbE
MjExPPkDvnx9RH2neqXuaq8U2QxX6N4xKNMWJTCfam4ew5lfKDGidgTUN5pV
x1kj+WYay/pbadMBnjpdIIeRlavZxtHAlSKb1VvFNHtm6olWqNe4hxl9cRDp
PFHDmMoftw0AaqlYudFPYJooHPXNJdYq0yCP0RChUVgqVnr549n8DFlvdJSe
D2KhoGqPsujH8NhLX/dqH96gAZsuPCTWROswF/oO9VmR0EQHxr7LDXWGSJUA
Dw0uoPFGEt0U70JkiDJCCYq9YoyKPd5r940W1LcmgW7LQypnPEJ+pJlC5lUB
mtR4s9GohPd6/FgOhtTEmIbrVd6o5WVlGP6FKEnSbJYO1bnTCC29LN4CfGdC
G9cpwZgym4lhCTS4UCjtRr7VvLR3OOxFcxa3m8Qfr7XFaj6Kgj4ESAnLdqEu
SLb7DKRGwVyeCMhi7YpxO+TK0FPlrGYcAt/6tP1orQkSrGjPMLHPvhdV8bU3
NAnZpTX8w17UmTJcCCygFH0lARXF37QXT2n3G1ORAMl1a8IxBN72Rq2VhG6n
mhICdtlKSHi+Afb1EBLH0BUCXTcJNCHXdbFN7QbcWrMvYt0kDKZjbZU+eX/R
1EWsxXYIyYVGbp5JlMDYBqtlnBSd9VBUM9n6nfkJJDytH03NBEv5zktNX49y
ih5jRbScDKKp7N90Z/uAx0S7i4nkRGT+2auT+FYR1ndLlDAJ3wZzrMnft3AR
zHzzgmOJhJsnFzMl65hdLZb5HGMSnv/WvveJjF0ZIrqFmfsVtWUmWtIqYHuN
vW9V154KvRrz/fPrAvtY6GLp+TqswXLK0y3GcnFxPHuqbbtnezsLvvCpDShK
rQjuOJtNRtcmKevdObyqd2m7z5fix493IEqdpeKpJGHyZ2LbPtB+gnq0bRau
2rM0CosDDBVN62+LIOZQRbIO+B/TsByC6TBcRFV/dIKY6RtCvef6E7Jm07EL
7Pt0Wv8Mx8UQoa0pBg9qRPesYYifXk6YXZFl3Osmb+TDyXAdm5R/WtKbJOCr
qddlpnomInbWSe/+UT8/HIJIN+3oeeM1Zl6ukOuHRDVnUGm5TSj9it4CxpQu
iP4scbVCB3paKIQiRtj88fK6fk/HdwhEWynE+nMmrTu3t/XYjJCu2BrLr3iB
JIxTsdfCcjel+/HqCi4o/4FJeQLJMN1uJ6AlU1SSgPt4BVd7nbgJOzfz8zWu
1AgS9U/K7lcKoXL+fn3vdcwwiZA9ZkV/fH+3EGbLqnsDVWMMxsHy+HAy4leX
UxCvSxZingButc8DJoR06re77vdb3hnCv19rLT6+bsXzul8zhsZBh6DixDtk
FsHtLFo1XlkFnbwSI/IgyIXMBMgveJl8rJgHNUHn+vzpo/0cKkXjJ3+f5MHX
lWYwT2Y3C/h9ugUiR5hpHLo4XDR6s0OzNoOGPL0hCVdGS6MHm1OPRRPM+Rat
t7CdiD0R3wOIjnPcN26PPp0uy/sQvLeHknqARMau5kig7S3ZpJPjp7cQpRew
a+3jLxcAQuLAZPnlWrBmN0pxSaE6MvrZrknKlDnjmD1SVNuLdzSR5nTPewv6
X8MIRDWw58pZ6yXEr9eKD5pxDLcmk6HFrqeULN6+Ukt9vzFa1lJUfH/gpf9P
5TLIgZd3tEE1hbXIuGF8yprFyLp5IQzFvzTzeW9dEXwzfoX/WOEFdZbImTr4
nvIgPAGD3YwIO00jpgMO5mb+1BC6hvhpn+i9wiotqYGrzlKd7ejICmckby5I
9kFfBlZVB7BLawULYkjPMKPuKJyUTsqq8yTOXtInntqyV/8IEAx07rMK8ZSp
d7CVNUutAMEVbliS/+4EdzWEnY0HFP6Aq4rKZK+yY1mkdFjBlbPrG8KGVLv+
0ypufnI7sQIR2w8YM3oiC2m/h5kAqSSINA1hLY7cAiaUhnsbFv2n2MjpB4b+
7GQYdWCYlIR8vL1eZUahQKRfEw7FsLLrSPaxbRAuLTPuLIC3MUpTEQVV/Cpx
lZhcmgkH9cLdzUA0SMdtZLDpyB/IkLLZRO8PgwbO2QrhDohC78ZPnnTSWwQy
uRGptBZO27yViXhF2Ulv2tkYnMhvkbK4NNed72souCelvH9YwomhfMX+ul10
mpld9dFfj9bU8RbBrYFnJQ3uwUM3Mtj82l0Qyb4hN1zHl6DYBJIppvbAL4SZ
UkKKujT+dHrs8XwACN8qW3ejk/Bv+vHtbyYqBzKX9ObuG5l1AMDFqxjY48w4
SqN3y8gAWAK5USMM4QyCoLif20YuE7UfSYZOM3zzWYbnrLoRoSqc76jTK3uq
/Kc5du5amcCgW44/VLQtvNBHa1M6rQfnMmHooo8ljJUCEtRE4TZ15Ohi9M/F
hOm4T9sbpwtEdy6uPRDnsQxoZOoXepcTRPU8t7fUv5U8aR7Z4C1RfDPVi0Iw
6zLZSNFH2d7+yI3qPfW9EqyjFXun7hMd6Qwl8OVkMQMbDgMMvASNS6CWXNei
h7yolJQrgqrxlOVTIDbG+TxZ8TMJFf7h91hShKFBG6GET4TNj1pzWEQL7rq+
rELLTjvgRQ5DxAkOG06LzS6grp6tUehlnw12vT/STQfrVfVaK0uIXEyNNMYU
muGhvDNp6xG0hgLBIZn1DRYHMjqOFVjmeMUzf7fHQnj9er2jzBvRi3+hHZht
wx0AJCrV1s1vmoVmfR9SlP+iKD7fmsE+jtSIJDc5PZ8X3s+NFymBAbwaCTDx
4rHMN0XnfsG6qfBC9iCLhVBt84t8C8HFroqgmdaf5quQfZFalsww1mJP2wj+
63kxOz7XWBkLSCm4/5NsNn9CqXbtGCou1UyH8v3rmfCT687HdAnw/xT1/cYI
z8U+dlz9z9U/UIgeZ7esjZ+DxvfKu5lawljYpUvg/HUIyS+a6EDmJ6qwwd1K
8IzMiBuZGky0tHvaxTYljW8elkgIk9rqW806Tf69qbDorVenzGgPNdH//OJU
dH1uKqF0aGwNvCHoNnV1E1XLnAqOgVV/f4irjzYrllOy1AI2O/yEZQmaJ9/9
cvqxyr3WAvZZDuZ6wpcrh12lBPniVZTTBA3HcaBFck58/sbCNRq1OnA2BlB1
t6J/QZUD8vhQPB03oCTqd9xtJxG/R/4E1JosK0a+o98WvRi8FXIlD+awnM5A
E+0vUJTkkNrO+EgKbhWJeJ1LDAAZ+DMA4byyAylXOh2/XPCRD2xpkInozaV8
6ONp/b+eegwLmmXID52fu9LeZGjn9qmQuGJvP6SPFz52fxA/YxX53X07DkX8
SIAkiCFYMC18jVXlDMe4jSByssXrtssp5UCf2FjLTh/hE6Ge+u1k5muex8oc
tGxpDkWmCoiy0Hq7cuSvgMpgAKzOiv9Onx4/N36qahiq5E/zI4PLCOOM3ajB
dIG9LgBSPnz82lSD9bSY3u0oOutODSGbbSXtN9AGfOKuKezoK5kYqRValGHg
+3DQQNWc+armmA/7VjEdcTB0eAYhrNGScp48yY/+cxkKwSirswUg8I0VfbmQ
F/7NwKLDvegjRyV5fKJFJ/F2wSBXUfLgpbJKXW+m64pTwAwc84iUfNnZRDeF
SRbHiDBhQzWaOJtGd4kAYTO0kAs1dPIskamBaCuvF5ALgmLjNdG7C/NLr3SG
ZG818nDZhFg8QIiwX7Yki2KdUneeUBb42a5dJNWVCCh3UJe354CE18D8S4NI
TEpOzvteFj17NzbdyJFvvcfcO4U4OgYTsp2ubVASrYz3TVB/0sr1UfxVhNHR
Y350R54M5OpH+e7jsHdb27w21OQ9zArzxa0Oy3K9mibEgPx5faqYzKjLOMTx
gTVPd62j1H5g7WfQJ0QpaFqOnqWhBi3s8fHUi+bqmY416MX3DxKlI0Wxy4hz
MRjOJFYajoT20FbgB9OXCbmIfmMDH+BdeJz3W2ex6jxvBgjw34WJhKQIMknd
hVoVPA/Tt/f3lMET1+64hZo37ocaYtXKQLLE0Pru/MGpNYD/6G6O6VpeR9WL
tzZEb/Q/Gt5VYXPDFjcBm0m0csFm6o64GRed7sTK3TKcoNicDglx0xPL1ZQH
BoJ2ERkYncmng2VbTM/VeO9/ZBShKEWn7mDvEhseNFMlKAdtQaWOnjX/dSI+
UL0ZMk6Qwvrlb++lTPSd8j0M8dMCDXVeoQZmAR4JempP893rEBEYo9xs+tqL
i11tMaNDGUVdBx65DX3I+t3mNEWlpX3VOz2x8lnyPLEi64zLnHRyyFxjnXZm
sx3gtPeOXojp5ORleAq5+W1BDxATZL5O9yB1RUNDw9Psp8rBJc5641IS/yYD
YCzro0IKV0gZ2MdrJSMnY208LiT33j6nSwCDR6gLKnd3NYejPLLx7Y8eOetH
jutEKIqkfV6ICiCT8aXr5DhEkw7K1A01pdtcYRSgcjMO5kanr0EHf96Kd8q1
kwN80np+cFjLBeLYXzZ//X5zBM4xhK6OorUpk9kJrnXfz2wt3eaUyTACBFqb
Z3ilhH6PotGUGujMApXlEm/Qs+Y1sNiL7Gjgy/ZUAZJuzEDsdqmYjf9dlNHm
QdZJ6KiGbDu2Jt2B5FQbA3OPwfCX5uyG4e3zJrk5gLpdRJSOLccVyFzVz5U6
JBmx9lri1gvQbkO/y+bir5nwlZ2+YqHk5T3plcdi/0W5GytMYvEv+eZUM0VB
6n2U2CzEnSv3/zYMv+GT2oVByyISfqPtdIvCf4eizW8315UPxp+w+Pfubd5m
Db5BBztJpfVtMhPy9Shocipp5b/w9JDVVF2DzgCGBbag7uGQHJ6ZFlFYqfG8
UIaAxdt3QD7L3c59RNTZOiGwNOd5KeQpT9BEFw8/uDu7WbfYn4Hp0T8+c7po
BoAOIcM7sETOIW3c+vCtX31SrGj9FFZdY7dGXEXwos9jvfFagUtQUGK7c8I7
I2pMXaRlsd0FdT3a1PyaFBYiRmQGW87ZiOcxA3eRz07tXpYmaOVd2QaQoCJ4
JTZ4Ct9o2kOO8TsBAx+HAG+sqeuRLhm6hMGGWlzJyouzFN9r2QVVHX1eDD8Q
+ETxzH45CgqanURuFy8xX6GQchzwVW6DFI4Zd/j8M4uslBrlxO3yvvV43OtM
X3b2IbNwaaSah6LQChvGn5YhrhItSx5G41dPx8f1amDt09CSLlGOhyD/dcLn
pPy/oUDy16oh5F3IuiGfCHKl+mVsnCESg9APfNkq++NcQiLNY4rBJlTragsa
yHlcdi3sUXOgwz2aAL/F3e8eUXpuoNVn+ie6gkpoorj3Olm1I9Cm5NRcqDf/
xsFez/2pTvChTQuxIiHloyJb0HpG5kZOHKJlYmR27IYMW6kn/BLYC/pzVsNe
jrFDoSbHOn//swEcanySpp1VaEO54ZTOvnn0XJ6XQPle216qO/zgYhz6DaR3
PNes2tDDXeP2kavy//b7zfGcp8D064Fb044TgrKOyX2/dK36WKN+Z6B0jxwT
5N7r145CDbxO8WA7/5Y3RF0rpXqRCg/ILb58n2L45S8HbqiI5xMRBhZIUTAZ
BdUkRP3GLq32aZszUTRpNFuhmML7SHs/Y09N9eLI3zXdzxXQ6bMOHEIZKIsx
20lDec1nxAyMfuy1p25Lc6kF2RwjwdIbbiiDjRESauuJ/kV4L0pTqelgZG3P
Fn8GQyzR5zLKV07BmouONHprZQAHe97fQmFZ0OvSBJS5L1wdENxo4sFoU8nu
VqEjl9V+lGpj++5Px38Mtv1h5p9IhiQ9ZA9yKND5b9tlszOr0DmUvuvVtLl1
g/idDwmIt5KcBRN4sOFjsrrPsgcPPMHe7aqdqpvmk9rAex229IjoMGI6INWo
Mi2RJw4VdlzQQ7HgoAx5hCHLVxZU0yKOkgBmGZT7QXv7MAvpy3d54eX9LKJl
PUUURwYVVeHdWG8XrO/W4HJj4OShVi9u4WaZ/9c51g1Lhznt2G2NSvwVxqsM
YxXvBG5PC582ZmFFoKpJozhvPzVmc0OqGYEn7hXYGyJQ6q+Zijx0QvvdxoAV
I1u4VD+ItGPPIDjA0EJEtwsQlVLdli4BioyLA6kHETJpXLusEeT5kYg4Zeld
Bq6tGpJxNJAtWnDpFkk7SDSec8p7EAjBx5njHKUc6ZadrNaRE0Ddtw3HPb02
2XuzfIqCIa3XZJRR7MTCY5r2F4n3LoMk9pTCSRVf3YpZRRfmF7YoFmy+0Co/
LVHYCsoJdyj/PAaCJFxpbkP9iiSE3TxLasef379kzqJ7Kc/+ETCWm1z4pxmI
8aAneivOu1Jip5Ai0mKl8bvUKQ/nCL3mQh9uOVS5pV/HFUdrDfs5H6Sjae00
p1bkpLu9QmFSw/GmGuaSw5YhPWp/MAIPnnA3LaVPGyr7PRhWbTvhyLoOq1HK
DoxHKgAsD+CAbpQvU+z/jh/lWYV/s4+I6FJjx+V4ZrzJRxr+y9UkoV+oBZk+
LF0ba9V9FM1t6+JiBAh4fBkUy46wngJI/zNu3z7VE2MsaFKasyb7nB7Gh4ss
eJyRMOjkhpjtnosy1/9OT3iZNyS8RC0Uvf+iE9pI0sOr96oniupljYOp9e67
FqkD9JqQt5jyLul0HLmI/tmb7OGDWlbHbREwtBRomcndoKzFMdeIR1/bVYMc
F1znJDOXJvLVBIAVnAxs2u9lFkV5KT1fl5XGfQ4MBa/QWWvSfXTc5V5x5Kw2
9Oehnn4WtTLUqThg3RkfK9HQVyqbpXw2UwgfJBkrDxOCpEiEuVp5yZdjBUCo
e2AwR7UPBRtI89n9CFUzdYSaz9dFM2aJDfig3iwd/huCz3Y8C4OUPqNo76R0
a3FniAu7fM1nhGrxZfQ3nhNKrm0dndt5zZw9HOq1jw2KX8Kr4jgbTCgRNfng
tzZh2hDSNlrfTRUPO08AOdkoOTqBNoXDF58UMK9BzejqfzAj0DVOsrfMTxL/
nvEpP9wVQcAL4XuwozX++fOYR0IRuMz+l+Qqv8fr662nvFhFE4dFuH4KxtGA
lyibpD+JGTj5DDQsOSYPYPQzvuidyoID/vQVRF6MG2xXpRv74rSlRuXwGfl/
f2/PoHF1cH5S4XUX5AUQS/cgFu8XuZ09iSB2g8aBPG1Tz7jKrTAJNCvr4oQ0
bRIA+nB47Z2W/XciNC5bDfy1CKACwKK6rt6Ls+/T39jkjQkdZTgN2Z8lI/XC
LAkwmURWnfQPXJvbtljcw4Yb+EClQ8xHYvZZQ1Ry8Bvksbt0F/LRzODmY/rw
aW6p5+gR0viqpg13FPdZpcTt3/DKkhiTVf0ZoWgbQP/Ucpk2WFwjwVOrOkIw
8sinxROxpuvFU9DKGjADaN/oI8JLrYeLN+ZhV4D2+u33VLYbZt//xMCkLQ64
kptn9O4X9xlqcJdNdVV2pUjaVFEDObyUHxG3OS4dV/xbgED3esSNS+PM8ho/
Z4mWkCa2/GL5gkn0k+9nFx8mXQku2z9JqC+b6neAHVh2Mm57QMbuo89WJiQC
3wPrGEbXFn6hWUHZSQkquK0pH/59rJlsTl2GqoduAeIhJdqI/KU+lKSAvjFi
O9CBJ3rU/Z6M1yBgMK3TOAMp1R0dsX/bTw69bUXeYwALx5nZdgXCIRdYKTNR
gYNxF4H3h/picQp84cwkL2VWJbhDfqVLjSf57NpbFD/BXoPOAobgwL/UjBjc
qZbMb7y1l19LCHe4TKRAEjZs15O3kGMCGmm0fT+45ANts+R95aC3cFQkL7I4
kqDz2ZPsCaaBOpgeMV85xMH+gBHbUr40dCz5JzfoQpqLYELCS0P1cjc5vc5o
FA0+BEPWRkSV+SEvNUwTvi8X0xxMfQucufkb9uKmLpQJFHAxqBZAUpH0uOQ8
tHGSqf0QjAqJ4oulKAWsEw/wNzne+FZMbxEje4YU2KD6RZalHS2Vht7MlyaI
0dG6ORJ90709CzZZ6MeLdgA+zj/APggpv7t5TezCe6pCCb+mRiQEIGWvJFwC
9M9MitdZwkOwTjaNMPTab0DTNK1LuxjLQwv4IGrf9cJs9woC2bZRfgGsPkvq
tuuJYxKvBemVOAluLjFbTlRMblFM3KY/ugcGvMnczB2/TVXAnyKgI40fYXHb
0037vmvX8rEc8FO4/xrrsIrScIOTezj6FowzmeqGTz3NQioW/GOGknT5zVWZ
cPeLUDqNIxfS0kMf7BXSXT+BtJihlZpQFTBqSulKPLVXBw6HdTv8bKL888Qb
CfH6X73p7BPnYkEBuu4ror9DhJr0cxN+UnNgu7ju1NoZmJnEGBnB2DrjYgjz
xmu5GGLHnKjyELiMszCSBeQEM7Yyf6SpPeZri1fBOnUzCf7xHkl2jBPZrW2q
VYwAgpG36J0aR/jwaVVvWUv7TNLG9gxbjXNIsqpviOfiMJpvBJKf0O9Ir8MS
XGbB5Q1P2ENIqBamlhKhlS5dwagPvL906r4cwCR3GwWmHlrGruSEpkkg2cps
y8QMcfaKoBNjmHT+UpEBYser7wclQWMeNYjl3xzAlDJMFBwTCfcSaPWZEKkn
uc7p2P9eg6lhb4WTrwnu2EhqydhRH6WfoHoDRBD5sa5SQCzjIQbVeuIs2zvW
+VkHEiB3m8NX3x3KKio/m4LCrQJF6jS9FCnowvuHhnJH2us0GuLBBHuIHgMt
blILBDykbqanjVkdC7EWWHy7OL1CRihvMdIUSiU+qe16Q151430YxpZLYakF
9AwfQHi4c4nci91T1fcRsAniOYBoKYbOOUMlJA0GJlCymRnSL38Xsb5/NZXF
X0DBZi9mb2dlRLHdYhNVfvcwH8gpS7996sf5NpoBc7fqQ75do2TnQMwxncRd
J3xk9OTUO7wvD1bSsuse6xHU69Vvn9svlY+gz2ly8MJ0XC+JMwuPBDq5+LJF
KjNSjAiBUaODP5l59y7soGCtobHK6aLbKSfa7zdtlZlbrabZQWl7+WTsiG/P
0jKHKgJ0f43ipCIiaKWyl6vKX3y302DRXoTwhhmIZ2oKzJDCKF3MmNG6xRff
pIMUrRAmt8ive61YXL1eHpUErzp090plVvb3R7SD1eVGG74KDXRchiO1RqyA
12x/r+9vDWVXTcKMfJOGCku5n5D19pj8CMATVhe+6cx4XX4b22oCizlgg9rN
PHmCxpL+jCldddMgsD3He2MOygjRZHEo5iZYoPzhm4quEmjwUIoscKio6kIk
es1Ed42tyQofMVO7pCGBHOitqc2heOxq9zCAzMiJkQ1zM49kunscO3s3cji8
hJQ8AV2ztnhm/tAk6qqiT1+cZzxohyfnqfOuYWGLvp2nb6EvefyqmiTeWpzg
9A+KElwYMTHnnXDaeMGEPWtA+FCiNKaDqnLz6hpsXlqIygAYyDYXl+0OgZ7U
NnOErpQuQvOzCKoHE6xvZqSzRy8z6B/6j6sPdGeDfQpnYYzcQo66rYprltuS
xl2K8MmFticMsIW6gzS9mUun2yZUyPkQAu3qrIoNscY9YthRVMkmVvXLvdbo
uFHJbajj6s6y2mP48QDDvIiAAQCkoVHJKM3DWcyNwEn0zmdOOrRRojdRJIfz
n2d+ZieMkLPQaaB/66gnpQImL/Kx1wJHVVuniPmRVifmzqN75Qnq9th7X6Il
ZNqZUVjFmkCwBfXJfs252Vi3cDf2FWjSYrWXgfgwSBgAw8vCctnFHLy02u/y
iDjOY3dQw2JYS3ZrFx8Z5fc4OO9Z20Y1vQGhrlxwTW/Sr2ETh2TaCTYoc/xx
ToWmi51X/iDjK/NtA19yhKVgleQCpKEWcL8Cc9BrDxhFfR+GEemItrtJ1IUy
NyV/LCByKpHrj+1PnoKMV7xzUenB9iMvun4+fVXUdp45K3mYfoB7DKHAkzmQ
mYf9KDuhU/HKYm/Pva6h+bI1SadNd62HfKGH3eoQd4onf87shtOqYUlDgyvv
WUvkEVFaWUslCES0L4qSoO1tDdSmC8NXHrmveTt8+Ts726wnyVtbo5y9gV5R
VUbIK/bSacCCdB8TUWRfEaMwYjAAAKCS3oLxCgt0fbZ3oAVhUEgJ+NtHAtbd
Xfa4l+HiWRcMq836pLvPEJT21jmmpaog572CMSFL0IJvXmt8hUXWf6U3z1u8
RTSIGObZTwfOp71ZCp+ZysYmm2eLd2nfT29m5VdeVQcPBf7YeMCNBkBmwQuL
b+UIC7kIS9Td2/IbBvyOjxM+kL9ZmEcD8T32n6fClQDOITNAeTvh7aQBq0FG
8WbsdNeGVd8rM8kXQ1nUy6z8vOOiOgUgaNFKxTTeEnIs/PNaKz4Iq+XXq4ex
8GN4bI3Z6gRcZIbbB5dFAaR4vRZSZG2pfMOa5TQFdE/5n4FUPJQpm9KLEgcw
beziOWf19SbgE9+ibL04laAiUroEd0tepXpj6sIKVYR6fgc3CFJt7oUV66gi
ZSVZLsW0vCzYY52VzbE+VUATcK1boaOVqNfdsIu6BNsL/HBbX40xwNj39TpU
he8F56aD0LresboFZGlfNKPzmWQHqUCJ2jvYP3NXp4NjMlBP/+95NwOsej/v
JTOt9muTc81xxkpUSml+m6yMwkjOlOkhHOJjdge/5Pq5Q36idKkL2AE1jzEP
fiZkRFS9uAmmB4tgh0+sU98G9y1Cv8s9JGOKjsgY9bWW9MQokm1ZpqhYNTOP
4d8NdswiIfSJnbqa7LOX6/e1PPy4GuKdbxepC8QqcHiqoiVYJBhvYcJiBozh
X2ClFn3FqI1eEiSti9Akpbrv8Sr2soI7+kovAnlCf5siy7IveaEc8f6PkeL1
CeRZuhpuypntHt/5u1NsPhsokvXsW6llln6fC3jQ71tAB9DnhYwQZZl649HV
ZdM27k2ns0HXps1tZXb34bhq/YHKmmVrXugKQnU83YQ3mIOgkntKkrbEQHpR
2x91dIQBKUbpIHxw3KbcqzM/v+/aTpH7/paY1Z6AFisg7C0rqmAL/UaliL9g
mESGTmxnlQnpTzJpRvkwV8ambMEtRXfBVYZEP7bscBwulJtNYdELoNhbwdip
Fqaceya7iSSedKk7TtvTBdUQRSvJT4PX2lzRYnI3FnCnfawLpDM+kceaBh+b
7x83fR+fqVQrtDaLnVdFoQ+1C8ZcZBVm0swczxIRcccTcFTTg7+6eQLixVIJ
YDXO4feOcD8VnB+fgjqhoqLfFAY7JiztxQpjc+fUJN0C5N9LDznQMYk0GHQ+
vZWGR1St6klbWUanJchBJISJMyZ/eYng3Dd0FOuJadnM7vV5Q6ZIrXYXquYo
50s1ZQUl5Z9IH4aUDK6vVlSJV6dWZO7BQtocI4g2srIjj1BppvLsncoCg7yD
IQb7uOMESR5o+5hKqb4M3v5iKd852Zm1Jb8FTXzKSlYKry4fx9CyYCSwhK8Q
t3bhUfLYrm45VOZLyJG40Yqgso5QazKy0DP8PZDbPkbiy8ezJOF4lYb3OCxr
mJSCGwogYc99GzTEYD/2Q+dNSUcXCxmNErYN3of8l5U8ngF8tb/8XKQcNIqh
UF4rjC5SpWr17aFhM9mVCf9ENM2Bo7b4ks+ULUwpNl4nnCaxQ2cGPM/RSxs/
old/hPU5m3GeRmBM3W0XtKC4gaaLGcHqPiDTxT08WjWez4oz9RKzOavyfl+N
OW7vhaWmkA4azTeoU2X9tUbdJDkYSdLvMUFmBu+Nr6Po39cDbKadCQ+WgI3D
Khh+b7dQJbskRyjx68RS9Dd8GKaBtjhBrck4k/MpDwIvIz5xL/Rdp3rI/CIu
oCAzC7yRB0TJR5H0pG/cGlEL51F9uFFjf19Gt9nqg8x+gmHLWN34kyMW5Nhu
1IqONZjOb1yDHICJ9n7ZT59pxD9ZPtWWIZEO2YW1L81mjfDvM0YiCdtGTiRy
BZF8d0TSpSU3LFghkFjj6bNf/y2MrrDZt0JYAF5FUe4jLpzqrdJXvTnz6QXV
ufctIbVf74TizWKQjQIrPJUnXfgmWX+g9pyhfTrZFPIhFnQl6u5GmFrPpASm
fSczBPqJmRxOGcJojvRYGn0bsOpe/21xRZML6Y4OJOCpMcisDy8Zg14/cpgN
5HzzLFPac+6tUGd9vKxgjnQhy2yoQ7Quh2DfyFa4+/n7qV+EOoyVPHmWKm3O
VQCPSt9SqUegk3fa0ryOel0/o/jTtH3PyjCD7xmv0dMnA/6O8RNCKgxQN4No
AP48Z8lxaGZj3GpdnD3qlnULIkS/x9+1mQdS+X4jq4OnAZ9biEA0TBEURiMa
2WXzUMoS5h8luvyWB99IPcPbwhVIVbKj44HBy7rdTGjhXr3l4UKUBnInREIT
HdTektEpVvDZKVnozSgpAWrZomwvWQsU+B28bDxkPCBG1tVj0ILToUaUxBvp
wK8TilVODLJZHcDi2BBTiDWEg+qR6OLchFk3jrQcSyXgrx1ZRYcGfOEd/UNm
rUEqAzwHQ5h6K/x3O/FLHqLvWQ7x1QV9zBd30+6TPf4QLkwqZpRlL5NC3sPb
ohI5lACboS5OAFhjqR2mLOHirrE6P+SRMtbCC/FCz+nnq+Pn8MLZyBkzFle+
+Qem53cRWoWKz1XEXpJ0ZEchxr/l64PMtjA+YcGWFezID7Wo8oJqZSoQ345c
UisrO2l0RX1ESMZf2bieHqYiekguwRnx36lK9lQahsAY7MitTglF2iu86gAs
X5c4nAWCrKZfwaEleKFDhpFt0A7eGr+AbdcSJp7YkqNgFcxVmoVqYpTjcKjK
a0o9ajUKYpJWnCHPhbimvshR1o2fC8WaNILamjqAqig5zRssx8+geLGWx3Zo
qLb9EL0ZhvrSP774EkAAux4l4Pwc+CkiyaTi7aaqy/jVdRWwM73zPbBFmb39
FeeEYMK2VqnlljJfVyBxesxbI8cnm0+DH5XApaA6DPNSveLriV/uojhbyAlS
WE6jyzkkkmaWSasOj48H/KSjGfspSo5paRGygdHGKhzcRSOObYxetER9oPu5
7x5bNi/RNYfhCRAxC02yMZ320EtO6JIyVU4kUtQ7vS1I9ICzPa7nIWue+2Ck
GfcNk7INhUWA+4NnZRydCrh6QR9cRhNiFiYLcQftaS6yXiYl7LILr5QQWtfE
theQs4+TfIVloUxO9zoroCLIuK/aNHYPQa++265WtnSIoxZX+MPqV+oX69h0
g1Y+i4n+le7u5RzhS5jCicIw1BT3RDrMkE8h9rICsGz861XZQG/Q2DEjcv22
ZErfSKjvCddEPf3LmJDJ7vOv4N1PChMr4vNSW9sGcKEbhesHuZltyg4CYWNs
zQghYF77BIs+NhZbMR4dVJUK4ue+5rHGuzHbHhYfC40YKu3bCljiSexGMyLa
K+ZekSVfT8VYKNQWS4JTva30UcpMKh22gPyk4tzdyXdAK7RugB9V2CG8d/P8
+CAr+aUj05fRfrFKrIzr1yCnDiEOMsts+zXL6EU1eZaIURv9Dnz3C1J/ajFM
/oSNi8sNN77HvzmNRVvQfGIN/QYLxbnxI4TyipIXZyGhmtvZtHpE2YdiljJu
1Sp98PdnNbPRR5s2AmxhCVje6hC4qpwZRX4dJ+1JHEGGdbwKPTiXyjqo+Mvf
gWGzMloKO+XeFMN37Bzb3I5Z7YJrr7vvhX3UtLrXn+aCPw8FhvhNOGw7Bv3o
8H0mCCROr+OFKR0kOxurNPH6qvAYgT3gkdApU0h1I9Me8m2tnrXSV4eEeFqW
FHBBzh/9nCxdCRMTCNVX1m3m7Hd49DmmdQG+KpalBgGluIWGxd6dDQBXbH44
lJ0445JzOJyi2bDAlPPKPYkdTvOKfam9qisvYO0sa391Bpe7VYRSXunXcKJT
jo+kWhNJ/7BMQb88etXhlGBoAWhvOtl5xgw1bgpffFWHfk6y8vVL9M/N44eI
bput4DUHkupb6yBBp/ClUl00HOuVamfqIX//9xRB5NeTgZLo43D8c72uGKfu
DvBAyUC+itfFxQ8dWj48R7B4vx9GQnicOyeU7lpX5MBiXHASsou7V4h3tZ1X
dlXexktmWxu1ulrWSqhllpB8bjA0fyCTQHutTWLI8odb4HNe8fjVt8FEY/ha
mqkfQRj2JC5v3ahxAH+26aWidcuD3IFCs1l2CJU5cYq1v7VQwxFIo9fNUFgI
dc5nQRTCbMu5LlUKYrM1npFe4W7M9wDljb5jIal2I8+GYfAHwMu2CQvUnHge
XFbdezDrSaEarzANI0MOZH1/b5Zcw2euZNJPPq+vPgnnkutJ3Nahl6+Q1TNV
SzCevQacqj2x2sCGkopSlsD+kjAWrZIvm3J+Z0Xj+iAhqCBouMabN7BDrhL5
qtdoHVGpHooo9oXAGkyXiRTN8rrM0bqr2aIQ4PtKpHd6lvsQ/M6jAisgUXhO
WA4JzNGJ7vjwM32pMqz2aQ2xnI8qhuWlxWy+XpOq7smcRJwZt49ZZpayBG82
XeXwfVVep4AlIWJwVM+L7aI5nv3qEejR+bBsUoG/xqyEz/JxBu25vqj1pZKA
7Hr8KZJ+ulnqUVJMdKLOxXXsqe+CARu4m0jOZWOweGdhruq7HbzKMof3NdNa
kUQpXwxKZaB/yfht4KyAVDajD+Q5TshUn4ncOTmfnE6o6qWpvpj2MMS0FfyJ
rXyg5viiaRH+VGjWqz47a46lGV5VchxAjKSrwoloUDBGJvlm33NFlJpgHWNv
4eDSuenm9Fak2f7OSEs8gxLYs+T4lZwJyA2Nm83U1sWaWFgGNEpT52DjnJCI
nX41Hg20jdsdCjvogJnwq+BSLq9caI/k/iSy89eGVH9ojs77U5ExCDMEeAZJ
cxj2NGp4SbitAT50OGfksEauD36mRsOIeQCAY8nrW1gna7D6BM3LJo5enhtm
Y5EuzqQW/UGll3F0J/VLSJeRG90EtW4KnGSP1Ewuy8fC8OEzDc8SOcUKuRxG
Y7Pbtz7j1098WBc/iSE+9JkqT5TjtaG7N2IDLBSeKfV5sZzF8lIO+wfdn7fV
C6WqJY+dJPuZx0kVta6ywmZyWBLP7U/yBoXrwpNiggRUdJ1Sn05lRrjZY/49
OqFz46WY2bxY065i0NI3s5Lcbp6ixX5gqbsH8rbcAfI3u5QSSxkHC7+JTkK3
6XZRJynyWe8Z49idcvs/eUpXQvhKdCPKECpoPyup73qKr7avH3ctyCzYnrLV
Txy93oTUSx7WEjXnd6JAI2din2+QPiJDvr0SUnBI9h2siNvu7f2EgB3bEwnl
L+5vmhTG+PjcFpnXtLIAPeCpAtjhzUM5r+doWmE5mHoi0cFJPefZMOGfugV4
bx8owmhh+4iYpkt199GP5nX9lyiHDadtk2qNGLlcIKfYkTGu1am3RcArcq0y
q8vR8/Kw/kBmCuWnGEU1qAF5gHbrJm89aO6iWaS3S2VITzF/ln5STw3zaeM/
Kr4WDQQxGdNx/TlL0IfBr5NaDMiZTXHNzTjsY72gN/bqJJ032hIhgkaVFIZI
VHdv+fQag7cFzXG7Z3U6m9+So2tFLYjJ7dlPuaEaf4w00AQwqauobxzNMAKL
+9WpEHDcJ2PAVtsLnxXDXSEL7GEcSoweMCd/6dJO5taT3Miua3SLTFQ27MIe
jEGaIN8bAcghBUlbqaMLjYombd6cXfwzmSGhvy60vc+MW/vu6lBK7J4z+ly5
BUZY7Y/W2cJ1EfZMyexs2aB3k1KZmpoaQ8nPwO2F7nmmDPQFKEAw94Ne+QKJ
giqI31lFsNl4YnlBQ4p8Z1FTZs6drnwDxLkY7Wqtdn1GxTKM6gqh35+OcKZ3
DORqqZTQgmD9YZvPYzxKNbr+s4NLdYGSJI2c/PTuXResOpvqn2DkizJykXMi
rw0Nft3b4LkPvpOwC+rJKmwyzAZWG4OZD9jnmEpDB0L2I7JfBZZfQDqDgQAW
Ut2xcitNUzMMTblM5msGqimlZk+DWR9Grv7EHGAq4T0oyzE0oRKFZf1DdTFR
kKfv2A+hmxSIeEPfjal8wZcQ30SRGiPFxVtwOn28jIRtrIiGGzK5HBN0oLMw
LlYBz5IKQxqRe60acKd1fNmrVb/yHX4fpGTMjoz2mYexBgYM6Kj0nx4UzT24
TGYaFV8Iq0MsPz731vHGwtEziIHeiBwPGkF/02Xjy4BJXdeIacIa/RAjOKEg
CXo1HbMvy9e3/4824h5En9E5zv6nmTm9HZzmTXrWdXzQi+eIKaVHi98ckW3u
DSwKCTXJ1TW80x4kwL4PKaMpY2YmUWZCYdYNrwnrOMAzHNw6+HR00HUbCYmw
0QF2ueOhtW6DZx7HtjI2DNUGexQor+fM45CLSEmOgajluMPOWkEgYI6Ui3sB
DMIXjftsRTDpSsrI50NI+BeMuvGWC1HIxjvw27eU3A3yG/fRwWIRchK3Omop
0ZzmSYynKdWRDkMIiC/wl+0SN/lAOfhxUT/JWmf3095nzo6nrgCMaUUpqKXW
k1c2U2YfpkljAHe9hS6XwcanLQ0f7T0BaXuev7o9coiMt5AHELUDFgzywE4e
bJzYDrMAS5GkctM4J3rjGL0yndokTzSKU4lUvMl1NnylvTYBsRpgt7fMHHE9
v25KpCwuqIeHwVGByBkylQ5HX+MGnWcFNeC03ChQ3Tiu+g1fXzjN49Xfx9wx
W18QGALE2edbZS1ZYAq5B/qmLWV9CrKvT28EN+rY8Zu4y7YIuFuQMAsPi6sD
h3nMjv1oZHV4DG/pvdXiRSpftco0+MEFMlNPffWS6uDwsHuh3f6vdjsvXKx3
fiQP8KS3zMZr9+qD4uzbz5VuFlObGtIknGZJQRLd3Eck0NtWnOVRxa3Po39p
zcvx+7oQd5ZBLQZawebH8N/ps5BjLyxbl9EQTPteN24b2GbxaVetewNk4Npy
KC3yKtMPYZ3LsCnjGT2AegBdee0354VOMGuadOhKRD0BEXiYR2Qi+JDE9W2+
HukMVd0Q2/023lWLGR5EoY6XyL4V9ObdGk3lwC/D6BbORQuyaA2Ho0IgYAB7
/zW4LYI71DlvMDtK3teJIopwdgGObfKhyEHyNaJb3i5NXHGvzjm0PHhmmWBN
SpylyDPSpI2pnZ6b5vsNaZM9kWLMBAdi1Ps7qj+02lq6qtg3zfD+Rwjk8B1D
aONIeNJi/SeGE0FZNYW+A3eYMGjEfrKikq6hwJ7nb9xc2iTaA84uVRasvH8L
Yo+vgMbzhdcj9Eme7OJ24MdIes5SJt4YkMAwbZzwJMgBTF4tLolwryV4SR1c
MzP7/NlTxQccJUwn89Tb4MUydxHtAKzuDko8iYTPEavem5NZukmlAQC1b1kd
oQcx7c3ZuraQ2rqKbBqx7JwLw0biXakZtOpvDNUYxcjxVbdonn/Lq+WKZDjk
KrgeyC0K+1aw82Bx8P6nKd4876pT1x/J8raW8fVcycPVZ6gBKo3qADBiRZXM
0wBM2tb2BFFryvgvOV753n8NHljG/tNA7wQFhgXiD//ufe/L8gX8CdgO1h1J
ahnHKrwwMZGZD/kOUhZrz6VGEtZo8q6I4oEoJuCwgLGCWXhqVSIoN3oYUK/d
wD6QM5y2KXI/eU/S7DdZeXGWWxjF+cg/wwCncXlfscEmUnER8g9Zy957tMjm
bYo8nIquQvNG7dFHcbWibI3z55LyuOplJJc18uhxL8Y0sKMIFQmyrO6H+Lcf
0R+a1e5d1FVPwNyEbmlDbMVH+3JSig14IsJNf2zA5ixVJF7LR5B0erFWXTz6
xT2nUN4Fj6Ym3vYtm8P9h6YzaDAvHWupv9D80SVc/mBPiNZy1m4+57bGA3Je
UcfZOYlLcRvLadYYkuO/KubI9Appunb8Zwf+tFu/dhAJ6N8w/ijyHIccJnJs
s7wpbwJHRMgzI1QViBpZwfaqXRm/z7IOkuNxTHTxV/azt8CYRvJvvT31RsKs
0leJAsC/Rrx3c/4yEVnDSxzcDOxbqjOaJdVnY5N+qdOYxNa43zy/5aPa5g+A
xisl4ZzIF8/0Nqj+fyRv7qLVPj3wYihIfDXfWLraDk56yO0kST1j/qBlWAqg
SdsinfpntaxlR4e7y4o97cQ45OqzblNaUTZUDb3e3BLLDhBkJnKrD+H0pVAw
xYWZRfyk4uYS1A4UeS5nVGlYYk04bGTVyMb2PKnzZLD1UtxBF7GkHMshUB9t
HMXjnEKA1Aw6p28vxn2N8DgBG7wtPVjv8a+u+tLssZQJMGWf1nYqzf5fNFdR
81tv4HkBYvThCGxFVGhZqIjPcxtIoRffFw3Y7aDqHkm2Wj2Dd3tk42X9oRZ/
B5DuhsgX0K9eOSD0FbHi28A3Bd2rF9n6r115Q8kQfzRDYr25trTyMWW9fKVF
S1T2NimPqP1t8R7iUvN5v0HKk+y2lb8mNBqzMC1sP7dM4Dxd19aRqjSSIZM/
ty9tan0C7lURMJprXf7Ox4D/bQjn3g1R0QR3joSBLBNPNAWMg2aTro12hoiJ
rCiB6/k4lFc+e+EQxeeflFGHDFPyRhvrxR5L0t0OBQgTeflGbi2fKDgvTe21
9Zf1iP0lVdgvFFZHNU03m5/1Kr+x86zdbvjmUkMieWz+VzLq5Fc/yrsZd0aI
WUjwcfvgS3ENQm8n/j97zRfffgO+UDwhxZ6wdnBhOYpjZE0apSC3331igqof
fgkEwCntAS+7aXbsaz6ez+qZA9L3iaXux7sBjNVDrA6Z6BFAJcMeQcbRb2Ws
pvJV97JU67uNXrlJlvLHDRTr3aIXS86dwHj9f65cGHPvbwLDJNOIXAwaBYp5
XUKdhdmp25h4Xp73UjPt4DrCjDh1yLMZrGJPdQwXdL4XjLurf+J13elFoF3Z
yaOKF2rc8K4tHgKoIV9YSsBQoKQ0THFc1pFwuTp0jgAn6z8pJy4XHxW3yA7D
yfntwvmJA/p6TeXKtlEF2V6qRTHSQPcijdZ+marGjzQm4mEqmN+q7hYPTYG6
s/ZOe4LDvJ5u+a2lRfUm1CBbyV6pltaIRttQTsrj52yMqBe+vk6Ipk/brG8U
atgluZ2BScrt4i21hqN6hpy3WezCm4w5y3ZXzt//dlaF7o9+06NAeXnhIoAU
kmqjDUwdiNSysM3B6eDnSDprc/h2D8zJ/Uhak62x1jPg+0LWnYW29L8rOKGp
LvAZsbVdNvh+EerG/zGx8y/26PIRRiFsz6mytHAvYYpIqVZxdW0pKKDy3yQX
hpkOXWyriyJyO8wJqlrsKrL2cQN1NJjSuGYTOoRimPNTqDOrV6YHIgLf+O81
c9VZ5vB8ObnGD0VqvHxClqrWNVWKWjd/ZNnFwR90CTmgOpVoXlX/uDA9qelk
YYLhOlT4Pmn9UNurfWT0pxnNzeTQx1hxOZwywZqpMr+DcgtVLfHqVyALhdSg
ZWsm9qnuC5iAQtQIHuyLee6c4i2Re445OaRvBozHM77OBjJ8slA7Q1XB4ALc
1ygJZDzVZ4OnJ7Hpb7mv1L7sytNhZ9vmj1Eati64YLKGhXrcBTsz7Fi7IAUb
O6PbgjRnYfnJ1tZ2W+wmlbUv4xsFVawE5ZGTDxBL98RwxmGPBRgH6eLHHs4P
xMNDaZfMRwQITyQhEwv0nABKNxuQiJxMfuMYscpG1EWyjy7UP2YtiRhk16Yh
zbCVmDpTnxoaF2udQLE+B/LpDYhGgAVakLFM7SlUGWB4pZDEuT+bftXpALcN
Zu7O5udn0Uu3AJCH0RDKLb1mTgYgs25ELZpUWJRVEExB9gJKAXc9UW9j+QW8
dQ+iOu57hezkkzOGPo+d7A2Yp/p+yxQo3FTjgTDHxXlYncbLXfUk4TTA7zTZ
r/NMAZwhfOpv3VAgsTi/dCidVgWGNPW0cp98W2DIKYe7FKWP+1XcFUzK2QdJ
CrHK0G7VxpvBRror14MmWNRIjwaYKJ5CwcBZSVyIiI0sEc+IxS8wz450B4O1
HaH1GgJSihTyJ363v7Adw3qSmIKyc4a4bXOGI+bxqXREWU3qotoJTaAmL5Ym
SIvTMPCEKra4w3xbiLU7IHe4sh6otL519rvBDbuANrVzFkH8aqQXv4EcbgEk
zz44iSr0Ekmye7tQBhVCLZkdSPplUaYKU+5Mb+YU7pc/O+Qhd+ca+coUFNpm
CuH7Ms+1hF1amElK+ZUBjkIIE74OFaOkfQvub6ImtIBSEiOseXsUNW1Gqhai
6dBRm23MItszm4crVvbCNKg1VDqrKiLsS0BTzlz0pobjvV1cOm+rVpnURjG4
ed/Mwevo0dfXFYj2YTbPeqYN7fgnOTlY0xjLZFN90CV41hXKAsVtzj55BUb9
0OZd7mQWyXE6/TQVNs9Uoq5Qd06X5xeu9fFBBa2rs2D3svIw5l72KPbVfJw2
JaxipmSW2xkqXrSaxadyjXNh+7ELrju8I8koXHSipbiZJk+7fYIKe9FdopM5
mLN1AeI1zoTnoptgf2FNppQukfVjwikvxw2wefbLxwYWAgLlro6RrrKpR4b1
q/EK+B4N078xS4B4d+gi+70Nm+r4QHyZSupkCHpLBGy+B1DpDuU3bei+FqZk
R0PHMY2XNe1/nv/oNvttfsTkfwt+ew3EPtHVkg4HBQX78klZRBdwLnKGEM+6
ZT/E1RUM5tR3lTL0JrsxlmaI8M6sqJkmhL8Yn3FX1iBhQoCzsZEach8GZjS1
RJ8yofAKfjThvTTepnRbUVgHz7v8OurA072K7HzwKDfNqZOv8pdsMQ7FG+FH
tOyz+TCMjTmxv5mAlsbd7CnpIZiZOaCNBTc6BwVWEFJV9u5v5yKaKdqt5aEs
VU5IkvOnTSeuqa7F6Q2hG39/oEa2YV9vGkeAZ5cuiCt6DZhzb/aGeqJaysqw
L+XBtDsk3sZkdm5/Lg9Gxdg6llxrq7HqRboo1i6xYz60ww5Ss5toKb4sBJM/
Xt3ddszZ2YPU3C8nT+DwY6EWjB5TUETuBdy59Ekre6aTU3sjX0HK/BjGxB0A
Ldb5bdH0lYOEkxI3w8dlmySyxbFiWtByJPAGm3p+4cyzPC6ezQ3UtJhMmeib
PH8m1LRYhQHoI59S6QLBL6pA2tO18ix6xj+joW65945lEMWUZY1FxevGgiCz
2MSonj+kw3lDPL+NSimPdss/1+zXA5wh6M/iFeCcD3kn4MxmUQMXd0FV9FI6
cHYrBCC9kFyI5LIh8shBp1S7LmRmx4RbcHs2+VPrXJuYQTS26tCeKWrtmJjV
ZhjoYKtBCtYUhrpiJsAdenmJD9zg4Mg6V4kKEXoruvy0zQtQsPxtlb4RPaj2
OQkb1KKfGbtcIdEKSjZ2DYs04d6sX8bSgdHmiAiCiFgifHaujP9lWemUonG5
3WxVic2R09dRENllzQ7lyV7bI9H9OM+iLgweOYtMjMvcxGCV6YXjsLPpv2vp
NESWsA8+YIU/vyt1GjOZZWUjG/jEvCXRsj1upB6kTOcZCa6UBkpfbNbj60k+
lOMOQ8jCl5qdZwRZTuoC6zKVH//i0u+1HyDradcVNYv8+UQErinjUesGteOA
vRCmu7wXri6vDpehSSrv7+DGaCViBiBZ1k9/C2rHKaTAsAdjJvn4S/q5491J
/VMhfdRWkx3TO7KXArit9j0Ums7RIIWD0BN/BMCEO5vdF0UK8XQ635LY7OhP
8IJgq+STFoel21p2pN5eH8mrV+BvBLzsIbHGfLEADI6zJpR58kdgmXGP9LeK
9X1zg2ui4Fu/Z8JL3gtfBV4tLlFhAPY5KTCEJTBL4qSNHhQWoJJT5ss+1CKe
RpoECdXHwiodANbz/ryW/OJy3Cv4yv2hjdoHP/onxwFWfoTysraqbJFwO/Qc
5cRozz5DbzeN2A87D8do8+qbwRbESpPWNeUEfyeJLIeEZaw/P16vcAIILAE4
RDGIbjtjKkpJutZbiGzalczSbWprzdn+WGcYjkdWixYQwxv8V0ibhyHWR+hq
kqN7fLOjVZOVMmHBFemwBngfHb4UtOj00jywW1wohbffcO5IShBw8jTt9ffT
WuiKAdT+HUXpnHI8HAKFS37BsgJhodBv0svDcioDTs+9Qk/8b9MkLthURdmc
8eaRVle4fqFo+zHZgvZVrgjKFEidwBi7a7VW8qNZZC7/8bHbX6LbUF2dz7vt
LxGwFW2GbJLeqKNDYzNToYC6jEf6rEShNUv9+zpqqf9tfFTuex/0Bis7aU9h
EwrQBjPeaqmRDkurZZ0WWff6xKYyT7vmpMGsv8WqC3zQZvKnyA3QbU5NqexK
qa4iMVF+EocdTU761HDZgXqRJxCGUQbFTnPVurO4sK7PEI9fjZfPcUOmTeGq
nBJ8ZHN5yExcD5hWBq+LDCidZHHBN2pRj02/UsBeNoMFh2+AOzoofPQN4QWO
kJk2zVh1Mn7koaBJnWmYp0OiQ/+VskzIKyZk4zH7E6ky8XyiI2ZLsV/AK2lh
MetTDj9SB8SwqqC3ZzWRXSO4uJYVOR1EaI0bhQASyWFv+C8nAf6xelCmKVZg
gz45jpxp6D1qTj03s/wn2wT/O4XQIVADoUIAjx8pKvMqssdY1gi84b6+OghN
8F0bOVVeBFfqVApQq0c1lnbeZ6gF+h6cRiRDcFeEQ3kEkAdUxEWf6pQdQLwI
+rypyuesxHLwmmo5lRy5PeMHJFp8Ru9AOBic15NMP63+P7e4RjyTzwkpBShz
x1Wq/x6Po/cgIy0YKis4Q/AkTr2mzSLyBmqnODGOHHZvGIHCZB+sCPtGQEgC
N1Ypt1YFBhba6mOrOtCJ82y6SSzBA2pLXG5L+w21c4v5ljF4U3Ob+CPnC51E
71CguVV8BbIGU/6jtjJeR6vFDrVzhMurnK6nzP87lDapnJHe9Ilga65ElcvF
PNLYSoX4kTGww6eznxGEyM6l64yQspuSFw5l2Zv8YmwAiCKpas6tkLcfcv8y
W1ILoWN1jg+5NeMbU3mSMMi4NibriqhoWbcG/4qjTkQkfqzPJWrdsqvISfLX
zu74QrJm1M9MvtUtDt6vLcd22oo0PF+wJkzjTltZN83p2HDEIeROT8pPgfVd
MXsTJJvlGDExxbCpnOUovf9XFin84qyjBhU9VqYM0YFxP440pX1SLV3aV+pA
XZDoqhIiQ3GMkQNKgjmVHLJd7JI/yL9XLHwf1Jor7Io9V4Sv1BtLc5S0esG9
8g8b5h1i4p812V7EB5/lHcjbLZRZEeT/wy0iPHD7pp+tJf5MBsA+SqFELgDx
DJ4bfKXRTlwuXNz6it9c8ZsZ+dt5ELGMAabml4Jbes86Zm/QKLowEKbjLmIf
rD5v2S697nCtmaQzJIwCnzilQwe3lKVUdnwX66cRBPsVI7rsLsr64uRtw1np
Gjig4iOrFsE0ShOK1Rp+1R1Fi9h54JD6SO1I/lCw7dUDn7DJEdK1UcIeoDex
PjFaAPVGTMXv9rNDN3Wrvwyo0sujLOw7rCMeyHwrx75/+DIE++X9GJhWQhfn
Sjc+L2BROYoQdT8XEcCjEhVjPsDjpt9k5HFojI+Yv7jD1c8aSHM9TW2FpC6f
1X8JCTV2MRlQZRJi47y/FrOwXtvIHa4jJrl1JJFq16VTzFnjJKhB0P/RYEYf
DQ1XImGgDZS2pbLxeVEpMK2A73FTJ8rSJINjk1buxo/r036WolmDBfhMBiLv
XDzuIRk/kPnz0rlVCAZpmZZsf3U+mnrfo3uo/h+yCTyCnagPUj2BYqp1wa48
lCd5XYeMJDogREUKpWwapkvwTAWdWy9P1TPIi/mBxmZPJLbNe2030WOmKt3p
/AkCsXWLPlJjXaMmaRURBF9TZFxwShb5oFUk7fn9+0YyFp2c7vBQss4xmtG0
lBWo0Lhrc8Atjuf018VRulWpfHHU9fUkNDQi9ZyBT1FslV7w/s8cef1vNh37
HKU9MUgTwtURcclqJ7416xEAzMUId7gtEQGc7uPmSh7wBYSuWJTtJaeA6PC0
nWE4ijpzzlFGchDV/37n3+KMx9J0mTIbbioviA4L4lhO9zxwWtgJaIh9dYY0
W7M8AYBGLov8uMAqJXiD0M4nUELpxA/fuIXA0flUUwYJ5nil84HzqBqIglf5
07IeCJ9Kpynh3GQM8cyFLxoHBW1Q4uGTnAhJVEaYkBEYZb9penz08vsufo76
b/CEHZZktb0YhD/xEWkNWJM3Var4ttGUp/d8TvUIDfll5PdQUBQ4wA/DQPmA
+DO97BTDGo+QJmbudVBBCpo/UWExC3gOGsr2zzEC2g1izVjvsUkGVP1IOTPW
NBho9KBe0NpejArSzY4hITZmHESjbF896jgDeNljilgef0WAIwf29uLqaQ0M
SqVFkUpJ4Yw0cBoLEn9xjOkWjJQlcd5mpaFloeW73JLDZk7ltnxnVMkGaoSR
LC7kRz/Bl0I2wTYy5kv0HLwaa35AwZ/xf+hwdx90n8J8e8EQUbTcTmGvtR+O
bD+8SJ1qNMiA+ywRHBouMf5tkAdbDcerTmT++1NWDwwU0yoZnBXsQnXz91oc
yovmHIDj8FRhnMtAHWtQjq1/B9iSMwXdju2wnpyP3k6vXnkY1x5TZvHa2+db
yA9w0Un/Iv1N/wR5+WOLF6ezUgmRew1dF1iD+zcgjnwo1YjKhQFbungIiqay
zji4tVIxklORn2FB/GTPOwviFupvS9LE0+9EgjHkXj++XZRA8Y0kw2wZ6t4H
S2xbXSDoH+3Hwmgx1l0Iog2lAkclxo91Y4qX+bmitYnqWCXaOKa1fNn49zFE
p96FSTEJrjQqxh+5eUltLsLI73+UXEtMa0f4bIiGscE28YrYMySLEuk3Eo7W
KrYe20uBdlYI6JQUpPjHC3IyNVI+BianQEc3HXqUal4uG18e2QBWnllbcsRf
tXI9r+l09kcRJ65JWMSXjdFNwehJuH8G5uSpxBGA8oPQ4Dxt80a0ZGllkKRB
76kvn5+O5kvCp4X4hamUpsoWjfHqR2TJyYolUemehuojYmvGEHef2RXdfYnv
Xe7BKSnKidcH+1PbxfUXECxwEvKLoxga4NoPVobznf73Vz2g7O5+U9k1CPGl
dIv21JuiIqp4x7SOJdqjoLiCU5hR0DkXc3aWNbymFPJKlTZX2jbyQtXr1w+6
vQFXNjLvGIOhn8vDo18U/hp1LbTCCg02KzZ40NGSiTdhdF3Umwq7zjis55HU
XvHVqKagRsvnuymgGWHfxQRd9aRFcaReCsNak9rVFt2WfOOZS+Y+OIaD2rnC
/B5hdZxH9BjYgAe59xR0KWdcX+IRirYu5gKq2/DzU8Z6k6hIKcLKpXWQRqsN
3Mkzo8CHWYXpoMMuorp9w/oWyEf22jA2S/pfhGu470GDJCXIKRYrqBAIrAYl
AddhNvTcgAFn5gDRSX7ak7uu/3tWZjoKvZC6aOiTDckC+lorwhi5+U/Eb7tN
XA8/vFQc2uCGysmc7IbtiPrsVa6vkogpI1/oCL80J3IAimkXQtM1ytJ39ILo
evdSYmtUtWm2a2waXMPVH5QmeSQMDoD/9JBVQjj6vCu+7bsvtI/TzmDSSBPB
Oti0QHGLZJEX/2ivnTe40nrqPCQktLu/nybkfAa7ivY8krmsLy/1T10IB/Ej
Sy8A4iJG9Y6l6wxisQ3/uAXJAveycv6WBejpvHr9Et9GLU21a2clmdRLqcsL
/0llQfHUBJP+haLq5nMtX/0fAMd8W8iCJji07i0+RqKEVgMZtPACF6BgLun9
Fna0UBaVxgwmIDSu6mGR7j2KxLCNiLKBoWlP6+RuY+tHmVz2vdE1m6PYZT1a
UVbhG8mROo9I9hHi2VsmuRgl/EuIWBtH/jSixSB80rWiwO1dTkjJauQ2sPZV
vN/dFlvq6i37bdfNdEAjVSFlWuqDUMBDjjL1v/zbCNqWUwCgneu7EYYxIrmr
M13nJSOfzqLPWdkxOaSciTl0h6qCdAerchoFVMN9VbFTOAr2o1p5RB9dhERD
9aMCNP/7tmBsAejA/SSVqqCBukhHzPdDyGrlYfglah5WQut3O/TRiHeJhZaz
NUV44kbOTcLKhmWgd5zjQJYCr5i/dIGSap9XxXKxDlhkCxrpYWf/TbBRFYGO
4VBAfOb7iBsJJP7z/ogKOtY/6FZMnhePkdKNh2BKoPIkjn5ftsbfsoAnuMzx
gIjjGkW6myFNZCqsy6jqFnWX/FcrFMUmzzmUVNosuVYUG6Jkb0+hAUtZCONl
ePbUzq7/Bwmm5OOUy0fAg6omUpA2cxkJSk2L/ckEaC0yslKnn4mWA4jxLNIn
TmzXsNLgYFJVDs6rv7gYJdtg5gRDJICnZBBNNMKeYxcf05b8ezwK3ZtvnGb5
ZcLRpgOW/sOz+24BWP3UTTJE1+x+l1NYO1AVrpdOGr2uRWoACTuCgmVWrk4n
HYWCEIjpN45ne3T6zJDEiTvhIhTLlJIbRFAu2J/0oCQwyrbowSzhE+d3zF2D
vHjwBH3J9/SfqMo1ze7TzYYahvxRhj+eHEvARfcybzyhpo6DF84t71RCSu+v
eMFnbt+RX1MmmCE1GPqD3AqfDL5tnIaan9Kg8n0HsGsAXl0B4yIR3p8FyENK
d/JJRc+/ByGLQaSPglgxutc7kANd7bW1iGLFmE99UG/fRfV43EwD+oPb1R/r
Am1TxTi8wZf2f9xd9GnX+yzL+0MfF3QXZUWEQ+G3tAP2I3YsXKaVP2KfeNxT
Wj7YmiTDzdBdCEiY27/pZcjUsE+3JcYO6jzA90jUWav95b2EJGrTbo1oGY9n
bHvuhlVmsUkzqy5NQjx/n2JBxNIPls/MNnkPKOLnyjFEgQY4kqa1UYIzVMzg
z1uSbeNOfhFoNSYguLj2lKdwzdy7nHL/hN2ANjt+0p7cCHrtm5c7kqajsDIn
w1k9c+ocpMyVZg/pIElf5RIv4OqoLifvLM0O7KoxQUhWWO5hfvVzlfodWR2P
t4DAOxSNbGI+1VgLGu5GssyFfqXgdTGCFEU/SPEq/lgVoLzKjEBzxm+AzmVJ
HjUEfb72py3pfai7dfBgaVaXBQm7JDDsYmHPXs9KVYMQObzy1RtcyJIojDqZ
3bk+uxlU+RQ/vGc9hZz1OL5IGEXHRe3nf9fz4KrZBdlh+oG3v3OyeF25S6wE
/QX1t7Y5gqJrPYfW3YKPSEB03Du6X24JDv4bQAVE3xlSl42fZi6ZNDlrt546
RIgJ2UUQQDeNuzTyo6SimUpGdFO0nCrDzDoJk1KyKb6DvdJJJb3q8vLM2ArT
gQwMnBwNjoHs/A613xD+PSQ2KF8KDf+d9Ol+kO8MSULV6EvSBOHBy535qZd6
VDC5N1oLzmG3AixygTNIfqdgfJzYvOwf3t7hOPI8nLSHtzuXXNp/JAC1yspj
3kJrA5F5EXkHjcIRwqs1kJpMOlt0RTpemjK/DTmspctU+hg499tl0tY5jhhs
m1ITS72Z1maY/sMWdEWUrEHHd5wXZqYy0AX9SAnFhNsZdMCaRy26lR1N0Szz
DjCmcVyxrav+uIZYDfK/nrlkihAvS7Fyum/mPjuOmyCembN5JwqjrfuTd6Q9
ACEzbUV5p73nXzf6AfqjAkQaG4MdVS89kxclQMvprldgjSgiWB1oEcs4VfGI
EQTDMcF7GYhs1wukPEATEz6na0xAUoaSojJidgTYrD+8hXskRhos5HFSEHD0
0iWjMnPYKoj/n49D63vVeRSClSxFyeM4RkAhn1Hj60I848WyUqyuDANgD8CZ
mKb/LsOwtcxdnNPZ5mL7iY1ya7NizuKdrARcclNUpMbn3RifMQb0NJ0Wu6lw
jSymuHY4uNt/4SZq5dMIihVRvpU6Mj2wVKqkXeHMCIRW2ET2t9/vnCeX0Ee4
fxJRDdg6S5ImQS6bQ2XhajhskSOcSoxx1iMGF1OnJKPgsy4CKsFAcwRya/8z
HbzaaBGXFQDDNloLvKpFvAfFKoU7mGnRNZsUPJGTLrMk6wZQn4Lm7ty/0eGG
ts43Tych7DYdawprQjbqyQVGvDS4eV96BCyBADFa53cOGzrkWq2KdgItt6ZX
LGo7g5XewJvqdDVmstn0VJjKh04EeJmJTJLuMDKjwLfIfLbjE8sQN2vtS6DV
UahahOsRnI4xmwnT4wlgtqA2oLtNbNCd5rX0bAADh4x0a669mWe0EPfo+VmD
kNrgS6AB/uR/Z5liViYbEi0iikYOrxsoIB3ChoF/Y3fOaaWnt0ApTjTztmYA
kyldhMw62vRj+0icKEPO9gpJfsaz+ueqzR4zS35+G4t62R6Xq2QLlKLmmJLL
twl8wb9LSUdPW8i0eUQQlxTdGKkLpNc0qq6QN2ZcbC4vtQyMj0IJ0w8SQwln
+WdjG6VB0TGyx0CrUGwtSHFo4Wl+1KQmUzSqvPTCbBQQBHKYPHT3B16fN9ma
gSLfcMwHb2GHRWw4V6ZyeSJl27M810W55hdntpiwYp1gR81n1sDPAtV5qKtE
eyu/dAIW9V1Nno9yFN02jZmn0D6UUwe5ulHTC8b3JCWDvKeyi4S/0LE4ZM/q
5Mc2AphJ6KRFrwisDmQHSOpNoP7EK2RyrdSK5m4TPCo6O1DYzjtP+Seq0Xk8
XnjPbaZ8N5tMO/HwrQCtIarQpjZI824MvZotnau7HnWERlbkcpVd30O2iH0y
4kucnesUFyqsmcDI6JdOkFD14m1NND5JD4ZXk4g4l+XHXidfIL5Gu1YfHMqI
PrCbKluNu7xKC2931wQkCOpUaMq6byTwjyEjzFOQgBqVo4hRofvzI8tGugjy
lz15gJbsdG8BwkGk3GtwTYarjI9Vp4iPbYoPws2XZb3XZG5Elowataj6lCp5
UThL/frhnfswk1zvhYafoJhDHfM7EZQ+tQ2Q2JvBjbPQZmR5ZKD6Qa1vp95h
4DJzfhuhYQLBj11dV1WKg/XnbBAjy0710Hl5MQLAVXAoslyh+VJ8A0Q7kBtw
oiOUY/6oCd9HF7RQm9RedtnmtXNCGjQSSP/r9KODzDYXZQ2WoAfVjixc+nda
ADu4kl1uW0tn6DhYE4SENwPpiNYf5LVoveNcJdjWd+h5Q7KutrXekZOwG2qt
SMGGuBxaKVYAhnTh+e/WNIXn1RJdHsPVnvN2pPiJClIdCOoeg6fIDIaZQct/
e15v1rnzKandGoloodtFFPtA65lJ+GDUjqAJafqYF5p4sc77YrrTRP3tRpdc
2L8xfp6tWJS1OPKCtMhnUrFh4pBsmO2X1KbMJIdvyHCnzLcdaWHw1Eo1m1hZ
cKEh4ZqNdHEQ43QNrGRj8ZLHU/tFE8qgnV6rE6XFNzlKbTw0myqRgg5F4mjU
Mgs8UPhgVzCvsyGphyOkEnFiKvJUp9rIzR2qNrlR9EqwSbjszBe9irVbu9Kz
3kUoc0lLcBXJRhxApr0inO8xEZsuPCMkzpwAtQAmALWW7X5S3ZheYwvwLLRS
+fJt8jPCT5H/UcWLgvVL3UVSdbJri14Y9sYZxdg6ilIjWunf8v82rHHbDbKL
WMx9BLJqt+xXYIgbRkeLfT3RWe/ky0bmPbFLqpwQdDQ044EYpiJLRVDm7tA+
olgQXCRIZpz2/o83uI8hCt0N09A3Ew7GIrr+jyedCIdx7tV2dNHDpZiE+1tf
eAh5CsBLkOWDNkS6RlaYNfwnrSwlL/kEjIFP8/JCkR8ITT2GkzM9bHcI5P9U
+TEaF7XDxPlTs+lAXgOec7rC25Vv/W2tRcoh979J5dQCMTv/yNcBtEQfL8aA
5Z3w1g50PCDjM7OEdJq7KV9IdLlhxpSDHt8cGUS6tM4l30R17LXd/kZ/YUEg
vCqzFeXwhS8HL1GkJNBXRyZIW2YUYpiZumSkMd0CzWB5qQ4gCMJ7VVOP6B6O
qqzEtV89MmCIkJaBZ4XWQMU+0I4gZ5QCzYlGpfEGZtVivAyzAPdJSf/uaK+y
ybIc65MTYsPEP1V//MKRz49LeV1up5z8dsssYzXej8odv/onh78J9PmET409
gaLyZrjIBsduUSbNHo05qjxo/AL6f3BtNxKqwKHr7kpx83SCjaE2Fodm8etd
YRCs6LTN8X//jgLmygAe6mTObJsib0OovQCv4HfLSd13tOjTmnpzGioNGADw
iGjKhdB84EdCX796MS4pnYCoz+/7VMWBa2kJvIVYOsjOovyYGVyGL3Vt9X+B
M8u+stzJea3U+yLVJncB1WvV4BhnLl5UXmJbVe/sEapIvJmoiFYeTZc6uBRm
JqxDMb2LfkFKEXyh3XSnDlYTpVeUXQpuZZt+KP1ds/mYrPF+BAVOCJzyDHWD
IQ60b2AQGFrcRiQE7CgPvnngvisWqRFLPEZjCM9e5isnfjYKg5Eky8yOjRb7
pY+sQIc4VsJy077v7/iAH9at0RG9KxnmGEZnz/YZTVYfO7OCz5OBaPoKRYcD
4lecdNFi8VKlxvCj01wrmEwY5XOZ3ydPAQHozUkONO6plt4QgUbGdTRaNiCm
usmJhEO/xk4oGR0tUKmCOt5Od/iI/6wYWnmw+vcKnQydk6Fyj/5wizWTPf6p
ZGBb3s/eQ34dRDNmHMnAc9hdNXJKED7hqvz/TL708a50LVT0RnpN5mrJVsia
o0t2Z8gIMiSzU53B+INjFPDEByuynkoM37xtf4bnbhjIlfcPLVvqeOsY5c+f
iFJ8Phrsrw8BkjIR5kgUD0II4gl8KwoGKaieJVeNLt2Ty1EauiO4WOiLmf+y
llOR4APrg3uecnEo4+3Xargm7Yjdlrl90AtfNIkMuSprhX2NmshXwx2j3W79
vZ0xMTKiNu/N7RSy3k5vsPq5sszr7ZCN3L4HZYLHwks/GuOrZcqv5UW5pbUR
Ac5c/RVjBbbpsWtYLv5occkBN0ecA/0vtHNcxdMLTW5Qldaf4j6CXzjYQsdb
+LoTY4upT+6hGw7FVZsEjLJaK0z0AOYgGOmtgu8RAl2j+p/TesUfiefsk4DV
xnVDhYnDfcB0VPexwqQ21kn0+XRTbxmwOXCaK5EhpGwQl0Ou2GuVFweYj2ne
C/zGXk1TEn6DcDg+TCMjkTP3y4sR9VNlyYZlNT/h6gcEsYgbjN5VbzTgbDdV
r8nPFCG897AXvYxT3SXBtR065Blew8bXijSGmRzQ3doZmIvzJUqSX5ON8AhS
NN8AV4SFr9SfqPl92kWCf5cKIVQgiwhl8M4p8fhkNG0+REn0LrZbZfT1sM8j
3a97HaPa9B7owli+4vOJfXlq2NG5uxrJj5p0Acy9o8+TO4uK64zYO95Yyl4t
FJMrdFxlp9GYVjKTyD4UjE/46Gckom1iN2ghFtJjGVs441bB5JmMVzF7Pajb
t1gvPe+/w250eUiUHl6iF7e0mx87+S+bAf6rc/lQPOAV7Qt1E4YzVggvfpFg
FMVyEedfnKnUWpgVrl9JAHH1NXRgtwkVvgcc/UtmcBxhSFJT4SCcGBWBwVc9
y9hD35ark/SFmbHlQiQ+7J4BFd6ha+Ks0DEHe4DkC2PIxkDdM3hkrOZ+5OYD
2m5+rHTs2XQjQSvEqz9eMlIDGoTl++KJXsC1kX6Ihb6syArX+NfJEgTD6WsZ
tcXmz8qhYymo6ekdYP87zdGeUkmfZ2zUrVc747ofsJoNs4A7lsXnMZi/DbTE
ndMWAq5SaJmXjFYcLVfbPZnxNkFm2kVne3vdOzJNxt8tMjNG+UbQEA4a3U+6
at6gzNZABbobiRPCSVXwHAjpZdFw1e6CXhojASR1jjHmqzeXO6UeMQsui+n+
2Fsr4zlQsUK6mKWE/plPtrDaIw8e7uYmhWjJwbXKWCKININAOWWGClTR02rV
HSiQTU61DbDOTDvO6R3rWC5+jWgAfvliAJ11OQkmPuHV9PZ0cyRtHNdl7xkL
z5UnRupGQM4lij+KyLSUbROKb7M1eiL1sScCzauOaxyDGY89XkMKSF2brPHk
cO7q3WDiAzIhE84PPOgfB8Xhpg3OFStCaLvtY5YOi4vKsYBz+M6YOuon0uUM
R2gWWkhEtmePAL2Zkj19cUQ3glCy8EUhtnR92RaEYlwg/uVgZNjkw1g905VP
fqyyeKpAMDHgFMh79hzbugbKgzGo/myq5wDNEZPXtyk69SjYRIpKwD7QvxBb
y1q8qucL/JsTEuhFtgm82F9VXrQLqKXQz/ApGMBJ6+6iUmcftIG3hE5iiq3k
quApvOE151FgDofAHcAes5757x4Sh0jDFI+6uE4t3FSmdyqrTv5N7EbYcRLv
CcLBIPZfVeUzHI/PsAY1/tiW3jsHAgc+y6jlsbhkLruz2+Yo9B9buXpDMX8x
sPmZMQSJCZE2+BZjNFaWbmqsXWNRxryGzOID1adOeQCoLv22VLY5IrlowPEc
Y2pe1Kju4I6bi2zk1rUK4tVBnBih++nJ2XYYx7ntc23aXiH9cTgbmnTuKg4a
pr2NATRiFOpbT7K2f5qupxyVodrVW8UN/KToqb6YA9ZS5d6FQEPpXg2spbJR
rS9bwjPmAO/cvZuklzpVZcXqgkvlawXOZdQARv2vZpraMgwIfTzR15/DQKIO
PvHNlZvo4D8VEPjxpNunagQ3lU/p+2WGK/INdwzQ+p4S6JfZPl27gaailGUK
t6OtpujrpPcLC/n1iqjN0UidTWG8e+qh2YKQZP+ls80V75MaDJ7oiKoSmfT9
FD/Pinpe8eYet+3IT4uTnE9qzSjjS6Rk+ktiUGWEf3J0Jd3clYuXf4pFs9yk
VvvBroUeh6OD8hffBy9feo+F2nAEW37eAm/84i+P98MB31OJyfU8uR8sdv3f
BSi9MjvUrtzeLzgNyPWu47sN+Zi9eeAhWgnK5KNA0ezs7IC0/hcPKBJHRnwl
sLXsowp+5nNMKgDI/Dm7yOkrUJxNd4NWWnTpeXXuglTJ1rGJsCrk/6OdqpeX
gAyLNJrR3NoZIHS2ePeFIebywCHd2ebBnHWy0CEk61KPbVzVyd35ZhLmFNv6
DXd1grFGNGDpHwzwLwD+BcxbFxwWkjUmKOYTLZ+DIW9LM5DiVEoOpJenV91u
Z4CdnEMmnLKUVD7K3XlDB2/MMCJ9TMe+8fS/46suOrEHZSafooC0X5crWx2q
c6xgYRbbvcsGxxLlDNF00llV6sT981Gs2cyAgPEQAZ3eulZ1CF115ek4KYjc
pn0D+ZMnSHUIZDYlZ6jYnvpSS7p6I3gBhRgIE2KSAUTjhAG9j39LLnWtCGTs
Fzw0xjhAehu8eac1mzmp7V7IZR+Gt4gNppWDvGUXNgQtyDThB54Q4zFF3LQ6
IcZIDkdlePsY5aL3i6jgox5DeQXSB1JjhSJRM228rh4xkU9+bDnLrOW1saaF
rZLhqyS5ASbBDR6J/RFBmkGak1QIiZlzyntLU6bCSmfmfGjPJv3F2QZb+0Ik
pafP8vQXPEo18hpk43lVUIbMH7qI2lFzx2DJYu4sQmhcs23o6R64XMynWtzT
I29Ws1UMzwQFogAM+pK1DEShgIu9hAuNa21ehGJP6breN8QdtJoRgTD0Oc9r
b7BWed1c6K6DcrUE463PbFPpQn/+4qXhE7Ang63HNHAQfpLVeP7qrb4pJpCz
CProew/xkkqrCYRFIyxop5WFAmtoSkM7H9Hl6wiKjMf5Mti0nvuwXx+7zoKx
WuGHeXvCJFLvFygXsRMlOApvx7vW3mo6M/77qUzz1QUXmOBaRO/rkvoyhUqh
dWsNVX95pok7t3YD8PWhCJbzF1qlwPcB488gx8krCuh6feLMN310lDivO3xg
QSPDBH7kS57Jq/LVjHLeUO4oDfAm974G6aVtqd1EXE0uUarsAVBnVi/wjVrg
lUnuZoPzgCCyYNOCxloyry5te6oU4fNIq1gYOhZ1A0a9Wf/ryrsY/EbquTBf
HADjdBQl4KoW/yXF7pSeQcIvFSvguc/i/AvG+E98iGyzQ+xlg4kSF+sfvGuU
jhVA3Ehki6l0PsBeNas1Oq5jGb7/OhnpFE9NUZ9JiWMc1Mc0WB7hqiaKHn/G
JdsJA9kQJtiuLk5JW4+SHyeL7GQAOnPFVrepWJn+JauPGEWIHgqWh1iRgxS/
PU/JnocgYuIEvVgWbtI5c2IIWoQFe+L682+V2fSL4X9QNjjVgrNfmICQbOnx
v+/O/EhxlrrhC7+bwWSKi0sqdlg6c5WIwEvwGspdTUPLFrhLM8EE2hTlcceM
3zzH1NKSTyf4vDQFfOgAPPv/HZ6NULgqeS7RC8gHU1oS/7eMrvTgtMVlz6XW
TatHuuFe08IyooCWh2Z6XJ/gYXVNCKUtxRvYCv9oYxRPG90goejcvlT9dyJa
WUtN/2aG9ZfnsU/uXNjXRcAwHii8OrySQzFD19cGiQ4mCJPHvUHYzKTcShJo
AfKp1kbKH43V4Z8hu6jBJrWH6exR1cTsvo4fB+uJ1GQbb8xdudRhzMq+7uzI
UxVpS2j9nkMi4WMsGAMrs6lMMO1BVyVbfOKEgW8kr/yvIkDi3gLURXc2bc5X
Kslgud0tu1HqDborh/jgCwXRcc7nmvLahp2BjndJ00qXbrZRwmhKvYYluHhV
jSkVGy6GEDbIZNeEhGfbRKDUiclr5JlrkRguHah3yd06MBFx8wxqQWjUoouT
seSPjLrroNySvgmzJXtr+NJ4ShiyAixllb676u09gZHQBEVLZOj5Zvg3LfKr
paaYTMFfxvPc42r39mHoOPZDlvyHtKefyw+LsfNVxdncDNEG80nxpxuKI0N8
vL4SeAxtshNE3R1OJTI7YM732zyfZV4zEx0bv3YX/8Qfy1C/mFAv5rdOV82b
3It1NvPEkvuKWCFIvoHqX0FesKUj2VNWi61Dl5NbjrgQDoCssjF0+CYW09t2
pUwGLoZsYBS+HR7AzrpI1zbTKyQJHqdbDXlVu5tIWtp9GzYXrgu+63tRUDNx
2RJ8caafMR5qhB3XRD0Yk1QNBhUTBvJXidW/2lV+Y9KAieMtpMQzjy1427oi
gR8DTURJCOQugaRpeaRYe4F4a6HO84P8KPfpV3AMLwim5soy+BsGQfayQZvH
jIILUMlBOJHUJboZgozZs5ZAkdq5nt6XGI8W8FkUMySncemQFj3GrWhtjM2k
0fNhVjhB/5ZXmsYn35QoqdEk9XdVv2+NcTZ6J2CBmy29YjRoV9hFnkJ5C59d
b8q8qLGnayLohLhSSPqYJUT0lQFke2HonxOI1KSrPJZVjDFiyN/I5J4dY+3O
5m2Xi5R8OwzPiz3sWPC83gPTgHLiqgYJGs6Cw/rmVkacRFbfjufmtciaeQY9
c2j1K2pGi7XqmiBmS94jOucjms2oWNk5Mf7OA0L0f1K5Z620NhPqLy2tmXi8
lrK5i8mkN94Pu98JxUMDlEqexedeLnl9x4Y9thCFENupM1gNCznYZXTTMAuM
bqHypGSXx+scCMH5rZqcFCJjOJAhn/0xurttFwcN3WVrGZ/q3mqKyK4KHPqI
WiRYQpYmmTEHU2Yui46OfaR/swLVugUNw8iTpoVlooNa09Sd2oTxy9vJwf4E
jMpp6ORM7IFoHY0d7pr7JmKpBDIn2n7f8UcbC21N85kXkLjsVmLBjQfpB80e
ZvKnOsxAV/lsvs6SQNStIuTQ0cm49M4JTOet+Ezby8vH5r8hI3K4bBQjV1SK
NbhBpVu3Z0i/3nRq5znQLmKSCvmmgpFBpvzib1N56HkDanqN73mZbX5vnuFW
dcxiOTBacjRYhFFGvVol4/d9wHj5IDrn4KSXTd9fvhr+X1Xr+kpj3Bwdjsi3
7R2/GB2FzXfsyRz+ipCscyGUOTCl04H+7NYO0NiukAQYPq2b155O6l6wYcNV
hhfo2DcyZf3hHyMxVy0N03yhysQy5tjFYDPwvQ63PpymUOY/aidrrSCjjAUF
DfAaCc9ti0zmpVbs9Gx7ZTu0k202hRhvl6ANFwfOnWZgmNx4y9MSClh/R6/S
UM6oYvTpsTAPDs+cHonsZGxSXoZPU6dLi+ReWe8twxeBfcPO5Qt/MiQXd1Jz
uQjva0T0TFYjpu8n/VMmYM0i9WVJPUrBd6Vz5D9umoeu1wy9U+53YAkWewpk
ppa+Iy3LccGhj+8wMsOyQL5K15ifyWmVR27SByAfpfx5akA9iaIWsRBT47hw
iY1uxmIyhboiJsV6mAsNzVtAidzlaxVnKect0E/wzELcT4b1khhMZ0MKKVWT
U7hKV0FB1FG7+ukSqzZkHJZdAdjO3ud7GLcOv2FEhRaZl4PE3k7mtNt5DFYX
/XkMvPHTtn3plntlK2G4PlZ9eUIjwubjdmso0GUj3zfbWJyFCJ0rMQaPGeVY
JBLN3j6ozxlUpteycIPbAU07dsDPN2y5UU/hg7vy0AGO7eDnvZXhIn+1hsmO
KcG+y2sMhz/o+gNxcgdq9VZGEmT12xDjn/j65hMB2LtknVYoBilV90FUdFuu
/YekxDfoZE2MRXPa3B0BkxE+77GTkrry8MSYfWE0aEDlHWby7lQDDFp/EWnQ
kMtSB0A3+a3JpgxgxawO1clKVnf6zDwljM3LnuDqcVl4DDMcjOTK/T22PlLj
UzoFC3KJvwDN30Xao0SYK8F+0VCan9wAApXBURqmjwR5u7bWWhYHoozgV4f7
2ZJIDDdFQ5b1od7dW5qeirHTpDZCoVLxw7wo24i+2JjmsfBJ3xEEQLtgkFp4
iZwnByOCx6Na9Txz45i/3UejetzdlFX4sPKMuIQAQKuEsgayTSe/fu3iDZ6R
NA/uN0xJs1rMmJZIUajybN2HIXhZGW9vOnAao47JqP+FPGJngUwQp+oGEKBQ
2Jc+vBrMBPZdHvX8lWtoTy0ocVmv+AZ0Xu9WvwBNE1oZqATEXaA2pfpJeKCB
JzUL+Q/TLSffDM7KZ5IMZWOwE4UOxxtvCGlUrLaK43+mnhZVdEPJGyf4fr++
ZqPPr4BfApEfbt3cJiIwrlOxTK8oqP0MxV+KZre2OqWKm1SPIPhli2nno+Ln
5wU7fgSh6QwWpRSIWDcO4GE7gw+V6pOKLaEXKEkbAWdYtJTHFu48jYeuKq3p
ouCCh9XSbunV5dUreQlFEy+YyzjTcytb+wNSSr4K9KetpLP7BLQ56JQ0fJWa
oyo2/Q53iyZB89niMa88lZNItHuQXIzMRW8M7OxPZlAFeYBlzp20fg646/TZ
p2YAZVDmuAiRNutokSyUujSzOOSCTV/nvs2S0d4oAfiE7tXqBRNXRszhNTfv
4rdTTT8SfcKtionllcAlNTfBCJlU5weeMElYyZcEOqeiQ95Ex91UDoz+QN2X
/FiUWv7UlAwpaSRZii/2zjGaOCpyH3z1b+wuXOh5GYN88gzJcScLvKhyNv6D
PH9KzbU14IFGSJ2y2WAYS17L9Ty8edqsvSGciJCLGu7gtIyWX8NbPpRs4y9z
6fEDZBQ1TW7zLUqv/yf87pPbHFXAXU/RsTcrdb37W0BnEXJnl+RwSDh0X+/W
b6o2mgCVZ65Zy+zMvuSKR/6Q7NUg+KZseERqFzgFlHW30k3F7BMbEZhbLO/6
4KSXYKBBWHlGsm0laOVTKUzXHQNpzEFw3ElN5th0FAGZcfYw/o6t/mijtBvp
VkoLd682QOlMgZ71Qmg7KzExaxfmEXNAtqD6g4h2COWM91NbfMIsDkLFZ0K8
N3wIKgGJnFfSPubiaosMBnkvN5CvcpQD+p54McvgVFSx3Mg8cbiFhYCx0nk1
/TkYx3ZFh2y70T2wof3O7p0N3+ovSr83nVzPkcro9tDCSQHA+ga8i9ktmHMy
bKYTyp4luJN1kByT8UDXKdE4xNo21NelHGFmG5Btz9YUiFl+3OWBFhO8au/2
NhrCguVdoBab+OoYAMF+wDwZhjFtOnTJvHDoaVfvt0M/tHMylFAg8OOU7jNH
keO3hVppx9fl4oUdhUa/vm8KSdFKwxBiyZsywDluTVCjrr8mExoKjLmfMjuf
vEC7CAefze/W+c4X/Ay+PhDeH9MztMmQP1UV6SsosfPoVblf8Bkbn284MFM7
Nj1uDA4jSyZhW0AbNqSvUFjqVzkqUE1pkHDmPKzdgq7uEbSpA9SJOzhpJFWd
ejSfJ07ai5Rl2dsBrdMYsJxOqX2rmYx/jsQGHyEq8zDn60paFdfziv1ljEaK
U/02/Y7Ytutvxi8yFqDE72qcD4Nwx4m2hLeY2qV8KYemRr2QDHEvmEEQDjJn
/xGDci2xvGNOSyGWkfknN5cwmEmq3EqR7QdT9w0WLJ+Z5tKYfBEaWo23Qdyf
sXuqWvdSdZ05mKYtH7FAxR+gz04fufwTGTE02cl1u4ZAeTrbqj93Tq8jpAio
UfZqgjS/Uyj23umn9ufGnF6OSU8mUR1673PxR8bHTKc9s6LtVq7X0x4InDty
th7pZy4X5NciGyhvY+vuRY461XSWRejCj+7o9rpqCWQYbgGqo8yx1aDradeE
gSk5ctOPwN3k/+jVnShaGDDJw3lExar+w4vYRmwFytCfcOQJy6gdKXAkkoJb
FaZQsYRNCS8DlN5RJuj/0GGAWPl/E1r0KeUQUP6K0MKLgjZ2cRZSMeswWRLL
San65J3Ap2bS5I6pSsvB1B/6dmKAKVmHWPO/qIO2nuYUDloFMsZQApU7TIBE
F2DjOvYOXgRPwbeZ8MjDQf1sTudtfEC1+/GPXRDE/OFdCedX5VWe9yo6707G
byoAMpFYxZRtjvg0Y9yw53ynG+D4RS7vLonoHav4YH1iYpEjo4OWWIeASHKs
IRpAfN9gGuFoWKxuHcD1RHKxR6QtrJu/AdKeE1n7GARhEON9FCx1zW86Orhk
lWu2xuCc/thu/9SufennA+sEjA/A9NlS7ogo+PH6dGRfD9CuWF6dW6yooy3z
DWSyw1GQZnMUA3lfk9iTYQMS0M1tP/JNS4YcQAvuWrkx1e3K/p0MgxN66Z+M
7rg2Mi1JBFgtnthbFc6Fhhcdz4t5gS4U/ILiaq2WMVxx5F51i5i5MpK7BlMX
xhEB0Bj4N6iwQDKy38+lienq/QueeveaRwjP+p9OO1EO7wXS4DFlrDlkG8jo
aQOFDHuNGdIMtAdflXUVmqakF77WgcRA9Rwx/NCGJAZwBvS07bfBOuEZ+al7
rF9IZP//3hUaLhI54jye+OfAe6osajoxG7zM8vhkkwEv7DKX48/hO2gD/M4f
GiCQMLD/ZprknlS2JiI3mAjwQJ/2Q+la8wC7IolR2nqJoOSVc1m8wynkzq5P
ICtBDlzKwaTSxarEfcjPJk9EDfd6kTTanKD48CldR0d14375cJHwQ2/uVnvD
XrxNrMCi5KFJHr5t2hiolmWRaxsabfNCvTW6fBIwNIaJmjmkvHEfwTJZwJeI
CGmx3IUlCUNgkFsmw+LPnPlbnPQdpnPCRwhkvltnnzXMmDurA+dax1HMqRGT
J0OwdktCPCDknyPyc2JrYSyrXqx5habbn2rmf4Tztgt/x1BLnsjBzP21TBNG
zZy5Zyz8+7J0dYS1YwbT8QRRC1WBDwaDOngzzBwgUfm7raejX9PNm1xxYe+k
QzJOfqQXiHi2ERs2LQp9uRUj5jx2ehqrIyXffmyAzIXbFMGm9j8NlUQmtlRF
wQfNcu8NQpM4krw+vInI4JxOhI40GZD/izQVcwMGrtciowAekAxKyzmAV30S
OmqECkILxVUjhTF9JFzIzIo8UeQdGRzEk5jPRmjAx9jBXgNQNKvXsheQsCDf
3F3ZxM4/NvbPWgUGW0wR0HqngDJzHMXEFHOXItz5Mx9b5gkt1b88BDngHrTR
32GdtowY6I+lVKvcciHwIzLlsGemBoz/w2SVAkUREMaRp1OmJjk8ZdU3DuEo
UB7PlLn/noSQUNteHevYza5JXSIIX6wRw55W5I3106FS2st7+0MTD5FrTKXX
T8p4kDKfwe742uswrjgZgY+vbeBlnmJocEb8WWolW+j2/1VmFJFtnokU14ZM
Gh3EntwmUHkte/025JsDCgI+PgKn8Vkejb17HYBrItfzr0R868juWJZFQ7cx
hl7E5tMF6G16qtoTi4iJbp/FTY9xsh24FgpnrvWb7CZAANJrFiyYvkNrNG84
GFXov4oJ7yUu/Kv6ekl93ISEy2p61MZ03Z7tfNFPl7fSnN+BcxdEwldM466F
NdIc/FsS2145AEj+55gZKHT0eTCM9L6XttCpKl4L38ZglrIe7KB3H0JIQzYy
p8mTJ26rf8vIPDOcpQNDChX3oM2h/eb6y4TBNbwyyC8pecON/AfYhWqUkYiO
5Qw/K9MYBXG7t3P+ZUqjsBkvZ5TpgrCWdUkdybSuhEbNxwnAwV329pVY02JL
l6vMJvSR0eK6CEMRb/IEhneE1wMhZ3jRiojL5vEpAnTa1rOsSgvMNsdsOd5l
8QZVRkkGsXRrnTIvbUx7KmMiRjxW7f5g7ZWT3gaYXH1slI/UZWieFNqhZzKq
DPw5cmqj9Cj8MrS2MhMju2zP/UWwxTqvZqulEf9m4MNNaPHdEyvhpZ/EwyXY
HjrDLW2UdQ67/O6De46scuhEi7WF5Vi3LllDnmhTMxkfAphgGUzWH5A7MEpN
Ift9wlzT28CXZDjNQ4O18U9zdhU4yRLJF+ZqYdCjY5G9s/opxr/hIDRoWoDP
ET751W8LPry1qU0uvJEt4RBKbpKXlwqzOcYRULhEHVnKBn3yC/xLea/iins0
UmE6OZq2+3meIsIE1sXrbgPZXSu97BKkAxYJy9hDBLASBbk5GbhZqPZzAVlv
IUTUIA2yfE3WWcopVAyT9wC2GOZwQpLFSzbJqu9Vu4ZwT9QJxGOipFjPeJL2
0R9Uq/OsBbp65zoWI7sv9cDnrs1QAyX+NGxqg1twIU1VnbkFufUXpU66J6hY
c1aqwupM+TEn4YC+ZvGVSfTHixd7kE5BW6GXJFggY66phQymgS00K8acvDEF
chGaXHJL5pTCdp3ZOBRmRMnozphkbgeF5rsVJ48/Suss/uImZlrWAkgSuzba
75ix+ezafnLsInBEfSCbQDX8tzYQLBVvx7PzkATxswNZFOKLPERW0Lu6MPl4
NHTz9Zl98M1LUdebBJgZ6XTY9zUgyHzWmqyXg9jZRSpond5273TFThmTp+Tq
uWDjUl7SeOwwkr+WbGTqpWCo07iPEvWg8KYrs7PKL1gFcTG1gr7dwoTiFxHJ
3vGu9aMXt89GIyP7z7ToZ7W0a1xZiUcCi8w8soDynMcigEyuCS49ChxquMOW
vj1h0YkMQuIQYrRAqStA6sJiIpuYX1iaMcfuv/UbOr62ZfZzhfA0nD20bzki
Jhr1s+tnI3hNbbB77Kmi5kIe+SKJdUfxq1HLqH2n74jxqOJZdH6n9/aDPZmo
g1k/hS3Y+sOi0A8RpBaNUAK3uZoNb/xHQCdavNBl4Z1Z4q2eG2t9CyNaNOzj
4LgJCgpSRwIXsc3GHYUzbp3hlPHcvqOgvS/fyhhV98SQVi8l26AtNXnqCHYp
eLrBOWAQF9anehM2vUUNJT/0zQMn88NaObO4GoiZbAorkdgocxKhAXJWyUhu
ePyaOt9ZEBZwDMpzi/gypN46ypKrF81fMKskHMDTHVIQhDlF4IhgmjA27U8g
F0nQ9qEsv79kEgRWwDh7bUi3RQO3yEjq5O8rIPrcGNbdDl01jx7TJKx8qbe4
IvsHyQCqufwiOhHrlqDf8JEgNSWtPcAALGFfs5vYGxZRRnOZRIofqcxS4Zov
v9qIZLSsfI4gLpTMAKA+kcjMMA8KAl6tsVPosidK13vxxq/whGe3Ae74jXlv
YSAIQ1OlUHCK24Wh6DiwgQavZTiSqVRlQer0zaaXyMv6cd4P+IRsgD9u6+lx
YAV/wMu8kOh55CN2mev6XtWzxRLMqjlHDvEo+ISL91m2Z6GW0booKbmVrm2z
Yeb9G55h7Q5Aj9JS1Ed5k+azoA65VTykHA2n0BAHEHcfei2bILJaEnczDlxP
3sg5AnOcj4Ykbkh4lyG0vrNHEXN5gletibpb0771BZGARd1+hUwr6tCkSeS/
gc6pEhq3A2NeTc6dSUrXNnwB0AkYdqXOjFyN24cwdkpvv8j6XV4qSZszljRe
C+38JOgeJzhHC0x4NMPgbwBKtkX4KRGqeWBC565BlBY8FXG3nGpQIWAYOM0O
L0ETho6DLeNd/s6ZUXceHOnEOK9hl4jIDnfZJIMuM2OIbilv97sL9at4gEvx
IIp+8nsM7UAGe1XV5uEvQ36vHS90vAo2Nulk/ZCYRy1UJhXFET/Q7Bk6qaXO
T7L1fzfWevcw6KVbjkO1G1BMJ/ApYZRaEJ1h2s7ZVWsNWdvuZcOZ8Ax02GO1
9cfqMht1aoyMfLpFeBltCwE/9qpWgeihoZxy96XLlFxwfNCTwtDYUTSButhx
MjyZyYEISc4u/nMBWqALD9zJ30lGBO89oBZquU59SR7ZE6BgidTU2rj2QJVr
zsmcwr45WEv6S5gNpoWglBhXTSgpciZ16abrlcZBUwegcpFwBH/vR0bHSjuX
nUWcdDzgFqpyA/JBr1idSlNukhKmflsYlC+oB93frKtz7tiF+9MuceEAeC8j
C17qTYpmnzOm4z0EV+Gd2DnnJ7qfSh35jLFjtixUoinXDWblmRyyXjDCb4zd
TV4N2SMXPiS2TG6JVytwBNSomDlnYQFDeiWpweUe+hyhxspGZoQDo7dLcjy2
qbVtBgpR1UyXazJZkIlDxhlDIIvOfgGlqFPDCJfjE615MQiwlbWjLeiyz4aO
Uwxiq10c8cza+PClAkkiWAsAa/+MIryS4vXQWWAAzstyOUwHHZNsMf73rTWH
02vfRVZ2yW8YOwJXzmep0TJQNjWAGVjNsuiGCr39W9vv1njLEXNBmS1mmVnj
8FgaCmgiNJzLktrQkTPiEg4unqz+QU4Nc3z3pVoD6M+8PSXOTHlyntlw2Cv0
tts8Rjw6xXDIHHLR1tPJJW6q+edj7x+IQi/Vxgwp6zu4PHPFGG3MFukdkK8Z
9kp0Xxp+6mG92/bO94ermDSrbbXIo4Wn+5ziMwOesisNTpTOQz58ouuTDZaG
pcM0zj/dUu1qzE6NbOhVGG09b9wUDJhy6UmJwXrUhSPO/kBZP6qLNGesF6ke
Ls1kXroisljT5UnF1Ffkle0035ssAJUw4lLbJ2vDwDYY+/7dvffVsqJEpzk2
1XkhOYbyM0naMh4IQPjLtO+9fE3ZVnllU4//1cDAVXw0iyURE4/oDIT5BhXS
WjWNlAmIp4+77m+0BOs2K3azObbHSfxeQfsLlFI1na2geI4aABoRsQT5fqXi
43QkaFsNlGzUoWfU3ptzKTgzt7nRsebgvJKhQlZMUl52WqUpcRMWWCIgOLE6
a4BmDnRPWVbn+NLUfx7P5tn770lRYmvFGeUgIgk+EuaukdsKjRB3ZCZT/qMI
wR/QtW6LNbHDOet1Hpz6O9Np68GpM1IGFppSFH1iop5FRBkMTFxc5R1gnBGy
u0P9uTwHYR2O5d243GuRvlzmMtFrqMQOJsvVrM55t14yJtzDzPGrTXaI8a3f
n3hQMWhsccZsdIEpgSzBGmP1TEs7ZiCRozEYZyVhfQfQV1ztp4rDbQB4xwpe
I1bUERtbkGoSnSc7Vg0g6/nB2VRIx5nNxqYiBf7WFrD06DhHK0AJSSHwub9f
E+uax3UbPu6IBjh7La89gQDgRF08ixT3jvSgXdblditxpfSNyU1a03cxlJUx
H78QFhqqXo4XygSNTkKrh2H/GXzXj3S9s5LS7txkSlhBGwUWKt/ciQK7BDAL
uafNBAALU1zUc6QGBhr3XyX9RTnp/jCw9fbUO6P0gJVr3reB6QKLleKrAT6O
owui+Dou91QQI+ASGSvd5kHgWWdw6zXepNzHMitzIjjwjZkY78LKwvg40gje
VR/YiBq9sB0CPNOSwb2ZlCIbNtrHCOgNmXVa8udNUCjZuGwXU124REpIAOxE
WbNU0tSFteLS5mdQyI9EMPfgBQXqOlbV3qddyNRNkN60vS9x/92KBCC+laoK
re0UTSx9CDZucWqLYJ1/wE/RPC4zlDKzFJURERmghQTeH/yePzntQ8mLOYTo
9W+VNgcrRyhXk+a4IcccRn/rrGwEQ0hhG8tGNLyDXpZiLn+7Do9zASGVqQd1
PErNvhFurSRq4cXQsUqKTWsF9lRYy3L+5D+wsn8nKjIkh9fPuV5LKfcp9MfT
Dn2PRBPJsmvNGXuqeMEpAjGS2IfjbYfg4q4hd2IioWYtV0RN7QG4HEW1U+2K
bC1mzNe8+0LhPQNdD+oBcLH8pJkByEVAxXn2BkgALVwo0psummtWRz2wiLJi
gw2p/UDVo/T2glzcGAifGbAlkGLCPqjsZvD1UkqsPmLir0EY+WTilx8Teg8L
Zb7wFA6a8Rb9gQ9++f5/o+dehtBaWkdzhsE2tQK3oFYvikggH7XQNjQycoOn
dupqjRR7dFs2yqTuy1fsiDEMDvGWbJmRUNiOVuq9DO/OFZUdN1fKPryINSlW
WH47k77lZI7hEdMgEAStFReJJWFAiBnHX5FHHWQ/kP4/uSmI5jG/2G66JSLN
ZVhObGE1wvFJBvN3h91fxwuzskJ3cjZak8jvRxjp+ZlQ9Yl9zdSWUsfC733A
haCbGMbXYwgsTg4O75HrYrb452QC52zKdmN8Y4ChOFVuiSQ1YV8Shu4K+qtY
PBDdEDDf/MAmYtgK2Sqtc/CnMyjfFTp8ZhyaVAF+Wrh9Lxry3/F4uxc6P84H
C7yJVWYSFJWOaLzPT4MwOTDQK9pR8s2WRoxvSVrP7Unma4Kb547N+Utj8pKl
vg/g/jYC6/O3di61KH8wcOX++nuK6+GavfLSLc9xQV006tQthUR1idmLCvaY
zwzosiry0zeKybz96VwUuXA0Nkhz8kx6kW6Fc3YVxDzIUJp4rxjlt/R5KM46
+U0e8tNbUaMP6bJdn5ihLjksavdGWRx3SMOEsqS/wjkBT84bYS83GVDqAPBL
weosrITEhHug9T2L4aP4p9gqJHfINuFV0pkxBOPOTfItJuIg6YjnTqn36wGd
CNHDCuxN9wj1SMb8VA78vK13ocFrYOkYD9BMoCSF4SkQ7zfwhPclFLmv9zuI
unu046wNZru5q0wMFILPeUTo5W6LRvkKmiGNpeE66EYBn7m+ekc/MUxMg7ZI
8MQSb7PlYim42uOfhS3OfnWwCZ//G5F9cNwPWjKfLAhD0VfRpAIKBF7oU7sQ
jfae4dy/HixityLYTi+Fqy1p4tS/IFayYMWtsabnmXwcv01T5EBf0f2gP1fT
WPyTwoE9J1oHCU0lgDsyaQhQHBaaByTGUHdIb5X61aDQ47Jg9915xFCY/A4S
+VG+YaF3lxogqSPPMsvDfx1Of7VdtwiXIM7Im+mMK6x93E/eBv6bbZfRwuZ+
VpSZtfvrSnyLxj2ZVqUlsR2ZyYKzYAgIG7cbTmTMJhXMPQUUmxBGxV54ldZh
1E0QT5f6sH0ZIdERgtPR2h4taUj0hb2XjeHfOnt+S6XZpjQ9Dd7zrf78Ge9B
7IAODMDQemWXg9JurcE6C/rQ7M53X0WqO/Ds7KbgvsOd6UPLxnUmMrb/BBzx
sbY1MrpZRcvbY5g0Ua1OkR/d25Qh8iDuirjMjTIPlVkdy5W/Y4E0oeUD1ZtV
usmpGWNndEEnZWULeeCNGj2dxjSp5XXZVsfGJwY4eol6lZHs8BOJxlzgndgm
HCFx1Aj9XZqnT7jGLpx/FTnS61kNZnHWpoR5m8H6jqyOVW8hTb2lOc3ISu8R
cXk8WBQDwtxyhhlhDULhtaEBm+Uv4bF1TLTCGEFtZwLWUwW9PtR8vQmZAmSb
do+9kI5yMeqzq58tmOr516A7XfLnY1x5u3OYCmLxL4cirIBJ66gflo09j8YB
xFQllViSrgltKpHbOWpGSOigSjINmBa7mZddHGTeUucWp9ytZs8sR0V2a1eP
Gvz9zOR55VNvzZodRVAr4s+oLpxYFvvZG+nWkqIBJlwGR9PSRqRZvTH4c0/2
ruHPtpWtCGPJ81NFc/ejLGaQ4Dzn0CmDdYgo+aSDySuAJ6V1O3t5grY5l8P+
Vd7wxILDrOUBRmVyK7/ItxmMLWjedNfrGhKG74BLaywvEkIA0GXcquMApp3L
1RUVcpyUTL8mldLByusu66Q6JfrOfeeN/J3NrJUA1quPz8gywf38VuD9xFWA
xeo87UO+cG4S+ezCkcoPCUYPY5wZ9RONGoKtVqe1vlI4ZMZSmHWTxjIkHhZL
xHlrpQIn9YnrZxza9CZKdmet64UAiACPc0nR/jnw/n3OLrfOCURkhyky+Yc5
tAWc1eTDS1zrfpFUXTlZ4tnkZ2XW1bv3y5NlbexXoXfGWEAmSFPPuzvdHWYs
3GACdLJx+9/xFletqta5/SO2oOQ9h+86u4WToI3RhKEvoYTSRA9GogSGkJx6
dIgO81ZPZV0otPedLlpfAAg0i/4/gMtlyzQ2gLLbtTuqXsbolZDKwDVR/z24
1ZSZwOGhghtvdPvoov2gd0euTzjFTz9Hu29PV8rLNy4SARqPVODygcUH/yrA
kwK3U05n2WbzS6QOL9jgni+ChH1OnWZPjYeFnVm/xCcgbWGM31Vl4XXJ6zM7
Lg19nc5sPOc4eAmeYV0fcAagGUClKwryaj5x8WY6/TitRqE6p/QcyOwC13nq
62VutNMZ8OHCDE6ETN/fuw/bdhYfM6WT6N2f9R7jTsrnezqr2wIwgVBWs2st
wye6iCedGGdF0IJIe+SrVjlDDvNLoswYKeraXOyUyaxneNhQeP/a9uIKUbXX
wMQOlvRFns+3TkwAqbjJUFr4IkqDvkefY9GKQYxVwcObEyHnifwYTMPrd2ob
ywMICv8MXauFVwP9QRqUz7h6c8IQkII99U9ZD065zszGxV0fHR9Yx9yYboPw
sEJc7+LV0CDOgS2esKe9gK7b1kBF/kRq3CmcpR8vRvqbL0Vkm+FiZmlwdIDF
DYxsa8CpaSWE8c6USsVvSGRy8SKj77vxkVKcsAZSLSBW6AgGZiePVDGrYujL
/tRHOD2XbruikLKFwVh9J8hekz0mVbxOJF7ZjdoN1v49eLxp99yaB+M7nkY1
FdyrX6hNPd+oCMo+uWLbbgMyL2AGAN3e0WxFV+ZMrjeUMO8RLOxGo+tJ+agv
nKxudo3xm6/PuW1SJOgnuGPd51FjY7oQqAW47qCUcAftiQoNEYH5rY6BiePP
8qCej5iSD+DCud61PIZHd0Z7SSIOCZjdfRjj++dcwcm+AQwle/LMH8agQ9BD
tlWJ/v01uvZdRO1lEJxbRDPy9VPHn+gXCVFbtTnYkuKca2ZOPEjnf102O1Bk
NtFxqEXLPrKwuyQ6MHzkzJIjMb5rRZpdZ80DymmEUz65ZdHpLVLRl8hmmNy3
MnHHWx/IWjn52A83TbiDxlFPmOZLPJ8diP8JkU/7ehp1X9ufHjD5EXNlzsfI
+p59BmEgnQr7fNnPHvtCDOGJdqwRcBJzQa3Il4rO+FiDfYMIvZJdWsDt+czn
cn0b099wRubVIveDLzFjhQNR/fNL4NSlZB9cV0oPBvWu+11D4ep/xfIuXbXO
Wa1PYfUFdTFFeFJ2HtT8qKBywQAaekZUGATpB5poUBVKHnda62s2gI4i/u7W
6/dcVbENSHtxLAnP+R/sv0TUkhZ5O6kxtyCbbrtV+3+LGm+CT5fRW4PYMO6e
6k5atXB+hwYGvAvVQ66153QGgt0Cv1R4v1MyKNC54MthK+pSAjIByjY4C0C2
e3TRX+LlEvXpoRmeMgPXWPwYIOLcZ8WD601T7CkxxkyM8pnIQxhVN3a6JDjF
ercxDpi3wpN6TiD8VVMhvX85t4ZatLOMt7I9iKRownA0cCRrz470lkLlttMx
xTQavwpuW07P8b/SPrd0IMNciWCR+5uyCrwWARtayKmkNdSeRI+48jlRVdI9
OTL59SHgdXFzdiPuGgQ7mQn6Vq9EV6OokZ34JF4K9bshTTHV/Dh3FXbQ/c3I
ZzxbzHhOPHF6tMXPi+Yu5NTESiros7LfIs2zCJ/PaqW9zIshtpqoTip+otpJ
NpF3YbmB000Xt2JHiviRhW5JEVrjgEXYimnCCz11VHCotUqxgoZsDxqSmGan
yOKWNZFyvcQHMdx09Ucu1qG2QCWgQEsa5/FLtrG43oUej5I6ZexAQY5O8m3Q
Vr9+MWI8Q62E1ezqrjgSfxtNgcNGbkbDd+Th6owqyVYP5DXW70tMBhfLGDXZ
+au8L8POaqx+xFUe3MOX7gmHllsPRPEiyQq6skjXjABA15JQtdanz3kFIrbc
gZhbVqL8jU3HcYGBYtfmQc37en03F2CqJ7weEHiGfp3KbNZJdT3qKUHH0G2v
3ozZ/EHoSyMCdQv5LH5jg9nbOb8ATdsClsUmSAyxKmXX7lPegMSBKpD4+8uH
lpGZY7CtSoQZA/CnBxwiZho3toJBzpG/TNLTaAHP3ZqZKSdT2L+v/5107yh+
JGb6mm5yVkg4TEvdSSAJP6wyir0ZC7TtLWiEXKqhnlgkKmYKvaQXbzZ5EC8K
x1BEKmL9i2akmlP4zy/93kmZqsmgaQl+UzjUiWWPlx772t13U1K/ubJaMM7m
hKEHgY3xx7pgWwITDAj35jdXJlrKs1r+1hJ73YA30gS4ishP1ihyqOjuxWp+
HU8TIxDOOuBgkDuetKC6VsP93FK/OW000gAEO1N33hVE5eeF61GQOcWnFYI+
nsXfdPK5+nNxTmeUXr+NZzc+iXVCQ4biYMo1k/ijV+LRZXQgvnK68jwzPqqv
o7nC5AUq6YVABUwk9oZyDQrLk67DQqE5lsZ6osMmPnLdnjrd95t2oZqfY8gl
UYmH1HlzlZWGqKZRK6Wwu7XG+FoxS6+QLeGnXLSiDpKfmLCBuv3uKKgIMG91
o7Ny03akIZ9WTmCauvfj+BwkQHqClRUKr6c3d34FTvvJkuKsB48ZyFF795FO
NcXmgyfI10G1F/ZkFvb1o1W6ZDOgjs+RYCUubnIBGDeN1JJSiGaPLmwT7CV4
pSn4P0BCtClhWhLYRTU5Y1f+keyve1n/AhAXu7nZTeD9+RIiRGk6Ncdaymja
rYjcKSKZffBMnhYf4VX5xAWwc2zWNc/8brJgw5VzP2XbrVhCbVLa/nVpzMgm
dJgEKasKexGEeHZHSchp+n1urJ6TpcWkyqq6xCi3YeD/yVoq9OrqCTBTqpJx
bbA+qbmgCqmTHFZL3ggCnQlVd0yCVjfaHM8ThB8PPdsZoyuY/EvUH91U3V3L
0JKdQZp9GqVUOOBdMZiLceasfRSxRscrT4yLB6AXAPDnV6UaMA7Znpi7WQPU
5/rM7NN3+lzrcF5eOC3PVzAINWnaxnIcVFngZ7vtCaw0SiUkMXoQqUXC9eqt
rtjUjGU9yh2+qBawbfayTNzTPAB+ZxP6xW1QHd8617tgSVdQr373A+Wg5K4A
hRkzGOs6d4IuMKiSk+ue6ZONEIyNIxiQsGlBiCsjYS28BJqumcDStafCrd3i
XTkEYvl1vpjOP6aabfS219gZoxDTMBWQwV6vv4HdE9XCrni5qacj9jQF2MGZ
hpjAGeiES/nVLUEaR0jJclL9acIBGOetRTp4+K1vnnAWEHvyudRJ7l5Qi0x2
hW2FsudIsC75KiTqyBS7s13yLZvzQrR317pBNpYCXXE7MUhIB34GIjlXJHVw
VGWKvGQbXC3AQCvFGUIgWs+nveT/cL0Tq8E0AJ7GdF9TtEwPsdehqGr1hi92
zQnbbpVMaGpAPEd+yna3q+nFEyl9QZPlmpk4toXht/H8/5gZGf6AOLdCx6Am
RzWsyWmFfKqhF2JzzR5uKRa+pQnlAGqFmOWa5PJdsxUquJOdtobtRzxYXPpU
ewYrEYZ7gacSzIj928Nl6ysV/KqzzFEr9FTTF05es/rRmNZVJRwBwfdzehyK
Q9oPATnXqcxWGUwWwhmKLlbROrn6+3yaZVHxxAk4jxBrD2tKsIrBSqpVE4W8
KER4VsObpL/mBQk4Vp/3rea24Z1A6dVZWA8/naqWLveRb/Vw6RxGbB1TRHFk
KSO6mKxZWueaBGn3/5THVsxAnwq7dnZrJMEnRYy7bAiTtAkDjXEa1VLb8SCL
MB1wLJK96a73Hz4FC3U5k1fAf2kUdLRFwQ0KJZ19L6LsZOgEEu2Wxdzji82u
HIkUgr1C+YL4/1mUgmru4k2qXJlyUJIBFXDyCjj9rWc63vN4EDK29DccHMg+
qVxYBGsDlgKOW5ksWhqB7cD02jxVma+sai5f/U3Ja11erW3qaccJEpKQ4gaP
qYOTbFSlKA7A2fuIQvQ7ulmyLDGOIsom5xSFwfUroMIJWDdZw5en4OELjEKa
dAauqK2j2tRuU1bN4jOjy4DPpAcA+kZJ3+IuIjN8jm/YPNScpnS8Ho0+tc2q
uEU8m2TE9nfAgAJSAUqr9nNYUMiopOrUa8JBsum3EB/LBwZO8iXsXfkw/13a
fyF0Ed40H24P5/a8+J3QXB9Ktiu9D1UZWMAQViKQ1i8ZOnz6HMIEMU5InwiJ
5iXdxIKHIc3dg7TNiSm9rtO/i7lQlqvUEzBWjceOWJmEM05/n95rPKuNtwvR
k7mjBF0hETqC3GMxa6q5P1gTBO7a2HQTys4xcngua8V/ScKORpffvnC6W30y
GUoR5Lq2fEkJOArD+InCcC2ySzef62OSpYPWMJQu0yL3AwlPKs0ZSulm7rGX
tqX+x1iEgXGfTIprZoLAgon2rDsoNrjeUAAp+qYKaQuhIFuJVtb4VRYIoEMU
XIiCZuX6RTWLr7r/cQnT7Q9W4h2F6RFfz+YOScow5GHzLc5ltsTTuffN67wC
y/euunxXgTmoR+230yOCtq+PRLitvYXwifePC266VD8jNAOeL4N9nBBqiKRJ
+MlFg8+Hx9onDojQ7bQlmR308LcU2RGhIL8v8FlHsHyfIP7obWwvtchi+Iue
x0UBVZxaFw5IT0oxZ5e/DJZWzOMJfSMmnDNNNMB3gQ1EZB4u/ObdnRJji1xe
PfIxxsFV/DGPPnjVvmREThmDiupwCBR+ogPoiuic0DLJ0+GPjLoNyAQIo8CV
55Eh0I0c8etY61+uU8xSHmeklyaLGU2nXC0yF0x2591Bg3n7ODqBVWxf6KaI
Aavks0DK6vwN6ldjiYA1fUFULTY3cPSAk/LVMpJBQ9OZxFbtFqMND57OCxmI
MBZK4I4UvL28TqnMIjaKg6vU060bIgOTlllovMq+zZ7kbyuwnZCZl7YsA/wq
OWOIdinDaUhuiCv1vJG9xXqnVdG049vVr3OFdkmHYzgCXucV/S9L5bIOnKZY
Czu5s19wllo3o0ZYI5/SS0+EDrVbEFj8oIMuijHWzhTl4sJAJ92q+SorOFOr
j75mP/si6pY/uaEIy48XBNd/Z/Qu/YENOXWb1jcpbzaEBxaaF6g5BRjB9W2u
D1k1W6k5o9DLhVNSWpHZEhtsyGcPC9JLrY9q5xJJxLAxbUvLDxov0tX5+kdY
KkMMu468qiEHG6rgYf35gbnvtOB0C2Y1Bov/kD/lRl6DrxBUEDWOA1ymPjc5
oQ4AWR0sdDNH8SVbhcFpy6+bO4zmHc1TGTBY27XlLf0YcEoI2UOr909jPajm
xtSOGa/nmErgmdFB2Y65uDmib+x9rZmDMmBtBmjvP6G/KpJPEU05TLdQreYj
ITHvBxWA/lvzCc5pGCv8LOc+/J6QSdYJsbfNcOUP6g8g1mBlqdNt5qdSM7bs
O+Av1sAX2eXSkI6dIk7qInQX0VhYAgncgbWTQLRJoJDFPySvTgGCa5jUd6nv
kQcoi+FnTqgl+6jSj5MABRCHqqI0SgSIPfJLM7p2Tsp6RPRrep3ZpLOEtVNL
xrv2BrwsZVINWS84zNOatZ/tAymv1CKOXFJIvvSicz57d9ux+qyQs9P+JbPU
ty8BZUBDYguU3t3XzKh0imKEoJpEgO34Z5cczVZWW7UlxLHeX8kEyzipgMD3
pkVnbjtOBxC0Y8p3mNUj8+iX4vg1VXdS+dF9ULrGvCNpIigUQHg6KGaJo5lQ
yXqovliohOdExfeSvQxzegMPabgtm1RAce+Qs6th1c6dXedrGhZ8jlCmVH7F
XmjwTXMppD3yzuzhZ0eEpsvh40x9lK4g4kQYzH/yASPc2bQWLPgJ2/JWj4qA
1ru7pibVrJ2ahwylQMZyxVcCv1GE8z/u+EhAda5kcLzgW75MECoZ5f0hgw9F
b/aT+AVAxHJR0flla2U/GhCdwRdvolTBOwZA+oaNKL2GG9GCPZIq7qUAWlyr
x+tpVrC0hhf4yKq3D59RcUMgurVBfH8RQYwXKxRKeu+OTuLg9yKqJmPPqeuo
hi44EjYDyv7C+bU5H+5swah5m5D2eK86rVOX7P76OyaFwkLnPSjAHbGYgeMS
X7I3yqcjv5pSbf5raeMWKfUh2z9EYreyaJx/XdFwP1euFBC61zL5orAXqA3v
NJoq9A66RjrvHek977dugBSQvFiSGDtv13KAcn6AsJtP/e2j5A4PApRL3yVo
90D8FdB18rB0enPH1GqNhg+hSOa1tylm5c3ugWWQTemVmzdTQge0TGcf3ek1
79leUzOcmrQEJdT5jHNRbB+S4Pc0n0tAwuognC9Jzek5Qwuap6+sEMu1d/MH
PJyFt+XG4AWTVRG73Q0MQSm7R3i2DwJJjRSEQRBbPD2ZIPRR87Us3PTyZk3L
v8u0ScgAcHEpdcNidijdUDvQceGgD92jXySE/PNceQz3EcKECHfN6iPIBDsE
XIl74V5OV3J4lGJpzanFHMvtvM+yX+D+yPaRXYUR2eowhEDjv1aQNZgzWLNt
qBgsDMyg9MvQTWiaDOEcHQ1XkcmucCGpnIKkBwwGa/D60Yo6FoyXIlQLzMQc
3gj8KQn2+nSZd7xDoMRs5tjz1dgM+RrjP2Lad3X/SgLCSR80cAr7QY4Rxzww
KwIby0QEfq5CdN4knVkQ4VlRyKMwU5J+SnBYCiVCEENUu4sdLBxPdwDENeea
dxyEYw8DOTtxDcST5DciXXPlNFKX36pWPu5jGwnBYVo9s9qJRig5qh4rwPrG
KAEIOTTXMncYHApVb5FeOdHyILF8NZzocn20YVXSnfBwqIPGz33eGnaYcQuE
LZxEUrYYU30ekIfjRl2vtmMP1fQOFIW8j7V7Gmld5pfNPoN53MrkxclnS2US
ek+o0CA4KPPCv8ajhn5P0H4Q0Ygl3F6vtonqFPFqKqt2qozuqUWCFBK2a4wf
NT2+fBPzHA7KGUcyfNMSsdwGTGH764m0cUZE2wqsPWspkz4gYKOTeY2JRvvf
g5XYDNNDdjrM/jey3qy3UX55nFe9ldi1fDd/1Rz/nhOt2apkmmhFrHkuaW4H
PSmve7/OH1T4LrdKfbr9MaLu/YSCgn93ItWRQmwNtaHd5kRXS0MG/ss+y3wy
xEJXW2i3g8lM7uIjEyKOM7G8PpunxBXO6ThroxpL71MCSFVGrhf40qw7AxVe
nYbJetvJgdIVAitCITXRqb8pCft193l6TyT3NK46y82zwGFAJ0EZv+RFG4bd
WHtEAZNp/V2vSsQXL9S0pp3Sqs44GKnwmlRkr/1QeJi+cPHa3t5iWXSN0xhE
TtildGPJggWdBpUAtN0/g0OVpjm2avzjfi/Rz7Q6tJArKWGVI+v+ADCEpu/C
3kkHBryCwXXPRTHOCKLGnTVa6fxtdsfwRlReYL0G4Kek0/bVxFRnPIUJasSM
bkuIDe+x394kUtoGxOK7eNO13F1P3BmvNVbeCGiTwPi9eQcs3oN2nRsIOX8+
7l3ErF6tPMkTAozdb2EAsEkMZI7iIvCgHjwjD0TkOTYYla+30b3KYjVJoZQp
4vDhJ9t++1tplq5DBq6gnX5PM4PE1cLf5P35QWyRSGrzROAFqKZYJ8jkSPLY
HMkz/SHD9NBBzVJlTpRtsKgtNRViUtQN8cdQHapvGibvJ7hIWOyvxzL1Vk9o
vao5MiX7is8SBhzDYu1SY92/Yv2ZrW5NoJLkKPJvoN0Jm8gtQtcBbadUP+e0
XFKGyvsYptI66FMuCww5Nedvi4ZVhqbeOHFxyd156yRPxuuOaOyA1xZLjTeJ
fcPQ8BvORWOheeb8L4fgxWvTdQ7hzocx2tKE7dc4AgDgFyJmLDcexq2U5Ogi
Omx8Zhh36B00upQeAarTaKN4SteKAdQWaFSQ+9mFkgZ6fQldppcmv7tS1bvS
teoDnx+8TgPeLTKW8qW/1NdXYeaP3LkXt7dt9uMjS36OVZm+hgscViqy/m8V
JlETT0lTWQZ+Wc/r/hm/TWTiO2CerLg1bforUBazkNvlEhMiYwM6cgM2F0E3
RzTt9EirUPCgZ6zdmyq0kBCKq7wFZNIavlJtsjpMxXcsLHXnst+yBlbBWcH1
IbM/oZA3OCYgNVlVdG1F5IyLTR2aCyjyR/Q+Mftj8nt6wc5+o0riOjuYQWIe
mHERbyu+GAqoh+P3D+oyybZgA8Le7Q8vS7THP/CznWkVLR37Ewm4vNN9t1tV
TCYZPoKDdFEEIH/uKTIHOwAuvVFbVPdDBUxN7NU9euKx4/snwJduwZ1sK+aN
sdQd6IS9CZgq3RTc2pRkpsvIE+dxMTfnQMgZuUAHQGZwN1CQeNSpjplZblEN
vbcN1Sb3S8vfMEV5/NZRMBeO2L9yFXyNjhMCGT6Ww/zeehYOvQA84m8wtyDX
SBH+CSUXBcKYu/9PxoZstXz11VAFnsVZYb0OSSW7BuRIUBtmYZF5fMY7mZ0V
p9jQ3Cl+9R9Z7oQ6IgvAeSxZtsJ/cEfS54OCwmL9BHe9S+ayb9N8BM+Uyw6Z
pHl4XOP96rHS74O6HsRoFMhWMrzhKbsTN18XoDHpYISra9OcDHeD1rZ2ke5x
PYre8Qr8hRiIBKIGl/x/5uiWIdHlas+1vJ3K9o3kdTaZeV4KqPXq2OQwSV7a
uyzuyFueJhUquGCYY9hTseZXF222HfVwIigVpsA/bhEI3wZauw+DQZd+VW6O
RES9xeKpzwGokbMsPaLKMwqfdq4M+eyYxTUOZU/sgR9YlLh18m7UGnQvahgx
3R7DJKO+wpLg9KloB9SG2jrmX3KG94T7vpY9HGavuaYOW6txjqWsfpYFjQnL
IZT7P+fc9ztgDSbVm48e0sF/SeB1Gyg4ZiTXLGWYcrE1cr27OVcBlDGGh466
y+9dgHm/4Q1KTG2yE4IPsur7iKL72METjxtI3khXHTNVVjrNMyWEzQqQB7Yt
FiDkYuPz/uQsQdSEyF14Hin2wyOWZtqKDJkq/9wWX1krlevp/PLNUGaNB9ac
2ivEYTk7jh4qVBzPyifMrI7MwM82v6zLPXaRl+AvWIDj/fLmx7XuFmsyqRl8
BkG7nszS1STQ0iqpU2Me+5TR3BuiB2F8nABXBB6FtWN7ilAhVLnYuI5Qnh/4
B29g95Y+AZ76WNTq+MrpZtWdjqNk1iKmQPYX6kVjgQl4Su/QqyMJ03UX3omu
BSQyswbuIWmvZ24wo672HZ9VtnOdQRX0iwN0rII5TImWeDXt9BlT0awo23cW
S3ZlAz1+OcGN3YSJ6ynbcyQI/AbzYAtn/MZ1NEleMUw7FJUOypaDwJ1kXWOU
E2p5MFExCK5LLNdSZGk8I0S6HVdXakLFnqpDbT2eoswGtsaXz36THOcBTSIl
QKLAcRcHXD6zNNxTDJ5/QuAYci6J2nKPVy52tgUT/+PH7T2Qu5z5WzXQP51V
ihE6SchE7J0ytIGCxWfw3aHYVy8bwoFS9mA3tQpno23tLJQ1vFtRJOUnVY5N
2Rz3A7q/gJMp39nqRnJWK0sxC0UxkHHcmIViM6FYddG3N/mfe+MWArHpNvLN
JxsDmJ5ATN9g/aFFbYiA1NbE3Bi0fPLDLfoCDsvaSREOB68npDLMml4Vap5O
AKXeT3aqbkRxvgjKoyg6zIpURVl8E2yVJjFojGgbVytyEycoDZy9ET+OcdD6
wuSfLa5s6xOdBNKCgN/dz9Us/oHgjfgKBrDZJ4WXn2ypO7ye1Hy13Na0CgkY
aPGBnJWorNg/6m7EFpJRYNjHzjxB0fjhG8W6LRa02tNgss1QlMGH9GlxwGMM
XMDsiRsCsBvuBuxmbKen1KrUYOydUV6TFRJpFhJBZhkqT27pQ02y31VVYTt4
ih6/2U/7YlrY0Z964RrNFtRC3H9BbHzMG/482sIviZTMjTNjv057wAdw1ar8
8WWegvy/ZwGeAWDpybMqIUDpRoNB1sZgaM4EUb86FjVH48kGw0K5qO2GTjuE
FmQSDMXPnqTqEU195cYxrww7dzzu0rQSXVjT50FHGV4tBTyk/UYi+X1Bcjud
vWj1F9Hiq89PerKn6MXA4jmLjF7wTw+ycjKSfb+mCJJTfAj6iFZJxovANKni
u5FuKQw2X/lzd5cbKcUAQMmSWmmVqhD7vO0ovS087/9UBGoZwyGRQ5T3Uxyv
EHdzcLh7eX9gizO5EPdX4MV2gZfhf+CoVAr91UwPt7mvY9GwwdAyzBa2iLhR
NqQH+9oDpmcFBGmrx8IoiTKfK9EOTltVAuN1M0XCNPEdQ6PzraB7tqEU0DkS
Q0nvWoAMTQOUVdKTdPSEQdMZQ1eA+dXe2VdGP00nZDCYl9DTWeflTSpM3U1q
54gipkzKUf6+ZTKBFOfVSgPpocCw1LwsfPBWfaKDcnBaNzvxDqc8Ghk57nKT
lOglqzk1hfP+7lJWfEd5ndhYjE9Jh4HlWcqhD6qYn3ZWLxW+gpHxqaFES+0Q
DGy2G0cxhc4uwe0z4E3sPqebTqvf7c24Wrf2ilVvWaSemyCR/VIPFBH2Ygkw
EpdORjczn0A2KjT+fOwC+DAUyBn4xxEQuZr7tD6CQLz5xGb/v9zrKIpbBUrg
zsQQAMiQCcy5v3RO+S1RVp0qUYLR7IHaVG74KBZnpKkCj463tJT8UoZA8FRe
2u8b23AxyGiBVwfJ9wmKY8HFOJB4gH4v46tv+d7/UBY+kVgd/tkySigYx9Ep
jK0woEPB2t1SQKlRPIhQgvaUlrYvTMr0zpHU3K86isx43pW0g4dD/S75f5LE
BX6SykleIhtNNzzqPYiLPtAYq12VCA50C9+7hCcDBBwbq8XODhRjcYy26NoY
ICJ43S7At/DoToqL58VbG92uGDnyF9Ib1gD6+afOsDPLzLVSZZnYerdtCHSh
DbPcyqaZFsP8j97ryTBQvQ3h1SDu2hrLBI9XvCJ8memXIO6VqgLXTB8XFeN9
qfpVllwndhpL2Ll+WG/ussHPfux68EdJEDcGIPXVF8dQV1pU59IkikS/DjXm
lBJQl172qxxG+BbYuWw/caFvZycCJYnH8DqFebkdjMDc0VVQ/Z/gPAOcVlUJ
g6Vvv3Sb0o/7JdIQMsEGc7Mt5IXf143LwzuQlpmM2x8w7/iNGIbeO/zfhonA
HLZgg5m5qG36MqU54ZoyXw1jhmNy0PkFPpvAiZqNcEejPzu1dIhc9S0eIh8u
Ide+ka/B9LpBtILAq4MJhSdOTdbVVr8ntKRE5iaZSjXAGmd8DxFqqOYr9Sss
HqdAibb+MGSFSIc3Z2hcIwAWVCLi+KBZDt6Oas6Q6kgI3cGQeoqNo6a9EGW+
JwanKIEWNjCccy88hu6ijAS35oRreZ/zv7RN2wo/CioiNBSRhjqIohSojnL/
GgA+gLdlQsj2zFHtPMpZwL+w2KnhY9eoEp97Au0K33wtekK4YfYXem/K2tBx
7MD6tz7EVI0NO/OIIY6WXsm1j/+pcE+b1PHO/EDshC+e2nRHiCQ23zyS1n0a
iRYAUo6b3GKgAduv89YgbptQvTp3P3JwDxsVYTN3eIlk99rWdfTUgzQtdQ1M
rq+wPw1fHQuIjmuT2ZlvgIHIYwL+v8tjRqopNPt+l5o9dmDqmhgmk4+nNS23
AhHTQucGq811VuSrCQxKG+VJTm61jvRlH7O680l8D//I0EyooIjUrgW5tUTg
6K2jzq36bvCy67g1EFkDjR7tc+d/tzOVFcj8INq28QHQA2qdBlkR6JMKKw+g
uDDALD8uwrQavtbOjSsrH50gaUcyu5VB0YdeqUM+DNAz4Z3+EZsGQDNmcmrf
jIrGQU9T2r1lD4mY6th0vYnCIUWfu2s5CH+6w6rS3Kol2wGSO/X5epMCTEFQ
HMsl0+4c+AYXmdmvQWwuvUtpCiv7OwiUhAMMIUAUWZ8tQYMUZhJYQ3AATCxv
cSChznQQ+Kk9OAYiRSEcNC23U5AVDncQJUWKKupEKEb7fLfL+vPqrdXtggal
WaeZ/wWOpVsZ0d0E9B5Ev/+8pbAxJ8AulF9pux0pLmvVrVx9X19YCIPZMCDQ
jKSY9Lr9rsX6LMpzt/IYhSGATJtWnYgn/gdAMAujp+h+1HmgPhPeiJCcQDHu
9I+QNzTTEPY8hXG2CEjhAc/jL3MNfpWXPPA5C1gfCNZuMHt9PPdJydFcK0Wj
1USxYU28lG+65PXodopft2XaBEu600ujFGLAgqPftxArvroGD6YZAIhBSWuJ
LzbwYIyM2LttXiV4hD/I6ye7KQ9VIYzGNggdIvlSLB5wpBjLC0IIBSoe68wK
bSYX3FzDBnXGDp7QMlxiQ+nL+NHvHbY3bt6FKiTtbJ4XPxER+blKVaEXJaQ7
V0NWtUq5soAsQ2Cwkvs8iOrMAdziUW3pke2UNLsPT79lc6GiFGHz78YvRcm7
q2iRwajc0AwXDwR4aneqLmPMPLSXeJRx4afaa9XhM3Ms0Q7R8m4cDlfTo76V
/y3O0jjt1hg/qf8vMPIwXJkkDNCfcQVOZDo14IS2it2vHrrpW2Vi4pGV9Ik8
HNavdF+I+MhqBU5VZAm4JrzMBEK4f0LKvt/33Oko4MUmSTCKnFIpuAye40Rt
+U2xjt0cHRORnnuRhuZEoGsNHy73DM8OWbgRZxn6hSFI+glUvxg/ROs5Ilyp
PkmpvHVT+ADeLtF15mrolRpo4NTQsTdy7Z6gHNFbcv+Ams1JGHaDso6HIEhR
Luy0unJt0CvhXMs4v43RZwnO22XZp2qs1TlkZaKXWE1Oy/DbeX43TiWtqIwH
c1TNJcwrnZDm3yq82zUNu8d86BUxz8alXLZVsQ1+5gkyvfiyWjqlAwOJ11d8
XRShdSupkAWVZ06H5H7yHtmNqUAvkU11gRX1CyAnG1Gce9fGAmUenhkWBrP2
JGrh4O5YwjqQ3RI7Sp/lctclFGx1vo11eatP5CPRmnxEn97VxxcN/Fx4/hHp
eyKQ79XTvrP8n0/SJqOTOGYha+GGbALyk+36MuhIpDm9jNVLhjftBY+t8cFI
A8ARdkdNcQ9lg/B3or6ZIjRMtULqMPpO8haQPag+MbhFJICdOxQQa6yeL20C
odZV29oJNxTOM6GOxTWgQhatYKAvg8blF/gfWNOYKTKcfgw4vOVdz23sDBFp
Tzpx7nGlCnprSseoKhuZIVe9H+z+sDsA5vrQfp/XLptSmDx5o+r2vcOPNgS1
w2VVRNtfMVNWkzsudXVtXuYWY0uIkKtO7ZgOwGKvl/5L/Lr3QQSz+emqIVnY
zfDjNBoCtyTvj0LEhx3tVH7VuVuWogxkoBDed1T5bQfFzapCng9mvJlX+Xh1
1V+tafLeZyoVVtXIaTwoaIhLARhIk5eh9q/oVuaux/vz1WozGDfHwVa4T1en
BCYyEACLL+rzTlWkGg0PDgXWq/Uu0BgDjJn29/IK/zLM9E0j7sSxcjpNbER/
aQ0xiMG5grrkdqcXSbd9z/nt+M4J25nb/k06FHfmmznPeKS+bQidzA+yQ+xh
Gvfpr9IKawXIDj+Xhc6JQhgTSV9Sl2PdYDcnpHLLEVhVDkFe3c0XfBOUstsh
eRx/3y8zewIcixKfjX+YgeTDoaoyCSThODZFGYtX/wENUxkHOoYla1Y0p+5Z
R59Z+Sj7r5gjv86QM1jdjJZzJxI8CLR2abo5b2jYnJbR9hqlx9iSWjvP+e+/
ul3ht/I6M8djyjClo0gdtlTpla1Ca0l10/FcXIOFN7hElPmqA6EXG8OtTxoD
vcNgdjd35eI1E79Ht4Y9e/jBACSlY7gIkghDZH77DD+ImkdKSB5F7hBx8kJ/
gRKljbmHiIQX8NcDJ4nAy0RGR82tzof44T3u4D0+PvaRhbz+kpMPm6fVWn2/
WRVeMUrSbMAxAv/jB8y9Fu7vhvV9lDAq9nyBC/WzzNoobRgdq0cyJLaBmhaj
udL4qMxwDAFEiLjQjY4tm5AUEdDnmPrKyf3/CuOqG5saHkEhUoYzn/8X6n2h
DfqkWUM1oyUvUclYdoGqoFRuXPJ8Bj4iz5xnMyWtAGfggKHWq4O/tu5Agkeo
GU7vVs6jgANzIgNYsmCKQO/zeMPBgU7ltkV7vRCiPDunS6jHK4YLa2hU/t7Y
bKmbe4P20cBR3OWUNIAOpQfrIAUEi26olrxplnDKH3FqMB3GU9j+fhEdRi0S
HQPXR9lod/Sjj2EMF/bKYtQvbtSR8WW5H+H7Ujh6+v/KaZFSEqrdQx/CyfN+
7lANdwmmuENc01G0eFkk5HC1kwPjUpnO/UoVVGmj0ZrrmUM9SmViscnR03W9
sbzyHcwUoAGD0eLNz1FqZXdOvtcn7dAv3ySKtpZZPf4oeC5Rjmzh8WkjIhE1
XmxSqT7lCatGbZSEljqB1WF9AmCrA3TPX/LwX2Wki7SF3EGmj4E9JKgm1AWa
8RFiiAksVbV5AhjgthPpNdIn+cEjlBXEWEYMHMIicXxfakEdWyVkM+bVlvZm
gxxXBFT00fugw1cHfgmxkLk0Z4mbA9+I9WBzMvb63DKGyXyLu8/M2k5Sn/7+
4Nej38CT2TYwv7mg7PFE7f/uOvMUkxLadHlfgaHB9FmAxD+KWRwyPQp1Mcjz
/wms81n57oawMVlgTZSnWjS195W0E/K5rfEYe8fTgxYVFmFmZ6qGYvUObqHn
5qpeOv9ocSMA0y5dlv7HsaUHS7VrZdDfYp0fiVIHwtkmIIg/1x8htz549Gli
u8qo46VGJmlxQDyktcCXZs5WyVbQTyOon1VVYRJ1ZPdLe3efZPnLhNydJbb5
tSl53XuKihOlPeoBLpg3wrl+lbVbANKHU9q8m1JRt/xXYPR+6kb46+QjlFBL
W/DQrLgZ4cin4mo4Xp2spowEByhNocToP+v/05It+tFP/gP1mi83LoADCyMp
bPJzd2QrxRaJB4NFPGqjdKMD5bpPqbR2FTJ/BGhfh7LoSR76hDPDqh3gwf8h
8+vavIXSOA3b4gmeJET9PWO2EJkQ9tVb+4L4OfnJz9GXgzmhaJFdhOrgOcrj
FeCz7oRQOp6XsPxSPsU6lgDF5P8y9hIZaxxwe17c7TUlQY9pc2jNjsk3L7vv
hvbCrKkiQ2j8Ba2EouWKI3+D4Rm5FXwOH4E33RQPdKA5o16BD1jE3CBAt719
fWXKFlhvOZgPuOAGJArImh1rhvsYvCgyUwO2Ti0xnHHVCegRIJhqwSAanxwP
b1nYvrhodzs+1rrnapKY8qGgsyO6AggwTPC1qwKZd7B2rfNr9MyIFWjD+GQr
Mf0TNAqW5ndNBR3DOl8U+rgaaaYCkQ1SM1/wttfkA7b/S/ngzWeovhxxnZnu
fjE90NuOLannrGs8CsSm9VQOYVtELt71brJoNqH4l2B8otOuMfT2N5NDGk+B
CCjuuToXVDW5d3Ht1qsPIdjdwRWqmPaccsJMX5zbMIgpfiijz2gR5QBRlDLV
vWPz2I79Ts4y/Zxqo58Hkb2w7nyUQn7znYsGNcydhkHSh3ib8CnoupHxF1Vu
dDHYFU32nE/mN33/uI77NZO8PPgr/NmBvBtnn+JIozrFsT88/kh6dM+EyCUB
R2K82nFahCD7I2h1MLv7p8YMeMzGUhqPEizwL7eAtM1nLrjExZZKrMtiN2r5
Z9kv/kfe01UL5OyOx01XwXFhFhyvGRIq3RaJb6iqFtOhipTEUQRSgYR2Qciu
PsS/T+11fQg0K2IhrBl3suv9/MJkFMFpA9iMsKLX7Ss/3O2ey3r4WwPdeNX4
cay/EK1PFqEUk9oGhBNmqLPwjCQ2Kg0AiqDVZkIsPbxCY5v6aZHlFfdPibVV
i/rwK9pNpbuDSJrQcitJk+CW9zke07NbjAhlg9MVisCQpeCc5y2Kntkum9HH
5vD+a7s7bSLYGzaKvwLkH6h3N4Tdn+1m4sLJOOt0CaU5AQNGaOBGM0of7DtN
sc2nFYjlbLc9BT+wPvUyRdUDAaq98JWKjES4+fJmQwq82lCRUq5OUS3uAb1B
JWoQlFI55as9mmTo2D0+o+meANcgyDvfB6XYz7Anr+BQ9TB5exwaRS3mC1uq
PmcVivzh0OU+9W0xXwuCJdbAMBd6VoZaqMr8m7P/t0428zl+Y5+PhhT3rWzW
+0jVSpQvK+bN9Ev2cjTTFb5D9Un3MAqNo2OACLkMIuiDA9+BLXCgfEU5c56j
zubIJ6fc69zzxoMHjviPdey2sevchbSNzGcHTnF/3U+DYEuSGCO5o24zmHpD
7EXzPzECrkYvYd9djEcZH4zO6smhQoe9ZI3Ap6rUSzYEXM6E4L4xagQWzTUi
6j4r0Z6oxQCbD5zPaF6DjwuOlVlCL1EE2h6qvZxYBtffAaooh4TX6Xv7vE6C
z76DIufLobbgh1poXPTCg+RuiW2TftqXgQUHfFDGkv0IpJsT4ebERWjH84jl
oil5rLbfvgXR64THEDAZ6Ya2xeA3yIRNFuZyib1PIPogy9vfcFR6I3wOxQo3
va/N+tDEeGopJKpTP7wbG7EErTXgIXIb1r7TrL8UqWkwYNq5xNbwbY1ZPvqh
6l5BVMmMzGOOQRSu7092ggaIrXKS7slIsZJCfyHvKVAGNMlcMyNUoeh56srk
rEZM0qW/u3R/9DVIAm3QOjmTqQ6k22yKXI6t4N8E3hW6KQwGpyfXsMN/99P+
zOEkOHSMInCVyewgXL9T3D23Hhoy4+KzGS5yF3LpEiJ602a13sFvnx6bGY2x
1fvMEBLtM6x4KzmlYoCmZtT+eEr3Q+hof6YqiNIhHUNC/ICiE8jxXUr/nwDZ
GKe2yKbE5YMboQg9Kat6OVuG+kZCpOcjSTr7gHs34VyAwrlaxcDLnWqbYgmg
bnt7vfug4sGFYnEQUIQUzWQkV8HfrP/v8ZdYXrcKRBv0+c+bWZeoMW+ahh39
d1hJ5CVNPytq7XNbDxL3ta3Et9s7F5cVPdDjqG4eGsRJOGikH2EIhR7S16pL
BwNXEV074iE3bhQSm4k6q1rGpOhIrMk5KFToKHA0we3hSBwu2IxwPJg4QjUE
D+D+Pxrk6uroFhTH4gM6ebpVrKNE6IC37+1TrQh4VoZrsMa/cLkkqn9Nm0aq
MR+NObFCZpj+0VcnUUv2cGORcl6GlWWkGIo8DWywSH60Q23Hcrd6KPN88pUn
56JUylVLl0sBGX5TXIx796RsCQIjmI/nq/mDcYg9HRCQLcFqW1y8GpRx3sKp
VW0+bQB3bfHfSbt99y27xucIwU8z2LdQH+kvrlmnvuWj/YOEWDPztBsfX9Jr
Nq7iLGB8g3p7ompiF85Qs4QWeEoszu2HZyePIuV9RT4vfwHFf/AkTIZwbQ7e
I3iOSXtRSXTCaTfEtLVGdFkXt4kEPn9OloB6MOZOnAjjqwVZeB1Ll2X1hwiy
e0PXQx9coP3E8usWWVSOuzJNvYN47UIA1svQw7LkAJFd1Bd/rODjImjkoeoO
ftiNlza2UUwylHP3FInovY0HZ6CrYW7+grJvuFi7qEvTgOq8CCtKTVKUFZDs
6adnbv3sD0EPHkHnHv96nFuZ0+vPCDTscgAQ+sttAPzNwb1IMRgzkXBhRacC
/Wxrfx/7iUbJHKLpv7W7NYsoZDIQKz/6Yf/UGN94KT/P5r2glTiP0xD/BsCT
/e7RyEHUcA4gA+3ERJl3ZEjSUkEjP165UKZvkLjBvZmKrzy9stwU3yKzTCZj
YC+BqOpo/jA1PqF+K7fNKAY0qcn3+tshLJW9LhbV3MMKl1sRoXg2tlJ0IHgx
YfUpvQzEgd4p3hkkYg8kTiuDgcHU+n7nBk2gwCKawZjlDpb74U+v6eB7+L95
ufEM24vZ39Ety3AG8w0/zhSDlt2OljPmlsGtns8c4zmiZPz3b/PaSMaWRe3u
l0iZ2LfMMfvWknGWByqbbw7Iz+sinOXYisS+aRo3iX3uck6WPQsQ692YNt5K
58aQ2yjd7gM/4WTjRMQ4b7LiN6IC6XP0C0FKkz0zi4TVMDO824nn62pb2Upx
FdLQkJPRjN7cipoCF8iiVulRNjHg7XZNnm4xVEAQCMqWKe5IejyBrijZh06f
51290d5ZIr5IGkGEYyaUEMVc0kgL44sxANPmn+JWwLYJLAIud3K16Ng77rRq
2dFoC6M69gkezhwzm+FAHquE8mplbpWPo31/jsVt+/9PBDDGrY3u0yAjDvjk
WbKIgsgExTdLc9cZhX5XneepPTZCmk4M0565aCRR6yChLgUo/AMP6sEDRqbP
Q/TG44frA5vbhGN7tNUIKhz51GPZNe7+GIaggHogWMqCSULlKXeNcbI9Dbb9
cyDO8rfJBA/BVEbyM/1AUQqH379UgadU7EsnpNKo09HsbxIw+G8HRdosBgmx
wHNsMjidUHJe7Yt+VdlRsCQWiOQmOIx+epv0z+DPZnxOd4t6LES4lqcwj20A
7Vu8RilPOR240sMCc+54HyaII/p+jLSQRb0eEj5Aa/PEn8QPVEKU4gosWE0U
MQSleVd8GyA9FNoG08eeQC8HMorDnsEqkdqdzP6Af3ea8nOHpS+5bHjdx720
zE73DoqDYOuzA98yOhZEJWxwCpWD5u5QEux8Fw7CIN/J8Tr9/RelglOmnpxD
5fsTjDsWFkyd2/AUZI4CF9ukCQJxkLfcOYfu+TqU2U9kyVyrK4sfBY0gNfh/
BQmgciGtkR+qcLzm84xj3yVS40aLG5loscIYFVOLaLs4e7HSXgiJCUBVOOhb
4R4Zba3mHYnE8B0xcnqpyenzCLPAgP5qBefLx1SHDN0FkVTl9f58GAj2soWb
I5qUDQXHTiuS2vj0/UzDPY3NGE7Qjj4vCYgi8IP+9XUnki88VSqG8bce9hJo
4+ltibIq+jAXCv2Rldcvzcqtbt3FoQmcKoxKuXKEndWI1rm6EPjRnxN9V4qD
AKHoxdEcA4OWnmGVdAgt/D9Q749QJemNyXMye78+UOtiiMR2bUIjbfwdB9XY
v4p4trU3eTizOCz8G7S1kouSJVMhWdOt/JA+UBhM8sAPUVyYdd0T/QX+VX8X
zLzIRdV294lhOlh9JC3jbgsEED9O7cdxrjASRmV5fL0dtz5lzKGnKXPvM9cc
vddBDdZC0lcJG8sT0z2zbD6EsT7Le+oXuOgn77gNA6gXlbvRicCzsTlOc6EJ
I7n60NmDBbxmigbRy60PwIKosm9zb8ux+oM7ubQfXqs4/uej8pwXJQcB9Tvv
Hpe03Cajd5UKac0vemKfe5kCqD8yBXPcYnQcogCxqIp6RqXoFkvbToA9A7aH
s8kiN1HaIghJ1T+GjamdWZ93qjC7l3T+CMNij8cBsjTzRPnkdEpTsL/iao1x
ozHlj4QJQAHjyK/m5VUPQ7qF2JpuLFSYmH5a6xFZOLJl4kdHATFd9ewkljXo
JO/Fba0xFvkASv469QuLnXGoTY6KWEuJV9MnojF6V6dZVYK2fPGIxF6Ss0OG
KRFrTpBFAFeahqE40+MXPu1kcffgOTFDV3jjV4x91r3Wngwq6Plh+fHPmXQH
HEDzzX5/4y7bFLZxLwiwOVeGe/2XgbCnZUyKY0R9udAoxutfJv1U/imx2/Ew
o27/x8XBpXA0cUxuIDqnYBbeUZis1i7YEiFZhDxCeczvHpIfPNyIK6zwXKlF
8kstt7qX8SgSnjaWmeO+fQl4+6PNIf4ow6nO/a4E+2PLpJ4gm0XVn4FFlz6P
7nNW4fbcBuioFOT+oV/XyTSPmZYY7B+VQC3yayg3Y86iW8m4tkXzlA4kGfRe
FFd8Q8wXKpCgyj8E7cMEB/gvAqWADwlEMMe935NtjUSvvxRm9SliaJRLojq5
hZ/aZHQX6T60s24hXYGHhMdHn4cenVb7VQaF0/VfHqb/nvNymCSmRm8oyVvX
3nsasmVeMSjn8yJNvONphsayccXWm6wc6VMf1PraKvnTPXotZqPsArqP1rVu
kqDMFFxu7JJHOJ8IztuyKEHZSEigvQZjFqwa19dYjMn+C3Nan4YjOs6O5Mbq
xVkyloAG14sUs6saTvpCVwpTSk5Hp93zHgC5KDE4hdkoS6uVdfLxY+bEJDb9
ErQAtQlictIJ1Tgf+5dFTXmJkrCAyC4vhuwEnoDZuPQKlAu94dKOLPjvyxE1
tQNmhDCBYpLhSKaFRAyQqj/Jk2BR9AU6PPPERJ8qb6oHgXWWVkcezekVVG8e
KKVaIp1GszgvLDioh5xOzaBm1TEjsTG1HNipIe2y3sxnO0ydinslwqlsU/R3
6nYIHAXrdKu4jkJLlGL/8isA0XfVEZGHcGHfzq/ZB8b6lyJk5Hu1Bz4cqUNE
ddHwbkfI9T+Bv4vliRmCWrK/D1rNiM/fKDjO3L6oEx/tjAjstf2yrMZfKQj9
yKxKFYt2NfO5iBFOUVA7ekE+KXHb6e/4B+wkR6YmN4e9slyCANN8uTSc/p3a
58Rt5vzAyP9Zv7oF8C9XgyXUVlYmPYGiAfTLGLFIzHm3uLfiHP7J/+TEx6HU
LM8G4U8DxzR1S94zxvWPu3GdkvS8uWAXmIrUwDuUHODdhIMi1PNx2a5neUlK
Nkr5osN/yVQbGc80Ind7uK5ajXb1JVqMzpwpDXTAs6PCQZsbzuZOnOl4kH+E
r4aS1mQEhY9wqxaxxTU9ozGB+wifoL9Xc0MLRtEnrQMu7ZsOPADrVjAWotzU
gC5Hba4n83Ogs2SYhfA6iTsLt+AeyniJqZO1I/tWLNHk8PYSHC3aVrwfd9oz
57sJVIBm+f3+xIAuhQfg3EhF/O2lvwB8Ad73J8Rkvo0Bai81wBTmTE1QXBH8
4PJTeJVUjE314H/LY+XLuXj+p0eysYwyN+r1wakQwvQvVcVzibGtNH1pWnW6
+ERF29xSdmw6g+QQQBOGhIMWvD04byDx2TRwrGR6/TJTRRpXh0nDcH7NYt39
Lb3jkV3qABRDw/lq/Of+PcOnQWYc/t7IPNoGuvEsOPCMt3R8Sl8EIKl9fxJe
Kdm6atJg4x+iabSj53Py5O3q7b5JshC32HizBYHYgmvVggDCm47NXQkehqbM
MJ/Hbgcdx1ZOuYpw4Iz1usi3kzInvs01g1NTa2H0nIVtbyha6Gc2l2hZzUY/
RdJC00hxHqDBsPzR2vbGyUm0/EOpAq0GryBsLfFMDXIxlN2UDXl4N/5DeN4E
+HLzJLTnspUkK8M3LthI6qWzRL+vzbI8gHZmLx6RdoHOVmMss2aB3n1if205
H0vpbqgVcrNKgeWV9HBnPpLYVpu7vBgzAyXqf0caqaFsMdmGdCEis5hcrZkz
s/l3AgiytTQBEh5lUEDMfx4tLRt27wRKaR/wbAABNeG13BRhNipf0Fw1kJuQ
VHfqNYVzthGRYRQ+3yQ+uNWvxVdLGh0dVaSMaGSboDGU6hP/l8CM/dZU3SGx
8DCM8P+/hwlf974QxgEayr55c+89+6aXg551pWqAde6SuvqkgH+BoMhR6tpw
sc6AaAwZpY74wPxMYMyIXt6HCSQmECtU10KF6NvyWwt7dtLWvzyi6fs/9yfT
88XwX+PjkPYWhAJ0PRMJLYnf9K0DdoDzK45kuvPpxriBVuFFEH54BYEumDSD
PaV3NdPoTFQps6C/91ShAw0Pbzk3LpA+bAHKJt6uepZLXoRASRT4J6oTzXhs
cXPB/1KUm44YkX3Rv/HjT46R3YDgVa1CBLcV8zd2LjNZaJfQmkrbcjv3aelt
9WqfVBGbxpsJdLxJ1uqdxp5Zjd2NKfw9QHG7kZknmDwzJgq3Zly1ZOB7jP+J
s/+6kAMMiDgZ4FF4NMWz8T4J/i6KX8Llbj2sDUp3ScaFQ9/sEk2x8B4/c6mp
Vo6sxK1+IRRM3ZqnVozfiCQF7SiymekXkVCaGnHw6/fxTr7RLeTTgIAbVfUN
WbwF8FBoDhnTlddo1/XLtHVmAfyZWYqWYh2uWCthps47A/k6VF1SuaZ6TQZR
t7OtpqfI6SzPfsD/IVFz6oHrsuxK4+PxrZ2On023zuqJFI7GxWR1eGNdJA4M
ekazB5ilZjNncNv3GW+WG++Q3dY87FRACYCdGQz6r4VT9dLjp4DUXGvoLt4L
zxB9JpfKuLBeTyRCUQvavokkpzkaOFLvhzcPkkM9hGDoH+MBTUNszIYw45aL
CV5xljU42F8S+emyEXSaJvl/2vuXY7LJYowk2a2JUEsrIbeAQEXq2eThYKMM
JocZ4GlCwUZEHA6RD6ch0dDCU4iPgm7AjevJYqftr832F9XtASL6yfgPAb0Q
+0zeTt9C+8DICbc0ZPr4gGqL3RBvmdI3Xfi5NB6FDuSR7+54rROesJyeZ/u1
1ltq3rlxE/bI7mpDSS+Qcji3/JwqIoZYNw4+PMIw2FDl9mMsb4tqpFkbHzZF
IBbK4MByQm6Vy3bv/tjH/1xPoKUihC6ewT3IKmC/g4nB2MXT1q9M2/pnog7z
T2NBSs7dbXEyjZHMZ52cGO/2XGM9NwQVjS2YNw/gbB0UPhScadFKJLoVfZTU
AA4pjAkZQpdUmqorzsAI833Yde7pQemgJc32d4LxphnKxtGybaIg5+ZPw65q
2ZbWpA7JPBH/7npOzTis8u6D/h/DwnjEb/LDCmlqA8wnk45WxGXnq+XZfSv9
SXGVIsG2vEZcmLMg2KIHMVhQC3TqhQnmBm0Z3DucVxhqqVnOxWwhoO4KAojB
WEvsChbjfc7AUxZneihrmWK09chmORBLoIXPZHAjiqOYbodIW3ejmr1EnPG+
L3WIo3k2/m0WcxH9NXPsng45l0bzjMftV64O95tJGF2pT95dX8PKnekIBbQN
RUuIE5cEVJmdvd8SfhCizHSz1vBON4F3XC5nOWuGJngaGzIlZH5OCCu2RuFG
hN6TK/eb1N+kgB5s11Fp8Zb2sr6AhRgK5K8/G7S1AyVZDgY0ItK+E4lrCv81
Sk6TdGRuFr65j/3ZqCCDSG+uDDcrLT/qdyfPK9pZZ6pdb3gjX0Z8JEwkTS8a
tYyouXmjwodwhNFLyQDDB8cb1xD7RHRd50xocLh3G5KccuqF20cwNs8RGYQ6
Jj5Kntm3XHrxiGK1v6Hvp+/ZAuy7WnFjaMDURDiUaxARtlz8V+lFIbs1tRwj
lRbKr89CdfPdorSDatqMwcpxcD6mUecSlTh0A9lfik1zIhdTUrSN0yInlgqv
0ttewsTiGJdNN6kUn56zmyczP5VESZW11P83dRjqokSGonMaCdUgxMV508lz
HdRmu6oHbPmT4L7Dj1/QAzHXr5+hJdaWuL7El2sXEME0FAKoBXY3CR0c2+Y+
SGvCGKmCB79nJJvKQdRSjDq/Wsab6Icln/G3xQRmsodI/lwQdtysy0MCrOPS
7RaUDcfU9WVCRbwg3YOIgBP1zIHoyGERo53RDOdEvPa8xrHlGJ9nsYgrhYaT
nxlHrpfPgg+G5A8bCsEHCcD01y9NyJCo+JoiojSXJGcfNkMqTsZHu1CqC44K
2hPQxeSYnCUWafYTRncIgOryDqYzby12uJeL5CiHRdyVqbtTpjTFPRGLyB53
+NgspGHnRM2aIev49opBjAGdYj2f2SfMwVWHMy+U3oULCYa2IGOHBlW76lI9
joKdvjV/Im6/8rW5efDLdZ1mxlOtgJkd/8Q104r8gWCMbbI+uqDH/81WdnRO
nR1MYUmF3KGjD0aUg5oDlyyZRSrg2Iqit1sOK0uMBbhdVrIzKi8rULjJLG8i
FQ41y5zyeGTJbDouWU2KyAfmDrxFlfPy1her8NhuOLXZj7wDO0/uIE8VyjNU
cZSFKjIFs/Okr5Y6PN+Auo6IJlH8c0ryUvQt5lprNvPrru/VjbXq9HMQl9wz
qkqdu+uS9QxuBA2IItkZxWH7o5F4e5QimT4eVAc1nP4NAMOWwwRaTRT+sBGo
2by7ZtCcozk7oVHDvsfAXaDWro6mY3dD/ADoBmJ6tl0abOjRoeX7TM/AHP3U
K7YB+lBD8aUnv4zX92kkdPZMmrIkw3g5qMrt9pHxiwHRjm7wszfIiR+uAlRz
tQDATmikyRHcTiK3C0sbLhVzI9TsCGeSQjZsAyvBnrUVW8yVg3h+s9LqR/JE
wvhamTSM8N7hg9m7FG0h8WNapuezJJifgE4lTBdmvobOW7mr+usLg1afFcFU
+cyY3edzqCOgnLby7J0npNAVC8ylbl2Ok4GLoVAABQetnl1Tp0NxZS4J+pFn
baqb5rR9HPYQrWRpHd//3rDP71w6xlFhkgOAqNMyWPDEs9USK88DQJr0qua1
ezn01oiMGxccOQlnkx/1ODCqHxL+qGnp3qEa0JxJZROQ5Db1MsrWtLR6jgxq
ydVfVJNL+OT0h/VwIjEE/klZRYHxUqkifJ69ExGSCfmJa8G0v1bscl0Xp9gc
mCnwyAVBsj7WmeqsMYLRtYdeHKhIU5+Jex2A2/aW3ribwdA8TVyfKNOzLUWU
/RuSbE3df78VpczOtrv57gKv+4WsNl6QMxrJ68RBkV4lvjbgkWcwT9vytHUZ
4udU3WJP2P/eIY5HB4QlczizLTCdUHRysXZks1Mg+Oj/qS9e8thvw6LHFSgX
HliS7MAQTZcY9AELowjKe2/Uq6JynVn6YInm6qmbv0E6rgm4xQvUfGxCJkzC
TQ4mDtZDMVolJdhzDLJ6w0fYOu2wEJDrsxLr7hRR2kuWpFpvxhj/0kWumXGJ
Ez+hCk0LO1EdposXxKtCKXBKkUagp78ceejX4IBlRqpiPzVQAFNwut8V/xxk
lQlWQcfZh+/Z5AMTprf5i43QmNeKIqcH8e2C/ZgAS9PN+egsJxLZrM/L3RbX
pTW5GxvfFTjnycvrGsCPvze92p1M4AAFXy1vJa5pSg4Jj55Gh7FxMjcEwuat
n7j+S/68x6DMuk77C4FgydoLE5OiXOM+duJgA1FUXjo9KjY/LLPb4wup3HqN
QH+1BZn4SwxH5Ole84Fh0dsA1YYuVV+Rdrxhx6H4q4YF8xFR4yE2sraIfwcJ
86fFkNoQXqiBuoHa0VMJgici1+bvBPgXRIsDmzcY8sAjTrX381yRwM23q1bH
A9seOa0CoemmJf8zf1Tj9jVshBzGwrcEXUH9grbH9LE5WiHJYqXHYdW699Ks
77+Mm2wFjdc7ozhso+XPIDofxklM+ow2pp4z1ws7Eql5I2ITb4hBA0CqPNoX
znuZ8+S0aFfyaX1b3iRE71N9Uf8oqpknI1kIShl6lthyq1IzLvYr7/823Z0R
OTWQZ6SQi3dv2i40iVIobhk3EkhqDH/etdzqquWvXF1FPnNqnqY2vqGgp5xs
r060vWNkL9YGu2uYaK07lJKdAeV8nYGj2a9XvJIhshX8Y+qhYopZQzZukgLC
Gs3Zto69pxe08v+QgNN2vOVXUbE94ptJfSqrIyLiVXNBGuYqDXxKBn5TlQAv
3Mwe0NGOQXvecRrFoIUoQi9yAS1Zc/RIJyq+JGGvyxxpDURGmskB+uo2/WUD
56JCpGNMLTdL6k+CE6ooYzXP31FQtWwRLBs7r4T148b3gQXq2b8XslTojEh8
ZyPBgLWkTFhEjxCAGSxA9W/BHLLumtjM4fO0rt29qMHbsb3xOFlK/XoqJ8Ec
Evm9FJ1dXFtUoAVVk5vQkFjO5sGEl77JDFrJ07RugojfJCfb5ip5adr72LIN
/rXDghxShgeWW6zFbi5qBgHjwRPzNlB8YvYNMeMkphgCS1TTBQvikk9yvFIN
p+8BHaECIKcFXGChpo9lmLxkMv6bS1p35bsa/WaNlwF4FDLO6VPnab2X4/KI
cXWETDAohKxN2kZUAQE7VAsyTBN242QsP67dBZRC85cxMJJnuVQA47Qps8wy
GweyOGkczKH8e2mgGhas32fG7f5Axo1+F5QhIRClX2tt20O/2i5Qpa/Kphre
NC2kPys5akRTAEHjnynLmbwdrs1IxFlqCiWVXfITVhp8muFKuQMwOXCzhoLE
G5M2jxy8IEsPB+EUPvIkkEEPst0d63SDERVdRQze1Wjle1VsHafCCestTTT+
Az5edUTJNJEkDREZEoLcm8FfsYHzPmxDABUyJgooXY4RFtBjPLGLKMzBJKxJ
mvs4vYHu694EesBK0Q3wDO4LXzm7pmcBwwi7/brWdPS5K+V4iyaRH7hhiVqQ
1gfSfmkGKqGUTdyNJjrWmazcGmMLUdex+o9sc0w85qnN2KY/BmaRzPCR2JX/
EA6zbzDt9zx/+iFh2PeUYsBBl841BxqKB0Kf0yhkA1hSah2WogIntXZc15Dw
3paPrExyCohpOCalWQ0dxmqLmu5Ms0cI6LrQeFyz9nWiYjXVr9/2cfmDThPB
v5wfM1Rxc8DVBSLTSv819gc8KuIlhh9JZf8hXz9ibMCjmEYW7FVXdVKRoqWg
E0drVAo+8hHXpajw6dctcEclzou8DNdJIbbdsdFdKGOz7LI5eIQBhjxZBocF
OGiQW2UjSxpBzVVdpRvqBiA5MLx0+I6/LQv/ZpL7Vhahz/pIIurHQIHMvGjH
7grKJT5YBd+X2vBrf/Qk7C/OTXCl6bWgcy0fIgkPhTouOuEXnY+qvMF090hg
L9+bSc457ri1c97GDm0r0eebEkkEGLLqp1nnvh49+lR3kQK1P2Au5o2MEAbi
KErmNugDj99epyaEYp3Iw2Nc+nmwocOeOhv/ZVkLorYMyEZqFS9DB07Ao5Iu
scK85r0fqkpv5CYuTgzURrS6sRi6c2lycb8/isVV+yuNorcUItuS12XebU/i
sooVtGMQf31n0XJ3FL+0nBQoNXvxAnHSkX3SnG9MPLDWgNtN9qvho671EqPH
AvA41Kf0Jvf2nQ1zTLyq5xyrYsej9Jq2GRzI77komVoZOK7EQMRiTfFPuWHs
Ed08AXWsxx2J0Znhfl3AnCodzbG51DewSE53DX0tHpVdelL5vpHbC0ZttsRk
U8rKHAAWHY0CPbRP8+J8f0kIqLR6VWlc+a800pILDvS+o7nAN5ufKNHRWnKq
oJSbR5x6ACUDqRvVwITnOtOYKvDlvd6fNFZk3udQSM48avR/j2nirWKqN4VA
yq+/tA9W+vWB+HUnHsCx1mO2pKdzUkk847yPzNXuueBGNRvrcv5DRjid4Mwm
yYKUEbMr5GRgao71gIhj+VVav+OW0tSJw0P2QydXizDQmiNsweoBhXVETULw
dpJdeUoHVcZWfpm4RiFEENt+ZeKoRxQf9MtUKCN6wGS6fZvunJCZ9tswR3bS
Np61b+h5z/jSpbfX+JbnIGbbBm7svtvlqAKZocnwvh+XdFMzSfzmteF0ivvU
C72rz1HvGlrjAL7VfE2y4/4jkeOVgidvuEHZfsODcPDtn/4lWDulMc2zDQtl
sG5PuGw1nVVvB8MgaATu0emebRL/fmo61YUGPD1ZqC0XbCTZ0/zz5xZuFL0+
wTlM3h7ExcYHFh4Datzd3Nv5e66NrFV+3b9TkKKO53BloRbNnwtMCqia7l4+
d9H0YcMvJyfr/zMna/fHrFOJxoD02WTVxj+9SF6jj4oy8atkELZh4oryyFdc
9dl8eUBonQteosGyq2NI0wSwI+R9WGRGl4tFnuRlxgE6g4iWZg1glNFdiU+h
jBiyxIjuozgg5tP3kb9DKbXihdmcber6ItNbDA4Cw83UDRcIDGcE+v/V0yeQ
UI+Zzf77GmJRhY4VC+EgnFbEv95gJB5KpIpAkGPJXs5d394BSVugRU2wJH+z
PbO3cAbHDEqUlLNL/6zvvKBYnzlmlrrTS1SI98J0qR5bWbCNPuAlAV20KV83
H3z7HMutop8RQ+Xi8E+w+lsoT+D7/zn4wt8Id5yGrG+B0WudBw0knHL0CpoC
NkahBoLPEl+6jbQbPyRJVeapfGvArJdwpGQBivapFqc6gTPZ9AGCrd0TmaOL
T1ib7/Az8BTlqNny95HJBmZ/SEfbrd3KvOLNBG0y0txTvPZ8UZGqfejKkKtB
RR8rNjquHloDk5iNU1SiCV8zQ5J1rnVWfmbe8qHRHyfuhg1BvPB2sFQ5u0Ky
yfSOz5jUMD97gEtaU2Mvpv1ijsSZtOvmkE7ApQNzt7Ps7xL1ZMCV/Qb5sb96
TakKxoNwANjEmsFruIu/xdFXiczUUeFauq2anijJsMwFr5rLEl+bCECwiphG
2q8amdYUmnQLMHdPS+xL2l3E2k0c0snb8F+sN94Rjb0zWM3RTNJMcWvZFJ7E
yLGd3ev4gGlA46fK/VlUdniR10sv84xIftzrmsNlG3rOEYGI8dN/4bwdDBgo
MEtT2c4SLYmZD46D3L617clcMOGsFOLyRlDygC/kECwyPGcg5iCQ14d/XUKU
2DWqj/5Ljq0XojuQZPdBSlxEc1HrdtTIky0e+x97Yhjwj3FUvzCYq81Intgq
AOLrtFiNY38mMnuNh5mpVYlm/lMAuJtwyhTpk0ddyznHuy4k4y38oCmOVekj
/H6xFiDcJ6SYxmQNSoGCRf0WW6TsOYJQuGYr3de9EuzjP7tP7Pp7lYsPsazR
9ypzqp1hiwTNm8qfej/igqKSGnfdEdTtGsRoH418GElWd/CgFvpsnmZGBBJ5
xIi1HCU6+le+ac+RyN+4QhoWiQdgmMruyaTTwAz9bHD15uUb6kYCu95AoKzT
nNpKGuVzqY0kPSPNxJqgt8On1ds1S2nQbbyT/VaC+zZ17VRWnUHPhuYikP8x
LNcPWptIbsmM98tgfPHfP/oA12/eiQHerR3a6d+GM1hSE7t2JAGwO73ZgeJn
2lsHldGykXWoUsVOhRchSO04PuRCMlyLeONT1FCycX9SshrZjtOISlTrbKsy
UC42OZL8d9fo75dmUrcXjQ2echVNyAyYC7ehrkGF24xcK2Fe8Quc3fFp/xd0
xmhJtZn5aV0vV+1r/TPWyhfJSebDvsQibxAuYp5jum0/kVMFzZncovAxuRBJ
qzFwfH63XVLLR/rjLtcj3pm7FGLbIuKkwh4PGevVVraPuQ0ST+JsDOE+o4eo
n61Z7kAlUCY7lP6HxCPkqgkPSR2Wbl+IpUPZR6GjwjDcNDMdmWdxS6PTVjyV
3UYmhJtkd/u+MX0houn8WSPaQkud0GQPgKq5OEI3HGNFgjmOpXYGrBa/WuVG
xpCW5zJuopl7hbzk3jSernz8fDa0opj+PzKsih1F/5zSYBV6Zsz5nje02Vm9
tzVrfj7oTyeyUKGWMDGhEC3XH2Enep3Q6G+ZwJT0vCPh60zb44n9CkKzn+Eh
50O8FYF9tYdic4oV6M1SgOdujMtiU7c2aqJy1OR1Pn5lvqi2mHOk0tNocnZV
woE+dx2hAGEE2QjWXl0zJ9oc2Ev8dVANmAjfQfCXAl8yMulmonPlhmXciV3B
oF0EJS8dKaMcejEVH5z+orP5okyx5z2kemWekZB/bh3lHdGHTH6YbwzDKyVt
4JW2QRTldyafDhn4oKqn2VLapTy2mYI4A9GPszkwjStW1uIhRv3ZowyVNFCp
92h0xaboX33ov3Z5HqXuErCvoDjJJ/WJrf6G0fR8c5jP31sM2HR92w7KIoCf
NBgPSkeSdv+5yDSvmGLS/ttqSK/6WFRFmuoTc5R+8825+bZF05Hlk+L/zivY
jpDJJxcWu8Sm8gXuzWFGwQRGQMjeaI8lRPnjrndHFeGbuYpKbjtVenB3wxg3
HZr/CkxZgcr9mY/JFNPqYv0VvA5rW9fV4P0FEQ/lcRH9OibO98hMgsd9BeWJ
0g98JXyZk83J7cL8KzUkYH/WhPyOxwLwHhK6PNJbSmWxi22zZpow9J0OJhtl
3eJsfr4dZla9/zEKPigJM6UHUyxrvW9MZMM45N7RoQs6qgHbzZIv/F8BuMlo
uWOK7p+Fm4bpo7yOdyc81lvPHsdjK9iMlXS2UdJdWQ6faW9FBTfX9uEGHwJ7
UdJY0KRGuWKyynNa82sGnBLdw6xgI9Sr9Ry0I4vzpK8OuQ8NUYr47t5ievY6
NI/2t/f8E0pIGMpjLa379y2L88gFdllVGlXyaYIC39f6VJ9c53ZInEQxeEKG
8MLJBwM1iDgDEv7hqykz7YwagvDmjW4giXu0sOLfFSVfugeHU9h87+ycrk1A
P75xVshDha8s2nMOYCsK8nOGgCyT/inOskIL1JOmgB4+CUNPgycpc/TIjN3n
QxwMtUcJdddiwIqGSGBBuJ9ond9Kz9wxIXGO+2DSLdMrFQaKS1iTd2jc1KTd
dB0NYGj8cNZYDJWkDSO2Ser/Xg04oq1CH1EQ48K/pL3uAzQrP5XfRVkiZ0Ih
A6O9TEJ0wwV0MRXcGWw4geO49Jey7CdLfd+IKeg72DF+IhkZQUVQ30W9IEQJ
bpfzDfzMdisNWKf1UaZU9yevNfjRoTVkrJXuz64Ml1hWEMY5SOq4PJoe9QlB
Ity7dDw0yKjjjMOwrDWWrOGsTOZ1TOKnKXvnKcq2tIVYxvzMggUHn2ht9/7p
QPppUIcGTttZ3+52o9i4Y8FhHrg4n0klvB0JFAfW1s72QH1BgxHPIUpDFPvw
vzVRPrmEaUmCfAmyruu2jqAkbS1b7+nqBqEQBIDvMrN3V07RJgxKsKTAZFtf
oDQW+BrHqe5jDPBdHnwcwwvFLdS8QOEzpLiunJuBOOpGQmuCr1eUbWElM7SO
g0//kaCs7+MFfdFQfBfIN4la8XF2l3dN7bNla3WouQCnQL7G2gU9+eADs3h/
O2dCyW1tcZH1bOrmmtKtFVlhYHS9JLhaFvLwNbMmztk+imxw4O8Bj+pZcKE8
8sx1P+z42sI+ajJS6v2mlWpDAFs+cKKv5YrCN3usDf94xNEaw3UfGLTnOJxW
u0KfFHwtzzvDS6f+srdArPuYJwOUOEshQ4ZR3HtTf3dOc3yQIyeugaITbca+
JWQM4rK8gGuqWlt4IDjCdvEDqtTV5eLhrBYqA8T8xg4IpFo/x+eSr0QZsuEr
U0NAtAckCXEwKbOW3vAD4BNXNboGYjIXAhdUUfN0hhOSZAnYEjfTZOsPQ3B2
jWrbctqHY0Eblf1wrk40YFvkCOP7rYTGT4T38g4gpOn8iDLUSUSdIEbaEgHX
ZWPJ15smRntt8P9+uCfH5I1KkHaFg323iA7Rp1suZaqBVvXMUAnr9HaWdIVO
4YZ1NscBKcM5blYui4xffJEluE5Fq13CmP3kdzMD2d7EmwVcEfistLvhARUp
GL5Zg5RGS62j+gJ800+tPET0OWQJQQLChk8Y2WfKH+yK8hg6Dj4+CTr9BsPs
m5IW9G+gBuk+Jpw951aoUOfUY2hZ5w68uqunf0MTXhef151Lof1LMl+Dl4I6
B6Wzv+pwMD3DbKUahwOKCFvra8ej0mSNS9XjJNgzLydb0scxB7zOvlmirJ1N
xMSg3ItRX777ndo/0/ZkiGWjmQrNjU0YY0vm5xwta5WgociuHUJUhSJJiDJT
TlKlyjqi3FwpELOBPKMHG5/UUUSXOVoym97+GvMmm4S2QI0dRfD2SfrihNdt
qtBeVLHq5mXJStWHdSdi9NRQgmWBeJSH7n2MtrkNrKa9qOzaUQKomAZHCwh0
uL4sPZffykZk/Hc1c2tTx0pbgvjBf8JQktGtDqJS4Vite7Tui9Qrjz5ap/jx
Bo20Mh6kUKjXUU11d2dZMhaVOYk9jfu+x0bn8ndPG/iEGXHTb5sPJxW71BUn
4BfGI8syCs7RyCeJbzJvw72BYPNY/HHWypiGsWfnrzm2wSGJPqSi7/8PqTP4
WUnQJQYfYYbrxZOk/8xC/mLcXzxoVha7zS7/V5M83qD+x1VHdJEpUrWIW8az
ckX3NkBf2xAVoIRI9EyLMvNcdXv49nCQt0Ig7T+R3yLhTlTs072W7XEdNVQB
g70fHwfcLEujE3HjaDQVhyryGVD105Axg6m5O8ZJObGwKY467bQLtwFC5xbe
8AS5mqcjCLMH5nNy/Xmlz0oWOskxcvTgThaFGM7dTx2zGLW5g9r6Z83Yrfbb
/yL5cAZcwbafdv/6R3Z2zVQLIpAPGMpmTwaEgfrEmnjOz61FBkW0VxeSuPf2
YNzbCMnbJSKTqLpeOKUZSf+sIbURf6LSiOk4kxjy+wk4a4qNSMayvJL1TbBT
y2Lq1qvAGjVGjknSJyJLqZE7ODka0Yarn9oKAv+bDW9zvdcxJhTNBVini/VU
WiDXx1L3C97aSA6ffix31Essakm/+FfGf/BySqq7go2UR2AvkW7tBrARN0nI
Z/pKs2ux/eeYkkV6zXuI2TcUUOu1OJ5UVpW607BBEQTBg+2wPuNWeOPnmgjM
ffAp05V7g2JLfySZdecOrM/AySLq3PndbM1rOSB/LLXAkVIci7mfWeeJNRTE
FHoCwo3R2TY8E+zqkevmHLyf8mxrt0QfMrvoOFVKLUqm9mP9WiFe0yoMf/SE
F20zgR4o/mnDl58QdXlPnQLkJ/1U0A7TpOSCk1ojGv/8m4XD3oZtWjtGHLgw
6+FClJfWVC8YqgweSgATETwkfjx7E/zX0JfaBXM/v62k+ZY2SBXFcL1wG+Ft
4qOks9y59C2z3y07Y4i1/wf5LZCovGk10GXjjf7QqwuKmsDDIJx567sONlvJ
6tLVDtNXu0qCyd70jFIAhshl9LOZdD0qWQmR5QsmKoSGcpr4RrTQ1I6s9Woo
WNjGpkotBFxJENgLit0SwqE7XCYWWPfNVgv+eLxVpWKIswm35qV7txQvJcC+
0hm1DYfk6MA/diPBkyZ6ZNGUyG6koj3XRvk/6h7cS7bR7Z+1pbHWHykoQN9q
+f5pSIUVznln5Kr9pdgnfz1dgkoxDVi7OXpJtG2FW32dS6Oc5OT2qr+LxMWb
flZ15xrfgxyxKAnvk8N3mtB7nZ09MsZZd5WU34RSYZrz6Vtf6RJcKnb+tx0u
XA30qFymAoSoF0wjhRToA0ZpHdrvghSLfygLcFfE7os10UO4b4Fgtivy4zjN
ETIqH+S3yEe+NSxYvpqOtybh3cXs9K12r1EJxEvhkbF9/TiDq4p7KYEbYwsg
CyQzC0qlEq1q4qKiM3LtT6l55NCDADmYPmWzKnwj+/5WavwB9Nqjh5nIOXCc
6A0vE44QYBjZowqR7XrOKH6lL/P5PaoNvwor2jnF3wNZsucDI3NiZbLTzKOg
CS6f4nJY5KD4OR/W7TFQAivQ7PZy41LpnrPNkZ5ilAht2CSVd7QtLhk86k1j
fsXk0RB1XdXOi7isq5sgsct4tqBic1WiQHylNMN66x9vIQ5VssQpibqLvK4i
bTtaiiCGB7LRKlTJynFnX+cW1rZ9rfqqzdBY4l8vS78jMcno2FqiPFBVIOEb
K/0rXbsXYW5G3UMaiNYuO1+Bt9/RR79Z2g4893Q3uRsyQyjviWyRjC9szHYp
q0+5gXf13zmnNR98mqbj/7OJDSPxpF5qnwFqDy55WuWHB9bZ0XVsZu4MLts7
KFZHRx+1UBuPma2LkJZl/XNxGbco3Tv2Uwc/aT53hW4JrvMk1Ppv8a7t/jQE
jaQUP0+2b/uA/P7hYyzY1OFb1z+4O8FCgm9xS+kfGziIn9wz2NIPFO7nYiJb
IczRIemzTS7zKOkvEcX6+4NFEI3d0uUfhVRbu4BHSzcT8uSAiGk4lgNg1iIC
/x8eAblGl+aGF/nFydDWCKk0sj1QSewTZdaYdx0ljZB0Of2mQ6HM+qnHjiiZ
uIVs/wqeYOX0F2H7nE5zYp8aak3CH8BK7CUSy1IcvGYIXUwtfC7TztnrpCfY
8ODkumz47S3WVoFVuZ7Xo0cbZeaaSRpsa1sMr3YQ8Mgw2PzT3jOypI7fcOPj
NdvyUMdyw2hU647bL8EPFNhh7IOBfsiwk5ATJ/HKPlIHzPbojPXOPvVYlGXy
+9i4/RjumfQyJzt76TdzGX/AXLul02AyHt+tZuVDLKu1TxeGS9a4Cntvut6G
K1biAIVouUBHrpHgZRlzuWQL5leg3zO6PhuPuDLHUg7psNSyR87pjMDUOyKL
MqhY3Qs8DAeWhJBPxUXhTKo+7SKwfjYMQUnRu+lix0yTmoqWfv3saowWW1JB
gMZ66Sn365N6ErPV1iw9oTt9pqdlTQKkxvQz1XQkPVo1lQwm1xwq/Ngodr9D
Z1C6rVHxh3bZza2rsiOdHBMzB8A7D61pESmcqy53EvhsLU6F3KsLSThZneTs
pTMgnlD5u0Ey3uDiXOIstJ/T8e15w10v/Cotu4EsiNE3POt1zJ9y3UI9H+4/
wFSX6fyS2c/KA/rPLkLieofXdmq+AJH5+Gai82c+q+JWYoLZnhG9h4ttouQn
sRsNkjftL+9mEECUA03HMWLOqhWzAKu91VcK1CNfFE2jHb6Wf1arIPNHVkjs
onX6NM1p8uSpOwBONH6mZ85NJjqLKb+oTovToAdmrkA39WOjQZmPY4Mb+HqI
gWquBy4hjpwLZsUy7jn05X8gGzQ2SgrybYDl4HvW7+fCxTgtXdcrvrI53ALh
eH1OHLMZnuVav3RQ1+PQORY/blxVwpsEYXm74GCYuf3ZjPxoiy6qZEfgp8aJ
6RhTI3/joJHBlXTnr8+rffBZ2JBDBOitqEQtjTxqYvzjztFHoFcG2ZdRfCQz
1X7RD6acwXUUW8U/cWxffHmjpgcOk+/6u9lBSlprB0W6shku3lA059Rt8P+7
VGevkhcyDbekvRdp/3AnZfoBEHzm+OFNWTMQqIjC3/V4KTcPzqFruJrryGjx
gwqpGVWIZkPvSYofQggLgmvVhTg1LU3acn9YQdSQ610yxSig1wZzkar3VVjt
sFaqsEEGteHh1rCulYR0L9WrCe31ANN6vTK/B2T0FZtimuZgKkhj1W581l0z
zlPpVLWtwOnbl1hQ4MfjS7gn0swy8jlwhCFLiWjXl1wvK06fO/mMyg10ed2D
i1euJi0tV/c30uZDvQfl9arcNZelbvUbY+vw8UNZWpMLRHh8qnXCCO6eumyk
cUTMcs/XPfrydQvK1+C/1Td2yyJwNdeT/O929XgWy6YZ2P3yZhbjZAGW0d1p
K8dNxNj//1d5a87rAtYmVJbETkPqXB2xKXYM5J6G7ZxTG9SD1DprB+SU24iS
5eqjy5x2fWGvyZKJOVeL80XAygoc1ulndeRun6++lHFz4Fuop4g0IgVhLKZK
aikMEgsa0VDnXRqiuzLLOLN+cSYAt6naPuJqsmPUNmKwOr8tPcBLFnPM9X1Z
/N65oJQMe67drinMHKk8h5q063X42P9w6pb2cN2YqxOP4jwnvWfhyqliDHnK
ery0koEKQYuXycjYpBBurX/dond4BbbujpoOYk98J1AtKiz0pk3X9NJVqSZR
5V+oIT0Vr3DalPdsw7sXFYvVrfUrKit8fqjYqOjyfnC+Cd8/i2oXta8ZOMSu
x8Vnjt1XhP2A/xgwO3SAdoTSd7g6Z1F891pOizEONylDbh3OzdXFrtzeu+nS
zGpmf5aUSxeznpt8ik9dG16X207RpXQtWkF95o41hbu27Xlw/YO8DqJ0513o
pGbQuSraLVRrJbd4xtayTkm2HfaKLW8gFeKxcnkC8XB3+qZ/z6fUasisEBNs
lO7hHI/lDzyEUHAipl5+Y5QAl7ChZnmm7m6XLHz4smcLEuXrijw+V1JxJ5Cp
CLLu/LQLeUlx7jK32FHUoEYMXwkpeKZvHfKZNXz1kSK5w5gTD9Oy4F24urjI
Qk33GpCfXDyrg8JxXIp1Mes9PxYXNptm/8IcEmiJ4+mxhXCRhbBvfj2qoIvP
aHLAeeZpd3K3+BQ15g1EJo4Jz7MtshvmFe9PlxpuLLJPsiNXjFzpWsyAtTm2
5bbu66aH83M85FmikOW0RpLq73Dyfp1ufAQxTw/OJZksxVc6gLLiyBAypcva
Qb/y0xrqV/V1PvBtU+vMi7bVI23UJLg2vkUzdrWnpLMaFc1kvHUSGMVwWqcM
Mi2Umud9HvTWK2q3d3Ce6ZwUN1WNaM+yHQKzeIKXz8LS0ZxrQwwSb8sLOL23
XDg55TVD6L4PhRpAZyPdNTT7P7yUYQH5h6PnPIjcLLmBknh56aDmpQZl2hUZ
P0MN+einCMO00xXZkQg3SNjMa9e/iwEQ+dbHz+kKe+VjiGBVvWlRlvzbk/BU
bBiJ34Pbvvr7H8BSzb8mb/fm2uZ3rnXmmb4wsTYOmHwE6R+Nz04p8kQwrjVq
wTfu5H9jzSWc+QLQkpedCP53VU2gKxuOoAunqjcSVROfjG+IVmGyej5HsXsl
ziLwHIJv5JrK+S/uH90bjdh4avJhYXdAVBMKyyMGR86q5ogFRCOp6UyU22li
gXp4yyoqxZFqugsBxwzmdrdqkLRtUQZrpZIH4gSrwLVJ75tfS4+XZQyePMbJ
vBo0R0VNZ4+53fnfEJP2lQffDUvMVe+7r4rP+oiHmo+TeBKhe5WDdMQ+slvF
2yTg8ULH3qEb15r9isJyQYYvCPXD391He+37fn7d57gRuM+S5ZDHyNW4OsDm
NxZUZkmZCEXMDVGtOkBIKDbse61muC0fMGnLkcwZ817L5ZvScgQzViJIBFEC
dkg3tpGAjIjRlYbgGJxknahkfw0zEHnKI+okbAH1dCQc2fClrWjnUaGZcYtB
bT+vATubGWbV/I9Mem6rBVKNTtLZYv2iSPkm0wlhTu+/i/RpfSOs4CDoKI77
eq/h1VCFMXH7jwI6tfFiXnL0B3rlJ8nILFSy4T12BOUi2lRpp7MZkmeEQyW1
l1hPOG2w1kzXEsXTy6//kG5eoDebH5hf/J2J+8JBI755vG2UFCa+tBwqQXDY
WkmifROlgT2qn8BS5ZZ5p2bLWumswEA/HDuZjdqbXHoHZ5oLCR29IF8MF5NM
ZQqhrRHoPihdOSG1OzeyEX9ToVNuO0Wj7fl82bykglv5VnMrm/O6zEmZwuMU
9UhwBQmcLvohUEgCKxUp2ypKD3am/aoSokeuk1yztyDKoRYEE7O24hARGNPP
LN+2HKNvT4PXgu9VIRRY9+j6KKbzxF15cyYUm7leGEXB3M8IGMz6v6Ex6FmJ
9cVd0ImHc3acIEV3GT8pv83l6WjtsIr4inrmsCFQ65EQaRAeFB2WChE1Ii6J
rT4LPdzrps+BEuG0ys8PKupHNooT04f3nyZklFpG7bpUtMLupNDe6T7qizDK
XCJ1evo1ibce1qD8ha4U4tIWDPOQ5AbpAAyFmiOIcYI5QEDTZK0Ly6kh6p+s
MG2sxXkWoKaAqBqHcNxa3tf9DC8vHtR8+LAUnuUYOwlwXA7/3IISaLn8hFKW
izfGSWTfCmArdVqYQr8LtFNiSSJ4DwAsC5ut8oUMnBVl2vMWFbvk0YhzM2iG
gYMHukTHvYlmgYxIBhOo0FrY2ga+5NeMeGRhUnW9KTsH8eO+1R7YsXzFBXb1
8Bc3NbGmY3sc5d1DHumhdAXLQXa/8GHExlOXdFZ0O0kcG5XIKSRd+H610zk9
HCA1GZ/JfIK+I3G8IuQBvua17q/Tf3lMjoi6dt72BvkEYvOW4Ty8/8hRGQCv
Vw2CNt03IRLAI1r9/wWYjHDb3N49+8BJR8QPMkBFhn3bDqJXgAAIhTBvOhH1
67yTxCJWOwpIaq0726px9AkQURluU8uTf9P77aN72TjUScMvbcpGK92l52Du
KriFray9cDAJVcnDUc57JjdCDA5AftIbQGgFVnOEEQPy2c/CuXpZbFjRjcHb
PorjMlIUM4mjJP5bVL27zIJiGcKahF62yE1SmFzjMv9mJt3b+DJdtXBmvchF
7Vt1nNjI2VZLuFTHwCo1z8i7N2sZYKGOlAtDMUWdXRjheFLzh3v7xCKmgviJ
wwvy6bOpMsXZn3uIImb4bIocSnK0gK+HGsEVAujqjhf7uT6uHUPXPTFHyYx6
NpU1R13AsDqD2zyWm9p3hivznCf29xmOgDS1eTAm6w3z4khVwJdO6VUrxXRM
rryocGrFL5FJ+9dl+9XIB14te9d4vVuDjeA8KcWvlR//USGxjfUzGeVBLEbD
2UPh51fZjgSDLqJK+ePOp9TCLlNgxd60R2SrLY+GRXkEC489QYSEcgFOvZY3
BMiCfOFywSCFGV5g+1DtaB0AwNFZDOU7eCc3zkLCZo5DxZGDe5bdwW/E4BXB
SUApR4k/E14K52YQo0K4wU3oQIy32zChnEoc2hILUO2yk8OS+pT6cebSDYJq
ygvzUhojrhZVefq5kvlkBtHNbILxJiZ9vdrydVtNQRaY5BSdyqoBi01zBZgd
IrLiX+wz47XRyRjB87kXktEhJarYYYmFtywzWrgWBqrPtKT4SFNQqLh0EGmw
wppkJhk7V2ivrgRvdfIJ81lk2kojoNGE2Y/qCG+7T7YDRjqKnw1vqJ/sSYgW
FSq7QhY8NfkeuV6dQ19TY0x54/q4XtizLvMgqk713lvjWoAlF+ZWRbB93Dc/
x02vMX9d936Es+It/ZQyI5GuflcfkPAFk/Rsxd2As6Mhi2MM4wWuxIds3Sn7
WqgsGTls44jd+doJ8KSgXxkgjIYdFJy7oRjmHEx3Aw5bZgXttvvIX6lJDy7J
PxbmvEnupwRaA1Ts2FQ1EZ6QezO+4+FzCgyKbRmZvC9MBGuGtIOCkt/kOMc7
v+NY/tvsvILy4cca9ji6CDX57ldznfgakT0X0wamaRLw8XAhrpguzvoWM+B+
cxInsvWhV4Lm5S5Ee4Yi3Zp/aEUkBklaQjnVs5CvdM0iLGYzCwwV30/c2rjo
K37YgaTRXL+4OfrQrba2wcthMCfFRdAMZqfXRu03jindWZ0Gg7MP+2mkd7Oq
5CnkGITrLmwBJ+gjND54bE30JOVx9z2VS5sQTDvWTY2Ap7uH53Iu5UKZHDG0
eMm1GZesrwUc1SE0qlVadSOPEk8QWDCzSSpMhYp0YRZnUXnCKLyQWyflnPwg
tUDLJmO714L2hFp6pXTf0A9d7rk4rUiAy8qClEswIPrltoN+I347UQyX/x9j
fhgNmZclGo42Ga7IGG9onKEE+dimr0RdnLKAYH496jWr0p/sAq3WuC9U52Sb
IlyfyaTuDCPiuGywvxdrj7aKpwv0Cdgoty4UyMGMoe4bfvUDAnXzwYMAOINv
eNbbxDFqHRcekzalK2Xh9xn6Ju8orf+UnIMJklFgShH6/45c2Is1h8rlarFB
I2WwJq/24EeGpfudr4+r3e7IeHwzMI4mplPUenSIgXfxU3WyoouxKhlzABXj
RSXP2YdH2S8KR5daZSpj8BHNqxuNVNoZSCyY8/BLMpM6aG3ocihu8+VvYQhV
leLpnrEXwXfAFxJvDxo+cVvS1wEe5IRLuO/iI8cik5tjaskVFZkT0tSJKFnN
p/IDJ8v7Vw7MP+kW6q2zI3rzJI4hJ3WW9hkMKai2C4ZXg9oTgmgzVVHaP1kM
B7+Tyr6yPs5qW8mKLoyRelBms2RTp1lHE2PQ9fgNjJt13BkpHh0AWNNC+WF8
j9izyLCm495Ji87g/yFq5VGokqojTQTt20r5F18FIq1bdKw+F1a6ena86k/i
+cJTP0yR5NDuRf8DATB0KVi+O31CsOTmSkpK5XE8Lum4jH7u/SxkpuU2zgxB
6cUUzL5JgceglRaceCaMkmPJHwranTVQMuDWQvbf7Xd1d68N6D1Kxi0gwDsh
iJwuJrS8pEPhwg40W9a3YHgXrhBV4PxRBrMJuHLCNOI4NbuCH+fwW3NjlBiX
vqRA1hppEJWFv/lRK82WIyuD1lT3rj8E6my+EgH9wsTm5U4EiCntVcvhhRYI
Pae1vyJNc+kEQryxbthNT4YFrXgDu8xMqNXY+LmdFo5g4HR0l+g4RYwPbjE9
IGkFWBG++sslWc/bgPJN9sKaOMmCKDyzZHqoDRJBLNArPdqVxWSIqpTF4I+P
c/M5UtzjcssJwV4WMj4eI2jCFv+TUaONjfavpuU95Y5VUyZx9VIQ5MmODKgS
MoO9D4icYDrqPy/DzUgDS2GF9ggHBlaV70FdocE9TtAOAZ4XfkyAO8Rog0Nk
s28yfLN3T411qGfr47ty1Z0Hb2qjolggPtAa17AQzlE1xiCVcDa26o582af4
tySlKeJmfQBnuPgmmcafkunP7m3MJOObk9xbTqlqzdokmaVVM//hxbdRFWmy
sbnFYKk5eTzHqnoyxQXtKNh76+A5vlDvrGphpkx3CO9pl4VQ6m9Qj035vkKX
xh7gNwFzs2cIzxBEiNOB4yDpLYNCle0NTYzP+f/eC45TiX4j8PxguRetO3jz
CK0dH8kpsV5iwnDZBbtpIyB+v6XReKTd6nAN2Ft4ZvLNbQXZulurip/jy0z5
T7+SZV+Ba1QMR9OM/IHpCxaUmPJEwKNDtPxJKNKRTe255Es7m8D3RXFQ0L8C
FKqkBWT80Tv62KtPibkxITSCCfQg8eRF7XkqAoBTkl2uU+pm9eYMbf1wTfzb
k3IKoiuLkecljsEOXgphmvk7DqvhhvlbJwWss6BPyqVq/zGONznYJiwS/IiT
9qJHQoipX/1l2sibqa6wEq4YqXdTPkxYgSeFyRd+z9Y9ccMMaixW9fiRQ+op
3SJiZhPj70DbnZ6locucWbN8bBDFwHB/gZRf7Ug8WYFxYcjADrl8M7iP1H0Q
EOJI5g5VyuAJe7Hg3rQEMOnbgdHHD7nB0OMcW43gHyEan+UD2oC9U6xpcPtn
IAEKgTUC82nLlDwKsk6k8RkRv4eXyxN2j73OlVMKpBZFH9+zV/xj07s/zLeN
VgVEWOu4RLnFAZOFfJW5hAsuyvrcujAv0e9ypwtQsqAfeCnuZYw/r7hC5V9z
yGNPs6gEmWL8KZVoo31ZqKf1JpGDYT3DFZMyGEojBWY5P5jXHfuCPfrdA62X
oMIR3XpK/DW2SQJz6yLrCFQaNRuZO4hVqxY/fhbaxn2NUbmtX7B+Io+Nq43M
rbPGmetVAKLcFMbJPqYyZlEX9z5Ch4mfCACQ3WT9sTQK2ZslOPw9EBfUObhC
dxr1AaTE5WnrQD2TxsDoZjiM1KQyRDhcc/HglWq36KflfPdAX8FmOjJAagQm
lRjAxYfZF3ia+F/APpovGntbkq0hpN8y6Df+9d2XpOk8qyO4+DEK5fW+D8IO
6/4CQiydcraqt3gflywO5IVTO2bzUC96jidDXBYnumRImPWAINqsjrfpeb34
TEEyO1dTj2hZHUQjbznOatOAOis6QgaW8pTLdmq1Nxk8Yey0V3ovpr0VrFx6
uIpCKvs4KQPlYivXkVqxQz77Pn6ilYnqayLnTPz7N/rIKmTESO6iA+noyr3/
PaIh1wXlaQ4dt9qegohgxdDq6Yvor9FNa8jwRxAX8pj/pmpoHBjd+MXw/NX+
Nl3iQ8USKydajHg61Brkd6e3SzhJQ3Gk2ZFziuFj9DKWUAUhWbyDPNoJAThP
jnBeUTUgZCCl/LO41kA/DUd5WNyCYjfn/zJOmM/VAeNXewwCyg/90h619DOO
lGjU0VV9TtpjZNJzXOmbFtCZm//e3WHF5syjah54FXdeNM55x+jreHjm7ivT
7cYqzo5qId8PhbLF2qKSk7HbPpyxcj0VNiBHDxGkdrVo1YBQcw0VWILh09g2
p/EFxsmtIDiu/VPtz2wLpMJea+6jYcHy1xTOKY2V4IMYD0VAy2oIla1zPASK
IaNikgFhMv2z9twTQiFArGdIsTa8vv6QmBBVb19njU3sf1cQGka354hoVGAb
AjUaZf1r3hl22KUZ7lwr+I9Zj97JdKOoGUN6n4/8CxBLT/OtEh23Eq4FdSWi
fiAzrPMgVk+yTSA1iJ58cqTLncBi39PLF+zMvG/MTtZHdTEFKfmaaVj+rIAY
qVxSuIqU2gKONq7vN3TgRWnaHoq8MsoolIZKtP029KHttiOj3z3BplX0bfsu
b9oXLfhYPdNTtGJ41eaYpnMNCsFZ23g2pNMFarQLFsGDV14gCW3jzXqfk9rD
OXgC1naVZxaNEeh6rsGy6qeBRVhztpcEjXIC0K8ssGyUGsFEpKCXRCheYCBi
PPPXRvlYfjy1a+GEXOYt9SM+LemS7m3Ahc28kQewKzqqI4gWgN8VVtW5mfz/
Dgo6QtkdId+c2fkewGDkH+FAv22S7F2SXSW8yUDfwiD6MwODaNYt2E7hlL1C
90TmMvfpE/mc4JIFVG43ok7eSBpN2fSwDvE6AHN70FGeYurFT6SDJt2xUweA
Fhy/1kVZhOsiXe18WEUB7K98l875hgnrUW6O/TSLXqhYH7fug0Ku1Tfc5Ud/
LhTzYA3nhwjUPfySuolGRg9EFBuccJFKOTBm7PNXNlIHZdKact+zNzOO+LRn
M4b19/va3ybf8Ppk21ugOZtg6K/uKc7qG5yFjmgt0UeCinCLXUuAPv5RidMJ
IV5SueALJ+uZkqXZ0x/NwL8wAaaefRJg3/afpGM0qrfBJ/APhjT2F8rWiK41
nPXDjB6qKTFggQMIu5zm88Da4uNnwg94wR9KqVTcao0TBDkNPyOc3Pu3NO6Z
F29JtRZlUOmg46EGCLMLykBUi3ZYpTF+DgCugo+MdXE9L8YaL5PgZALlswVq
FTBvg5R5gGI289I35W/HPph6FoEcKrzvIa9cZ2ClMHE/nuiQfyWaII1Xs+k0
78oLTaz+eL/Rwaxbv2ecim4LhqrCA+e+khHrIfkK210FdMaFtNzmsBxtnp6U
P08+KXoxTZPxXlBLl6USk2Z1mulGxd6YKRz6DoiVJs7v/UOfv12MYufQs+e3
x96XSS8F09HXbylMI2n8ahdMFCMoCfFdMahttLMIufQIM3kRDlWN2wiE3q21
ULknPTjQjUbIQ0Uv7UMXrVzFsSXH5rlWbqQunkYyJkRv1IoNW3qB3dAmbnfG
rxJn2Q6o8hIynr6dWZhygodJWl6oBPUnhS6/ooYnUzO0bhdSkVSG2nbjWYBb
Gjaw0HrR9JqKJ/evA5A7cO/EmX0LHKU4Wj6v3ZSU/s64Xpe4spQCMWNViqqf
M5nXC9cgghvpgLSetrZHGGF5y3zNEwHecapJrQL8V7D5HYovD0xM+nQGbspl
RnO74wsGZlnN609E7r+Ft7B64an9XRdzaBJ+MrWX2+j0g3/7FPYutUgTYGya
kp9hlUUvrPMSqYnd6DTWGU+N/WArGVq6b/wj+ALlpb8BCsHBhramtrR2j4/E
OvS6IP5cp/LOgvvOWwErTMT/k3QTOm/rnCnw9NMDx+brWNtMN3YRkgGMeP0N
aeMRsuDP1lLLMYV7F6wqBYdfZnqJtIVIrPMND1AWDFw9UdRtS8pc3P9aMrF2
2sVSklXX4PYcuyGfJ/LdWw063djnSQoVspG7k3Qyoe+VbZk1ikLGJBb7WN2e
67J5kOzdst5KR0M7UPCpwoaEv8It6ngVAapYtWwmf8t+rY5/P8TYhYTgjAJ6
yvinKNZvRxZq+dHq0a23QeH9iIAeZamK5FxDxTcawqLjj2RYkk5f/6u4gaYh
eKA0qmgA1OM2hZlEUd2Mrf2BfYAPuqN2HbDDsEPsG22so1WP/qz9bfbW8Yao
4lm/PLvLb5UmypjE7llC3BCocLcfemNhwMAdDfM2Cdj7+KDtfCOEz+yejN4N
27D3m117hEjEv5kwbY4Xp0S5unBLw6MLggfuLB8YKlhG4iOrZ+YSC10LQeTS
HmeEkxYDhe6+E5TZzlwVLGaxDPV1DNjSHsajHjWLApaHaeBbuIW7LdzSdQkf
CHMK63Bajg7lsOEvkBLl8diXhJPgh0KBE+K8d+nRQj64XoabM2MrORn1VO3X
Tg2YGAFYlSdGxLqCBjuGAx07o1nOAKiA5ADchNbmHYaG1XGyKkAlAOOB8iRu
rXlUeg5mi38aaBWJJbcOYbK8vadV5fs439YbIVxxUZx15w/DeQeR9qjsREuS
pxh3pJ+ckkP1nzaG56n2v7zjzDZ84VK9lusnWj2rpP7gDgNHmzaixdLREUaW
2Hzf0YWDV3Eh8kZ2UR/Sw/o6nX+if63dVAR4Hczdste3bELMX3KSznvHmQe6
k8kDMgTd7o+AjVR7ViN9N1hwcjHX51ejaQ5t+mIaEvpUTyPbmPFBVkjqQ6r0
iA62uzndD0ViLQhcYVXMdCTsEUk/Y0Q5SlfRl6ndq4dzN8KfsISGapozda3X
o6PN60wPsmRe1Lc2pZpnQfxw+l1AZX3oN7eM/ZyxIW6rUWUIcdTfOqs7VsPf
CxfzqdtiQESHol3eAl/bbS72pWYnr+x8hQoWO3Ntd/FXmNGRBGNF8pKD4E53
GsrndYLqt8oJoNutaP5RzmvBFeTpaQh5PT0tebBoRk1Ir+E3+RpxyYFcTQVh
0auk+unVpi3HvBqu3hA7D2pEMi75HgI6Rklz5pcXKSIPNM9CuaISzzR1Jhip
J1a4dpELNgWlezWbpS2eZM3BDmykFfyrTx9FVfoW0aTRrpMTESKVEmx6J47r
cOiE6BN3lQ/O3kokW43VJ8/UkNwaEml5k94xWwVVZw45Vrj0yLiVBihKGLv9
RlKT5oUuwmItLsO5hCcx29SrmQ3OCTKCN1As/5skgynCSGb0s8scTDFk3L+s
HgRWkDlEjv58huOFImCzuO3h/pAnsPJtokQceKTALuaYHFClHIC/1mwt01bG
OaFDXIPHQEhnD23AgZGaSOa4R/2iEBXnDONjZaOtg5pNvqocvHYHRZAdBvA+
qfhZlK8rnkdJbls4JPIjRViFPaYVyI1j7rtccjlMWrRLKciCbPC65IWDA/yL
Bf+O6B86y8HwJmb9kagA3xF46Atcy/C8MIbp+ae6HdKFA99TWB0teEMjLP4O
6QhdHplSrHKlokpBJ+SXvpUcv0si2laOPnw8IweOuHDidOGklnk3UhfKaJIb
qAi8es1cN5pZrTGQ4ufpqX40dcV6PO5AOTF3QH9WFUvB115IGte8KvXOxkXZ
Ar1RGKh34ItRnHUHZ+ALcWSv0yAO13wZodThszKXvuJn243hDMVe2O+v/8wM
WhRVmndUKg88tgrGC2d3xphG6wg2RZR7japjuhw7U9dXj7gDKsDe8//Iq7qy
Z6lhf998edBrAM4NPdN0Yateo8Fqszy4ZVb4CypHt9Ac8R3NnY34HZhnOwqR
WS0YmmiGux+bCQpzUWFh7osC6xpGpS/tTKUE5H/uhCQxT+8musinWgVDVwzm
JV4DMAu76cTK4TZsKD9Jm5m+q8soFVJOe7VXptt9FDn2x6l6VhuhmALxc1c0
VWhJOEom3r62nUVECORlEkbQibwygtRRPHVVS+OaEEcr/NY5HUl2ALJqzgsr
h0R3C3uEZPeYh9ZYbNB4XsJfbRwsBRt3zPKTxq8qWjRffFvuKtZNV9kpkQoO
KaLi5rCnV0cMghrrkZ/hUDxPXZj8aMNH6WTYNrDCFI+HJY1/vMtzo4B6jNUj
uENJoBz8EJS2TRxSlgiRx7ZKyrhwFkGe9w1mchjBP5aS3JIcxmFp5oT0OetW
qpXrzV/xz4OafXwOq+nyzZTjTe+H6wYE5Cpzs+NO3KNBgj43CF1rh2l887MR
4GiVwVgkFQkWCt6ExF2k7TtnTtFvSxgritEi/eJfoRdbSs07Y5QAOyY6MYB/
e182qJrHrwHjLjGNQ7XhWOsdm2/d9OnQdUL33ajtJzTPhbxpO0slsHxpIzMJ
HDmulNuzn2sYhVe5y4RK7b+YAbxpNFx1m+ytV/rZb6mj0hyo7A+sn6GQVVIp
kQH+ijwT+Z7FU0zQqwEQbZ4ZOEGrZXWsWPKaOTNpMfdgrM5QY/xh9P0LU1Bp
JyOEup+UgfO39aXjdD6I5eQ+S7DVFquAh5txBzzQHABvzbRPE8EAlOPm3hZn
kCNjudU3bq1fS1tz4DNlViBZ5qGQCbLv64c0n56SJAnJ4TSYBOGH/2IBrxn4
mCyd2wfNOtGm+2z9BM3qBNLz480n6nb3iEjBFnI1BdySFlKLgN2lwYGYLmYW
CUziT2IC1Cb9Am8nM18HcCSXeNaesvaLylG3ga6pVXmdM2sQRgArsXLudNfa
AVy9w3GMnzci6rDvOrAS7tIFPxzt3xVj6Wl3C5WMomMOM9sz0izrudt0ze20
GP08EU0qNWEge3spE8QUFW+ZZTbNGNDKNJJ6Qg7pGBP/PsuT4ZqFFBeHNut9
AjIGSyeqny/oPIK4edny1qXChu76oaxNd/HQihuDHzOT/WeSauGTS7Eu0qlP
KsSLNBxdeYrS3mHl4vCafLZBT5mxCh3qMCjc9tOn7jhAHWdekUKcTmeAR7SS
p9A5J4i7GMbaCW9KrDiVG38pJo9LuDssd5j4efs4P1mZxu/EPT7qp4/W8+vi
wvbDMXJsydGkKXYNvPTyFlsaPP6iF6VINuhf56qh37XQab0nvEizpHO91KQr
0T4ScAhMnSXyUJjzmYbZ945EOCg7ho9oAfRRV23c5dhb4EjJojowvrozQVHL
wecwdHbeZ0RUK53wHNUbEZyv5mmaXjGLLU5mzc7A6d9EjimToNoeTRrahI3v
tZ2Hp1mhpoRPWZP6xF+i8hAN+f1r8Fo9f8eIU3WC5VUkxQn4m4rRMOwwQvfr
YbsiZvOgdI7JGcD0QhpA2hG+xrsgbh2AZUk6sfemu3Gp0AMtXAmbVOEg0cg3
yjqCWcLR1clQOxwt7MpvNd5tLse2CW6umMc/5F/PaYsEAXSUFkhvRTx399Nj
IaRw+tFgQYOps6dLe1aGLH2KTTIMLVZX5YdvVMiBhe4yFBPOuDKG4UOIMZFI
s+0Bpw68wQQKrUOxp6KO1lsx+9e4bqnvnprlOXZBIGMGEqWW1HAg9m0GyaR0
uHoLYQ+sVWtQeXYTMrfKW668T3Pu3kTgRM9n3KTLYcT8jeNmmkMsSghh85Ea
ats1GfPSodvIzflIcUBMAwu8edtkBXI3vYipgpqJPjus/KmFSfEO/TPIJwR7
TLPtS+q+n0UUfGvgV/TAFeMBfUD+XU4yNK9S4qezuJ7xmJ6vCLGZaIVKfMoy
hIAySBxNWUduWEVcl84vyJ2BfPYQ+AOqI2la5bh5HlIOE9HBBifBLsm0IZY5
Me7LUkQ49rT5D1SNvr0CqahxbE1tBxam66wu99HdN/4/oryiPPUR03ldNyOp
Sc+Wa3ey/2Y+/pyWmxRWFWr9q6IP/5XpgTPgoK2dAsV513i271Co1O7FqCi6
QULQyIP04QMgX10L9I2rphBN1NjFs2pb0tnOzDgRCD23HTl3c82/9FNFD4oF
qGAMQhX2zfvsLZSWHANNyjwRcUIhhV4eaeuHaHOkV2ECagvPkj0CI/6Yuj2G
zvAiCNSfMhDW+RuFydmWbWWpfchffUU+Q2fB8ZU1ucwYSuRU16Jzm2+uZJJV
R3GivK/EsS7sAzPlHnEtqwfBboN1K3KA9FfgeSKzqUEkXQd/21XxwvLboh8J
HPKw1uqLjw8wzwLtP5ftHzWQI7cM7YVMyNZYf3Qw9/QPgXJjniguwqR0qPYb
l7vseRTiu1woBwvv3rwDRVSPfdNHr1Jj8TLpQ//fAmKgOOHozKrKiNafTk4M
4QdirazfqrCEhu5cSaQ4CXFFxGO3b5M4ThPaf0H1cT7ozEt879/bekhxOGH6
uN8re7u9Kpr+6p/tcL8QOvU3DIiRf8e4/Q3T0AEatMVpwNzDtRTMuRnWGPkp
FcVRb17HsR6RI5G4/8lHtz2Vm4Hnx4MrPZ2zDYUZ8C4W7mWOAHyXEiqkn547
N6t2L/6s8+IodZNSIALg5xNksGYCP3FL2tFgaMsVzPMalC6gmUidm7ZUE561
f24ttXfochsADNIHxWyWnf7D2mvz+pRfSfYeqT4jRZKBmveNcGAmjbME7GjY
TRwccYK6BRkQbywhxHv26QMTjq1EmbFNqNQeZ2gm6LrQH0G5+C7ZjeVw6rgt
9V63gbfv+IbnV3DhcvIINB4pOEx1/l1aLCRTrLWLiMTnBjwaSF+/E5qvYUJu
NYZ5tf2QCCS4pMRAcMMAQl/a2OUZ3gxTZpvpaP1ItKbRJ0A1iD+KxfrQdTWM
ewepbJ8SRvUYOOdm56b10ItV9q/Psgzj5MMtF0oVFHsL9l3tUSIz7KO+2Wdy
vrpbBA/m0Ie3iJA5ejSxHqi+qvJLpjLfsWSMep6U91eBAC1rGDunQwglXFCu
o9/3Ajx0s5P+Nep+7HuiRFUso/21XfQ76SJlZsSDeiyvl/fVe+GO00BU+PEp
GQ1aTA9H8+que8cdbsKJ9DIOsb6G4ZtuInmrWy3hEgowC0rKGFXuiEtNKd1+
Kjm/ILH87wvG8owgdW1p8HVhrDE/0prWsVI4H1I2d7FLUYFWQAezzrtvHgqe
fv36ATz7PuLTMFdQ+vwFUGTmtRlCfdqNjxqc78zXYlWRpkLnWVXx1ftfY3+d
psE8ByRtpXP+6lv4xL5DuMIrzC0z8Z0O5Sf/W7whiIYLEHxw9P7uWn5JAe0p
WxBvnh8lHHlzqGOWPuLtCtJk+mfwVxjJ3+8kuNL/j/V85o6ntvd5GA3mz5Vb
P9LS7W1sl3a/JA1azeHxJVXFnnMfAjdWchv2zrX5T5rCfUXhY57Ey7SWnLpT
IOfGb7/o6FjkqlTvtemwCthtS19TaMiMX+wNXH5/khjw+uG7vFMpZ6SjlUqX
5pkJTAHFMH8tELo0naqtwSvMI793vXcWMtX15mVh8mgo0PRHGPGJXmAA2WU6
g6fDBqJY608ZmktfsMVyXIiUm6DqWIFhdrdnLbcvzfl544Xup50PZso00TQ6
Tmwycyx5mYDooApGqoiNq2Ldpt9BWswJd4VFKhIs0yI0gkIZPK8ucZRWue8b
HF6tX0aCO/gMuAhB9YRnquaGbEzeg+0Sox2xmHLH6bp+XGUuA7Gs1mmGX5h0
0P3xWqvPWhkZ1Aj0MaemEf48GRigpDczpdHi2hQq4Kk+tVeYmrhtPCxuoobU
O6Jw0XCSO23zLEcjjEHjlQ3AMWCDRGOZYWfHbpj5D3UHUYpwQrGlMiLZ+1Pj
eN4gZGwaaRkGIp5ZdcoRS6fQU/QLwDnfzt8wbrMQuHabZF59agE6DKd4ZW+p
Prf5VlnVX9qESM5tkp4u7pI8fjLhlWPdCBP7WO1rE5JRA4mphdNndzI+hhhg
ttw05Z09GXfZds/RnI0N6fhP1oYRyejQKFyXkg8pFPw4N+lNQHg9A1Pkv7xp
3di2nTsf2aqzNwtP1miQLBllSSPxtyB1LExu3MBvFOUCoYr/eXBRUIZiTDwn
OvlDPScqvX1v3aZRl1bkODw2gwl4k570W+Qhvea6ZJcbleDQuWM1W3JCVKC4
RbgadevY+YokBXIz17LYkLfqiYPxG4TYxiLmgNuFlFeudirqSNYBf0P+kTNx
DFlji+S7U0dP1qYBr52QK4NfDYujTltKSeD+xHi7NyQmdGlPW117mSSFEKrZ
usU2rCAmFf+v2XgZ46p/UlVb7gHwm1ucgLnD1HZL0dBTS7vT9v5/oerjCLsn
nPkzs2GSvgwrkeyTmab2ruF+LnKKHG5d0jLXM2XZnmKJNXaZzovUSA/aH/SA
tBTxcANNKZP0OghYExFj8fMbZPWhxkFqeJTxWFrnNi++rbGXEI4M2RquimiL
NaARaxqmVq6vsPM9ECSeT7k54hQAF+phiIO+Ssw8RkLpUSm/jokhyztLAhuG
Xdfpq9n9NiCn+5TPKNmJ64JCgyfqgiTYuz0Pug0PDvNYhfB++XsFq2LSjnaO
yRD+fnOb/ZFw/NBr7mFVhu/9v5Rj5fnpqZ+wdq8MnvEue5gK8fAbQGX/3/Pj
LHnc3v15q4G99RvQI5X1H7QBbS7Hz1Jr/oFS/cFM2nmydG62r8BIdlcfa8UD
q9bcgnueuzTosNTBvsBzJIWR6VUYCN3TgvDIBq7PV6h01TZ4jYhXxN2XXcbD
Ohef3hWqC4iiudsCq5k5ngNbAZzLodwWYA55qAzoXDpxyQZKFhFx4vmXUUA8
/ZkFD8K/4jA+W4HDipDryLzld1L3M152OGSIBzX63H79hIKpN3AFWePhQRmn
14DIFMijqMoKNIcj4s6erysbA4nfo7gvdJB9c9pMSjA4HidKx2rngeKQxYj6
yWiH+stFXQ6peztbjgkC5Pok81oBTZdKwDOxsbqkHrab387gfHujZW24XRC8
P1c+X+Ezf5gl3wdm/vsS/VBFDi03tAweg3E7+BevaQIWeCtVQ8PiEmzJ0utH
7V/cfuSfcO1wT1aZYg9kxew8/253Wcw9d3A4AgNB9wnhBhGr5CJdlLb+bKRw
5Xf2oOaVDrjSlWjkrnCaZCB+s7oCVw0VUGdPoKubnGTqxOQNE3VycDhcUgl2
sFqPbUM9+9XvdhJxD4gc3Vmvc0OM2Q/OQiJfnQYo+SOkqBJpHsvupFNi9xul
QfY1E9czEQWcdEx6S5TH7TCYGbuURipbC4VgqUw6l2Kwn6bfodKjxLzYEyHJ
TiJ0pbO/lR4tWYcWVm09xor31kHA4c602acbbn2sk94lJmPdzX+NmjpcrfX7
fLYNcYfhcHc71BS26cSPSl2NrIrtXs78x4027OEJlcpzGnPiFRcWai7IVKkh
uVmRpPqRtfBg1SU36tgoW0EX1LbE4Nsg1cwqBA+dknPeVEcnn/TYoPWr2rj+
n5TXB+0br2/4miPykFmG6zzMjrc2BijLsnkpOQH4uP0g7VJ0gpZgncIfAD5+
lHdWhD6J7xDeE+xzpQ6oWel0Pr2oTk82Ck20soaUolikkYrn7csoY8cOyQrZ
MTAbluLRyny1RKERe//dg0tGnxmEybPJasoueZXqyziI7nnldY0D+LDEzdJb
0c+I+75yzwikbUis3OzZIa3+k6Xv/BWF1ye2f3KYvkeJfDSWEnozxL3icU98
DKKb9WBsu7BhCQ00wXcYiUDjG26qiEZTKqj+6X9ZA+2YnS4vce3Kf0Jt2XfB
Rz/kjy58Y/zHxjx42hhfVYFAKGSC/qYpxD3sps3vN9LmB7szQQlb48eGUzYz
hKheyiG2idmpDzSSIsN7JcutVnv9eUPP5UeRPbyJ7WVXUDoaVTLdsWoU7Mlb
+r97uvSRpp1LO4gaLqX4bX3qySANTJLcEPHiDSXTazi2OrMKeysSwBBZquEK
2iTA+bOVMra48Uvrmwapi6vzXTzOcBD1QSReiTVjThhC+NY+qbFhUHJt2PZd
kq0lCSmIhEyQUhDZqSxZ3RZKtL3t0yE6v0Xt+Q1E5gHqwDehXGK/dPU6QtFN
9odJ1EPcVNPZAN0vsI5VJjLoIMWydoaF6DTPaFFDBeAGma5PazKnEfTGeYGE
izGjgbFZFIdEWo0mERlXEExn7IlRbeSH+mA17Yu0jv57AA76IMxIAQJFDoTq
LHeBpEE9af7jsCnxgq6pGuMOfp1FTCY3PaAHmaqOHLcSGGZShKL7Su5Pdcko
yKKtg1A0T8UWqV9BG8nV49QeBD5R0Jl9zPsiJ6KifnLD9q3l5G2fErQ/Z/We
P59LjwMmpgYHdf1LPQLPi9+EcVMkD5RgPWG8dYikfJUYykjSrwQtFC3WyCq/
NMm/38/aOJx14BZRUFYWkKaShsvTf32AVVYc12h7vP+9ejKjwq9Vok0y1ktW
CqH3sCHNihIyJQG4JJXGM13L6XMzkkqR68P+iANNaSM3OPiY9qLFGrKg0LZg
DzkL3d4Bhjor9puMkgfqOaEC3/lfO1Im0RoIkeR/erWcGubQw2Mo5BHXlSt1
4jG46WaPAETnC6D5GG43vThC5xD7ByZZ/1aO+RpGvRnPopeOljfUTMoqVAZt
vDPWT0YiY1zuBUyP6OfzDJRrAiZ1ARpQxDSrf/0ebAr2mnqdCqZzy2tqNNlw
Y3pxUMQME6wXAqZMaJyujzhYv+DtPZn3SiM51K0hXstnPAn7DHcwK/CT/rCx
v1st+MjCQ35P5DgZVw3uO8VxMJCf8i52J3om8OOS7a4wVW7yWmrjAdP/+8bZ
aWbGwLkSBwUv7CT5K8omMd8egPm2gxYyvkR18gs2S8rxU5lCqk2rXR0tIZVp
v77Ljvor8nKgSCcbgWqVAaaQi9W9vTT4F2hshl757yMnZsk9QT1yCPH7F0gX
lNjN7fmAmz833z46sVEoAFRzGQv7wrurQ5rNwPhBwedhFTlpeid4RKxLbIPY
1tIhwWePDlNryIRefzR+EgxrFp7zjyD+7Ft4gtkcFIXzhwJ2v5sxI1riOqNr
4wu3n7b1heRhLhSWgn1VA1+h6hlOo+APxOQmEyrBKq7OqAf1Y+Iobsd/tI6C
b9WFhJ38Y6UnVS2gNXPPkt0ZaFoid3hZOpYWIefKMMGvIfRkB8alu86Umv7+
4NeyINaJIRWB33G7GkARKn6OFIENnke2EOARKJZPa4g+MgowJazB19//vq3u
zS3t3Sc4t1tt6KFTFu9m0ksNnaRNLIZ+QPK/jbSDCvlmg8HABRNuEmqZeyuM
Vj6rvMM2MOAzsfoIFlivc3LLtTJ6ClHPZAEXUnlTFW+ky8a/ux++PM5ga9Mk
OlNr5stmAM+xNXaV7BQFiJJbs62uDwya9fC1yNqQnL4ybwx/L2sToLbgxh9V
M5/ttHLMW0dH/wg4sFit/CqOgtZDQPc9UZD9sGsMXy7HxGdHNfvi+HTVmohj
OFt/AaXJZ/MB0cCp6QcydUmpPJ7wqb/Uuxdm5X6O5Utvfu74sz/7wkTmiA7n
ya66VMwecs+1SHiGIZZ1vPAHTAnjZ6xLlrMT9pOaHxlisAj7M5cc7rmM0hfv
9FneOa0OPdetQBzLLUm0e5+FZe5Fb/VI4xH9GZoJHMgiObkIJlN48EkJnYhT
65OkRXinE6EQA/bg/KSw9wCBS6MO69Y219Xb0/mYNQUXFEthL3DRGfQUGrla
y+89BYGOJjDJ+pIbisiZF5nC1PYaWlNl16Gmi8hmfz4MvJyt6KjyZ3upj6B1
1wghya+QW6M2PQLeGB/banYtnd6FpzUNUlZeUF1nieyGuHOJDkQJ7PfZ2KNa
HuFCyFQ1fKKRbu7T4liA7VnhbPE+jN8KmZV3C2n9sbvQQLhzStzBPZ5d1rDp
qMgThJY6N1gucezBdOq3fxWEmMgT2tzaUhAwnH3aEgwC8BzUGrPfVu7hF+TS
tuMsKdGm8OMoNbPD7lTGmUcCu5YMReGbrz/iZEZzHsgmVOAcc8O2nY588rfo
FpTWHINNaohVf+NSknyKXg5BRPGfISLVoMnfst7g5Fu+lQxADPU0DEVL6jX3
7CGIB+jBaI8vw9UEPLfWebmiq4RJNi1pNbApHeBC1UoT0CRTuk2dRzsSqcE6
883TFNdeZLLAsMmiEvUmAeHVe8jERkw6gjm6w276g/TAzFr+IXq2nV/cEzJg
0mOTd5hJxdYovxz4+a49UsyS5D4wtdb/LYPhEVYaTkGSUVIOVvNgimYl4mKb
ACdj3NVrRnjbdxp+PZgrDiFkzK5dAdBvqcHZyDEIKcODD0krDwVmQz/m6xM5
jt60NJegea0rX2lMnqjkhlBVHMe2HfjG3ziBCk35sxP29a14uNFrHB6SHL/G
R2L98wpWsS/fBtox6sU2GUBIvX+8Dy4qit0nx5T8uVyIiuKwWLSvBbfrNuoG
19aWCdiLZFdGI+IxukGBxxIV2dpz0c+WLJ/W+rJQKCiUa+8HIh3Wrm/yMeQ5
1T/x607HAY59UtduiE+mqiw/K/L+FCKFOO+0E/sGEanlDRGXcB4aLT6+pSjV
AXqWVzGfrjVhx6dm1+HS/47WsgOMbeSqXNh0fh0fIYGUl+UEblFXdy6OjtH9
PJ4Pp/tbbdq6YO2MNCSLjp5GgR9xahgtFmZIryXgwNCmGBYsPHwD01qHxx9l
3y0Xmi2q5id3ngXiJ4MEco7uRaWL/K8WYEobyCUwM/Rk8cez5mXYjc1Ny3Ma
AP7S4CRkQSp7QJw4gHCZ9DdOxPBcc/6w2AsH+3fcCqTEVrzedsakbqDd03Xr
jE8g6w2Hupz2Tj5J5epvL7cvlcMe4ZQ/dFnCiTTUwCFpuFq6lFFZfEjaTsXP
DyVtS2xc5HSvs0RE7EKjAIOJZQIydsHLtMPvmyO7hA18prPdLTkynBmBGQMV
mp5A/dqsfBh54V9AFLOq/PsfaM88oOjUMBnQYZ4S/QMVYTmNG1EmxXPjild1
ML2uVT8PlQlX5QklSs219M4D/NNRGqTYhXksTy6lGKOnM1og5fRF9T7/j1eK
CW/AKHPPCbgNun9mHWWCREaF+IGe+lFsVD+yZZaEOhBWq/ioS3pHVmxKGF99
gDaRUTzBtVdCFm3m3Ew/aTBFx4E6T1kzWOEt9ZQVJc6qwyYpgE5fn16Ax+vT
VMUn0a1kIKOE/Yl2f55mWCBrvMfOMT73i/EBO6zwtMwqGKDTxlbMEzBW2FBn
Q6ZbgpaZfTUeTe8K9foYm/mrxTaCJWVns5xPOJdlLhW4oa5XMBHUUQVxvsEv
u9tC3vo7QSglvFTWTUkAjDQxFExT50rYpVWXSmINOdOLWGNstUlWNfPQxLok
ycedQFEa5ddKLdl9gp3p8w2UC/yjRYELwRU8KvqwUMX4tI0XwMJ7DTJ4wDgF
QNTsYZnQJvI3EpcM9qYHpRACb5EOfMg2tVKlWLygBQUOYvkmqi9aWPzpJ9Hs
euSnsQcpXhO67/5kuSL2taEJqEdxlASAINP+j8bJPM9ftT34NaVEKQayFMP7
EgSD1VwuBqopQB77Gwme+aZk7CASlWUHbeT2fPlLkSiz5a+Zcqs8DqurOVeo
i5CfmNrjCRwyKND9ZJacBX/0OflqGtkEJ+IuhOkEWSmsKG4wZ6YLKN4Jab4N
GNYH1pO6lxuoQ/YmT7RBM2c0EoiJeOB2fBh2fR1BCauwFuJ0i6Utdg0trX97
VAkhNEdZxGgIvTjwCd+BXV2mJm16wrKr13r7MgBG257+A8Nb3wUrFICAUNRC
SfUL/G11pthDfBdwEiH0b5su6oao8Jn+OBNQvkFi6xaTBQ1vKevO+n08DA/n
klBO0v/PQNtOZ/ZCKp5PlkCQM9VU8F6kuYszqgffNUNnbQ2b83OqX33xyx/y
zYlrXkSTwf9Qyy1TRkYugx/9wRSBIFBmXSM9t8n09+x7hhBcMkZoCKXDidt8
LsiD+BucsfjMLx5kSIrLxhDJNPciZLwOR0VLuaDSuPErKytmvkKKEdun4N6A
yOoNOr7PZ4KkSyEw36MqY83lnFSef4nMKWvTFMZ0gSIfzU6uUS17p3+IYuUp
xEQFjA7PUXipS0gm8pWSAbHo9UmM1j3FDQUwbjC5UH5aMaI8vI5ZCrSOSBK6
UP8c0eKQoIsoIqs2MO8n666l4x8q8KjdZEp1iPb5qkN8H+l2HVQnEjEdkNh6
sSRUBgJo72w2TZtannvarctb6HVzAgHfGqMB4Qn+Lqnho9ktqI3zSIAiLXs2
lKHkCnFEQU9faSKtgsLOzAD9KtrxFnYQC0ijcARK5tlLgxVbaWoNFcVfkChj
n5IHZeDChhjkHTtVxjMQGyXjLXaeHs3JvSCZDZSZx84OBrw7H7ZMJWgbhdJd
UHOBF5wMXdzQhLfsokkBaLemqlu1XXEiTXPwyD8GFEkjJJYTnqEoYMybX2xr
296kjTpOqV5TwEub0TGtmXpGzKpBf5Ue47cSb5A93gbBbyMZHvVhNlgSrmYB
IvhqpOdmxAPV/r4iuPGtNkomdPAy/11Ccjazi3gLn1FWnGp4qO7hY2rCPMWM
oqd0NSR8EK9uwTa+lx82U9B90FBG/yqRx8hr/iX6/4qG/Ty2Dye2rwTOuQ5D
B2kQ3BcNV7EeQAnFtv8DtJ5A94oX798Nm0LJqzFbn3ehuocLc7B7Lq83ds9I
4+SIbyIxxoZQ6hkrspev8mjpHV/d2OxTUCI4L/VZQi1dSE6HkfCiku+2Do/+
rdBgT5mBygud0aDjbtHomqk1ur9ReM1xTjN6Cl02E/EmeDnvrD+kz6FSelUk
+nJjgecT4ijLhTxlCj94Sh5gFFMDHu6xnpnpDe0Pnc2RyAPArwyEm7eZnf5p
9lr3mCK/fSR99LnZU7Nz4JraZ5CjIs5SzSaXz53xnE2fU9P2QGcgQS88mQER
Gr3QUvo6+ax6mf2G8u3CZXQRZ8pr+mb8ab7agRr7akgWYPDpZJl1jU1uuxuv
1uDhxAU0bPUWKErYYIVzAC7tIV/HiC0OzSh6sPJ+WJpid0pC/uw+us8M0AXi
iBFnyknhZyqGY2Cp2grF160KXwJJ10qY7LUxHy150fUD6vGCPcYgEQlkbBfA
vDuz0Kw/lfomcTQRsiEuykpIEUZqE2tqx/rTuf0i4EwcyT8MPIOjpvHzKhAa
ZFmo+N8nUCTkmlrbHMrNviCgENAqIVdpCcxVLxGcaStd/WjA+WRRJGtowAnq
k0io8daqgh/8NI2ojxBFKtF9oRY8EULUtym0ghh4wWnvhNf7ETmVh0/kQRmB
8jJ4Hy3P2wgF1cXdtyK1hwhPxAXMWIJGYIi6tArJz/IH8AOam4B1PaUF67E8
FrxMByqJheZ/DzBcmONjXJibfcT2y0dMXQ5dur0bx7Yxv5GRJtT2YLJFwpHD
ZHhz1BVyhQTr6crj/G/KYdluvSKcjsJyVpvO8Vaw3QtXyY3HB4gADX5yJhBg
tMN1iLHuf4aql+2eigd25r2qCLO0WwHpgzFHoEOPKUuQhHPQsXdkzq0LIFEM
iH8A/mjuNQ4euH+xqwOevlIQ19UDcnX9gh/SLE4qDVKXAc2rX/r4NUJfdMeO
VslWNFLL2WppmI5Jz2bi6tnkkQBntYK1dgCwKhblx1BvvPYuYP+QrnjifF/M
wsXZGVAP6YEWdaXR9D+WCXFtP99mERW/WDQCMFTXykTshvbxp6bgXQagk0is
eiWCDX2zAOHtvjNOSzeMZ6ufL/vXcM2WnHf6kwXhKCcwiONT7Duu34bAh1J4
FlZ27iHqxr2Y6oSYf/quyCuhr3qiqdlN23CYRBN6+mAyL0zXfypMOJddTmSg
IsHmIiUzWJGtGRkgB6CvcqzMEJtrCAYBTYThM+lADmUlERi8697IpfJDcveI
CYSmNhI8CInVSdvSCcqTCZg9biNiYNumqsPjdVV+Mg12R/jVGRSsM7NNJ5k4
f5VAZXHnZosBT8z0x6yu5xbNIBy/yHniCoXTH5VZiA5l/oECd0BTdj3ARG8g
D4E66DapKHD1JPuFutY5oH3mKWdQooJHCFL0QkWLrbirWm4k2cZ5MNkuoFgm
aa3+R0EyhWnBqfaaf7lxG33SYBC0aCE08+JunYuAgQo2g93AtzFVQ371LkVo
ng4vnQQsF3Dj20vV8qHhQ7iAzJPVt68lzo6DfzHBB7IRkst+shTiNyaK0xrk
ZQ+G51EmEJpWdVIG38BITLiRnjAbS5WBg70TEzzBkk5qkYpPYBDVrvejGKoH
zd6fJrYRwMGtUpAN3e/45F/l1U/DcreXdWETkrNI5681Ni4Ksy3srusQ6ySD
6TTzOXKtf+pMtXsVxcK8roBq7sZ5JgVWGOqPU8Sr6X8wB7bxQQ5CxXlrg+Jb
+/jVThC7Z46TgrSRF6QaCTn/hOhjr9CdMLorqBqYweasKfLAVkE9Pio2hMty
wqYVTNcHd9iP0VG1+JL6ifFLNHUBDf0hHZAFbG10dGSN/Qt2y7dozvKX11F6
PgfxGfKmVULO2sI8mW7ufaYNlv1w/5hZ6Ms6Nxh/1t/WLEH9tbGHejEvJbQh
lErXGsOFXoE2fsdALU/i0F/1yosSJ1cfBhx9Y1r/YMPRrGwZogoXlvK0ppsA
PtomhI9z+VRKGfwQK7yDLQGO93OZuMaQbCz7R/Q+xSKIf2HBuTbSJ/8olsYk
Kl4XnuoTfBNEUY25SlmOiywaN1ek92GR0NxHjaosj5Bprpom0dz3vt2iTVEG
zpOp8I8g+vM6NA2xBt/h++u7scSbQAUFtikf4Kv9zF2fD2mSlytoDIm+W6NP
yR037jy83Jt+4Sup1WCN0km7XETeyZTWW5JwYESA/zt0ZPX/PQHGvWlTplBT
NYmMVMWgzHr+RGJauruFyGPTWRkeveHt6SxKTczkaaqP2KO91Xmt/04JycrY
Mxzd6VlXeVeUrQWaapZw6DOT8O1l7rFGDVJUg1WZ/+cJ3gdKtdJ3MgRoBJ8g
fBjxPjhqa+g1ZiC9jB4BT1byh4mO8FPs5rIJR41FGOEYqpSv75N0rrX2eEZ3
vllP68ROHFBjD9twMR8hXN3Cc6SLQ2zdUz/t9W2f88ChhjoboX4vSWM9BUmW
//FeTXPIsoy7OEaWpyR7D39iUhZ/lfpHmvsdAYqseiseqgqtdnIaYz3LYygz
S90c+f8R/8Xw60U2Ip7mqG2HFCdz0iFX9xJ4JbnCT2re+wDw3a19MrR+diZV
85sk7gE1q3+bV4Hdl27NShCUwC0g063MQJ23Yx57weVArbiMrcYSGUCaSSFM
VJhWqLsNSjS/AbpSnEz5VacatYKdG+kbhIYn+0bbjukSwjEgA44iGhGZvzME
YfLwJjEXwJ7xrip9j1cCi3JFvN4xWCbgSVmf0Jpl76K8wc5KiUt4d9r9dh92
u5e4uXzmYcKtAmlpFyLgvZeC/llvWf8vaJ6clyWSbJGF5RY7/NxqW8u0Ksaq
koa2DkTChYbtuMLB4/5NKrQMvffMZ+DBZ8xHHXOAkwcRgRbTdShOpGHXzNNs
aSf42YpzWQUN4hoiuNF/YxAvbvudIvLvUDoV7NaAkk6zUIUzgeaVlexW1BOg
qVfTW99clyBlvJfOYg0kaTd3b9JqIs0kiRvd2bU+83v2/g4xK/wGvZAfmrgj
bMVLuK7wUjgiV4MKD5qoue0BtgLxEnSfOMHW99xKkth8Av516AhtBtcO93lc
Zc/dP1mrHFAEtZShe+jNIsKRzYtlZ9yKqnOgzpfDgszGVVZhzVFMuKKdCE/Q
c/tsnCTFDEjp9ryG95d96HQCgIBnJQL5CkecXJ1SUAWRN0ZhoLFdBDSc+qRE
PJKLJutJNt40hVT5VQD1KmY96FdN9vt7yyAbq2PdWUPPF0jhwmAd0pVdbyBu
SnuiHVNZCS5BXywcYlonB2rKjn19LXKdKbwWUkZjhRjDeIqtsELLld+ZwTdC
/zwB916Q5XFohsQUwQODqDOppSv7mcNxOIAmEM78orz4xXpg82jzOaZO8ndr
+IftVGx1bgdtEH2Z9M3WlL8Y/24emPMwjiM/Xbfl3v5T0ARBKnk9qN9v26eX
rnFMaVDormNcKIcp7IIPueR1DPI/6gaYNi8gY6MXyTJ/FfIzzWTazKdTtvya
fRRAyu9YLFuOuHFw+BXhOMk5Yp5PDx2voYwfofO2vZdTgkEsx4LWWaNNhFUo
MS47zzPVIbXI4hNXg760PfUj0kUl4JQq6Z66s42UKsQ6MKQ3ycu8jMiUiuj4
SAIylQ4bJQMyDZafHKdEc1qUwd4RYk2ns2nFzarSNlreFisVO2UwiPALvB0R
oHlL60o/ya6eByDHxhaf0oC9t1u5QtntOgjbNNsYFEegE2rxKHhkZOJ78fvR
dASgFZ6ykTUJM2ubJfV7uSycnT/b7LaxDRY+Ys3Ak3y4CrB61OLCtp/Uh8qb
73c34L0ANkcZDUvvHu3pBPoc6pCaus9eW8D2O7GOQqPaxERApW/GMslW7zaw
mfj8P3MOKNB+dW91qFBpZ40kOU0sOWucpdMssO78Wf2zhB6xq2y5qloImXXW
rbwirAMb7kN+eGTrp+5otrkekF3iaHSJ8lF8QmUOAhAGQjdqp8uBUWUkjUqq
SIXc533G4igc2Nuqq6LeLoA52mFRrH35E6gOk5LW0Y06XnsHc8jSwX0cO/DC
qf5YjE8oLeWBnXqrjNdJDekQxrPVTpOGE6cJ3JMMdrEBsgCNup9KQua5Am37
4S3EAhj5g9Z9E4IPRIqwHp6YlpYg+jLrYdE39yfh7aEFU9jlQ9QtDNlRpz+t
+1pLC9sCsw+g7t6AW0fm6oQr5xj4ntcIEF4ldk3SRYyCz93ESaIOapJBAyll
CZRZs74CbUrYil69cZSdw4+xah8+0B/OfugILA2s5jMRsFWQ6ghKEAxbj6Zy
jk5qykS0Ao3o8n+hqf8iM1WanPOhiGOP5KjzcI95MYyb0vw/szf9QKzWjj/0
iHRDK7KW//dyfE4aS0ce3iWwYkSHQSIzGCE/eM4k61E/J4ao1un17r3D9o0E
0p1Ma4irUeAup6ua2uucXEKEnEModNOQgOiBLJgU79b4sv8BdfvIWo2WWu4N
LjQ5tPMOHRl5vGoa42SU1pUaKP4E1s6pm4YwTK7yD8wqzjkBRn4a4GmdySnn
m8eT2DevjcdLf3ne/NWPle9yvfIDTIcKbk8SAKv72cL8fW2G1U3FQjHXmV6w
0kX5+LItctdeqrxoFgxKA44px6AXhBAlrSIAgk5CEK2S0CIWVYVECLLqTtfn
aM/Q5e6Ik6bQeOxVz6/6xWqYhlkqyl82ly0DBH9YVALETcYOkyftN8TzQern
BElbUG28Uv83EuYIOQ01jcCY8OPHQk+0SQdoOYilLifRBraExBokWdQE1GtM
MgTcY/cZ/HGrpTuHkaxCKJ6eWFx+LCYE5TOp24wT/M05BI+Pf0XkeJnvLD4q
t3Doe8ujPbifSRUIgWU8/QyCHWqZHfVXqK6y9oRWuAbDxdQpUtp0GBPyng/h
2+uZZNGg8XeYXNhM2twueoHg0R8nsiaAdkJnYTL1dyd+F7SMHyY9MOIW4aYA
bG+A5ixymbJhJ15Iij8eD6JkNSIlTw/bXZno0f12qXwLbeQfyDIuTII1MJsj
rieYc6jZ3yk6PLmEIjrhMQ35t/cE4TQOlBZ5JvVb0DqaNyMAFauqSsiKdjpr
VxdiuPR0+8KXQeyim+RwC4OUI73+R5yDepxPthnC7hsfmD3mL73zWybTyP0k
flXljP9aIYZISbZEg9Ttk64Itlya6qOYQ+WaSAuLi59EjCEDSzkwhHxufEeI
3oKzD8u82YjarXZDFDTfN/GxC+VI7b3Aqi9ooO0X4u62T3zE7umtRs3KEv/6
RXmg6SI27hPJ7Nuf8khZTFWK1sdlRh7x8dTwJvbgCmx+G4NF1DNWya8yQlVe
Uhfpxj3bf77XqVlJBBvhBfadPH668+BbLASGASO8pmAdUBstFn1ezL3tca0p
xNnA1+YU/pphzUf83XFwRTeAlMNLqmA0i54IcQDWDfc2Yv8eECoDEMxrfIqa
0GEPD5AKiCy6VQQdoJCGtd+7p3miLbSQ83F7DSrOZVJDSPltMauZta0fuYaI
8iQSKhON0iVMB2Z9Vsxg2O7OhFQnvZoE/LlIeEahkdp5ZHzYMpfv4znCNQo5
W3Cm4WJgglFYxSqroeqXqtlk6APkKyQQLW91t/8o9SHVuFlLPUmqwN5Vqvon
FxdQqD1YNYLOrWp4k+WVWg+JvWAGpTBUCgCI0+5Eo6VyJ3MKxHWZzsylRUBB
Fo7JaYXb1yD+U8sPJp9AZS7bqcJDy+UeW6eNOMWikQC+TKXAUT8XIHGz+6aP
pFvB/q5ArBYwwYh+ppbK5qYTZNWoGHH8BtcWkxDkN8zjKmcBmVdnZ7dN/Cy2
crvYSc7A0YgsSKs0VKoqukGqZAqTcAsiXDtF8VMecvlAb+lzeqAQexLyd+ov
p+BJjaD5GDmpfh0om0BjJAu6x/KwjJNXjFZ6XsStTFfEOQb+EV2yTH9AtOdL
vdZ3z9C3R6ebut5VS2Q4tF/pW+bjKR22MOi10LyFsECY0WQyfaox4r+TJgAU
q+pIiCWD2ax/SgampRc3plt3KML3HpDPuWYf5M2LYKSPuj/2AmZKZhLSzBlL
EFZMC+neNdSnIzUIU0c5+6BaFDfGIKtYoWavLRv6xDE830gOdgoa8I0bcUmy
NPXoKWXtOyHHuVZ/A1nJ3iawy9QtYt56PXZp33MN8TIVWEo2y5FnD4tSnW86
ROnpowp0fsQpBN2bC+KhEoNJ1qRrrCH2c+U2WNmWl2N7J8TndN3AuvyDsXfk
vXJfLs5jgccpN7wYgb5ZS4IX7oxgoVzt6g15PgyjZONTDGjBIjBDK6h+qSvZ
/Gp4NwjH0mZuC20Mua+Lx6tWv4WXLnX8H3LfJnutIVt+8F7hQMQi4s991+BI
5Wb8ol67ATxKY05sCM640IPwaVC0fJUfetAqhYSdWu7wdknZuwKEie8EtVxf
351EJTF1WB8F4TId3RGoTNGRdGAmsexARDViCkORtpvIL1a6UUyliYc4FrqG
p2A9OnrDvLUi4MeU3xO3A48eUol7/Uhw2SRlgVF23fw1ZbmBOz9U3sO4r1PP
IKq013szlXLZWu2iTlz4lOJkQesZo++NlODaqSTowi9MRh1tquz6NA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfRghwT/w+TyiBD5y+aEwROvlC7xXvATMjQKg30JpPFogLCpqs+osAlMcBTI1mS8SAVlurM0PoxStkCSySniTPBgkmCEbL+7mS2epUh7//De0ASE7KjoEshwuvD/PlAQ8LWmsIlZ3YGWugSMXL2tjvh7SUxLYvHjNm6DxKwfIlsRk4lNIcDzVJ9CsjcW6ZbfqnCgh7gi4lPzlrV/JirzIEXsrDZcQ4PEjBJT2etD8Sdkwfss+9OmcJKgXKOWEe6lygd8llV6aJkvCT9qIkVbFiC6LGdJEojJf5SuYfLpkCdfnCcwU/s4YgHSXWOdXmRXGexXR6gTva2jMPIvMB+QJjInZ75Qs+qdH4lBbPdcZXnsTXVk39CyPQpgMIHsxa31zljEU9GsYNzqU9s1YauYtArwM5jtkgVRhzOJBWQVOknS94BiA+JsLmUYW8+Y+7PQHuh6ttLw5U3LQKYh4a/KYM9czfbFAeQTeG4B6NsE5pMs7N2A2NVlHaHLiQF5spbCnCLycTFD2eVaAXZSNgRFTSG7waLvHlNn0IZLcbrSQMfeOysnnqZtHKUuin3PGOzp67uFYZOrHdTCyE7EOAMJKPKTSyxi7dpfVJ7bFzsNUvMeP+AvqLd2YrXm6ecTJw2hplpGpEcTrUFz1FlzuFn56FAb5tqtTpweGt/Fq7VBGlADrWAi8x3tzmH0FZpRbNmu9OuLWUeT8fzpnKh2SKTx1zWnpEj93rORPQjLgRfyLHINJDv/CjlwVqK9PFJiesHOHQh92Ui8yFpDd0W4FxVVATnJ"
`endif