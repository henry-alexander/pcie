// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
sbWPjWq4Gih++FtiMrHEkWKEa6l5akyRAGg5nCGdu8iI+wxQVAeXHKsPpuHD
5TxiZEFXdSCMz5Z7YYa5HLG6TrFxbh7GqYwUvXcar4T+uNo0F4ZdnSCdfAXw
9Hyzzg27+36//K2QGGRkKM474Fl5FLH2AXrA2GkaN/M9G7+NHhNFFf4vdsSd
qZ9XaN4EIeDq5qyMWHmkAov0E3uCRfadt0r6YPcJt1eZEEH5k8VC635v4FcS
5W1ahz8B67Ar53S78YFv+T8jbgLNfxMyguxkZXCidFEZiunADHkFN4Y2x1Sl
jMYxTfFeN6eP2Flsfc+uJHm4f+N1lZeTTuxzkbKbhg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
k/QhRrAA958pTu6aNO3q+JMGEog68w0IgQXHY3oFZAxA/evLBzpNhFymztA9
jcyAa7gzlPrqWjqRyNWfeSlXu5Wv72en2NZ4/6ldaF6m1h3A+gRoCLE2ke7v
J93+i6gSNEuUz9Uaxb3lSaQCS2bQly0PDfmx+peORcG/hGJEaA4XFZnyKrH4
K9U/IhFKlsGM8K+PRiyzl/4p2XnC4PAgFQstUKP65QjVo1wYoZSVt59gjYS3
PBYyiHAQysUVgCH9Em6JVT4C7krH9vXhSzvqA18JNSUgd6Qe7SqSX3xjK3Hh
t/i+aHeTIQ5kwX76BkTV4FTu1OxXJ8qUCfMnvpV1Iw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
gsCMp3+0chvcX7XbxvtYHr02KGIu1KKP2LjYBOodNjNgqaSHQJWN54sloiga
KJVQm4hEg7keCsUVjyyomZIeY0JEtSGmWdd7li0CGVq5WDJ0fslJGKaWqbpG
oaH/ASpjWo8VibsPy/TkB7jOugs8TzjIqRLRqE0LDEF5S+j8w+GyNDcMJbea
TwTKlRwyyGA6u/NpaW9DnSLtTInUGiIo/bCZwJhynocIykQ/QuvmXYApJpvf
ZjvaGb15NSs4m3Q2cLiT4yqnEJaumGCbDeQSC4u20vnaSurDxbnFTY/WHzTw
n8Kl57sXIemM1ykTCvIgsJgG0/aXQ7pa8337cbr2jw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
b1lA29KE9Jsn9GMl6PzteiLwdzzyVlfn6U3Os5aVv2DXK+yLlIuQbTwJpbC3
RO6UHJ61ySNdRaOy8m3AcP1xZi3dgwREoJSQAm3sfyD6he/h3f0eXJcB77N8
UG4s4XKs4ZvNzydAbVI8GLJB594CyQoU2WcOLZrOtwJBwQa55NQ=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
B2nnrLw2Pcgf17ZFHUsW9UtaESW376HuyMwre984GOobiQcjJIILtMv/hQ+B
aY8S3PFZcgA4iAa9aJWP0gUt6U79Ek8rxi0ORdl9cP6VhDVBSxahiPhgMP25
sxWnLs5ViBBD5+oeYv5sPNHVni2NcAxdCLoG5LMwrd6wct0qoMExFX7w8EPt
enEysGeiOFRz6yJqD1NKSBTb6b2gn3PahSjC/LX1+qCG59iUTxD4UZ4O+UnM
Tg5SlIlbD3uaOIPZVaHle3kVMjz3xn2T4TM39OklXGzH24ssnvJzdVGCEbvO
VL3IjOmw+0JdbTXoVeYYFlkPzvisf51g1AobywLOb9K/Ezii/DVj19C3H2hv
Rb1IsmT9h5O4ZIjhsWdw2nz8cC5VqjMirLn+NcjNl/pyoFOs/75qnEOaTE6h
Lm38ZU8D06hK1xoltk4YZcRM0hQ4rlm+OaeyJ4isudmVNgxfzLY+i+MkWUwG
Pn/d0EF1BsL94XOxQ5jWRE3/ONa+CRje


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
mjqq7XzgdOOPUkP0csJR8/YROplbZ28XAFhIIBz0PSIp6RlsWXA1AK5lPhyC
C0t9QOvTKqh6YPFkXz42pWwpdrzkTi+6Z/lJMTPWDPNjmIcrNE48DlxWHUnT
TkYfpMJ26bgRk7reRvxCYUIxeQa/l8nI4y25ZcWHUsDptb77bX4=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
MpKzgIn9U7asdO+p2nW8yRVx9eaWXWOM5d+dNvcyrUmlA1W3PqMH8vtFWaSC
fLRo+PAddvbbsRhxGhhTFkkTmJGMaXvrLADQP1IZzTC1aJkHou6DrtAACVj0
NVYyvrRRx3fEOylDeEGdgd/zqf9PC6KMqEkhuO0ZW2MIflGqlc0=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 2112)
`pragma protect data_block
DJ0OEyHjW6gARf55Wt0/nTgtPGstC1/aSzvzV4i+PMlmRgTxnLK7ck3eQE2L
k/yL3VnGzIaKVdhHirAGpgDiBy6wXbol7Xx3ZaIPyPozGoGogNVDGwu1BeCR
Z47U9P1IHNpIaZZZv0DHXEi5P9OsYjrYwgjNX5h0cklQmtrY4j7nucSD5URA
gjvZN6WF4oCICFCLvEBSk9njzsTNGPKgNIGb/lusjrbQr7IC+ZZiw6V4DHK8
thjb5wN8Lw6bAOxNkKU95VshC0tUDPh7HuezVnUuCvJLIX2Vj88WBDUXFun/
wZzmQjX/JW9e+e8Xn6l6wVBBNyEVf+biecCYOdNzqtVZqrlKvPIUvP1/bnD6
QlOJDGih1EY5dVLA+o8l7jW4GHfGm/IJZYe0CHqm19AEHDA1w9nwxAjNwh5E
gBpjkS6qgbzDQxhaoY+1+XQo3uSSF0RyW7y2DRYLAu+qB4biIOyAmsp+6Uib
kJ5sAxWqOHTZwflB+5IRDcy9PaK10gZl9jGdv8CxRgl83H4GK5hGzdH2b0j3
ISqKLrHdCjuBo2pkvEMcgZ+UfYpXPv+nQ6sjrlg9vB4yP4RAMXvojFqFx0Xz
zYDub3UyiImFj9F22M0UBgdblqT3mmiLSTcmZ2bYKrl0FbopaBFNrVS8LtUS
Hw27oqC5xGqhzfrJD0wxzKRP4Xvg6WaS9kiCiNcXFIk7Wue5XrmtQZzsl5no
eqr50F59q13o93iQwHNfXilOGLOTqxS03SxI/xeKccnklYqbwInXs45uxH8p
/wDmObjrZ9WYDNHain3cIL6iS0Ll2D0Bs3mrUmlq0VpGmcS8u9NYW+6G2qts
83DRIKQN1wC71CLiFBSEOwfEDGpHPqGr2RkX/mxoVXNoiccdnayeF5Hz6HBh
ENN9M99l5ZMlNmsF8mk0pUQcI1d81aTFlPXIfu3b6lRqFjwFiBebMzfwxhIA
p7uKomV1KvjGRZ4/jYLvMZuzXvT2S1U4QcGPXvF3kGartA3kUhbl4VJQLEfX
Ft5BxCGhGzTpBKQugWZoNy5Z6x9H2qJm56zgp/vSCfqBU3KFg1esBXckX4m3
bumqRxzymNgMFaVEprbcIK4Sbu4k6Vsqo4oFhZCj6mZ8KXgyVKefSp+ocXtp
WLMWx0lQLNidLGAIzMQA6ms686pchvZ70h0Hr3yieyZf+6pTIWMw3/8fPKyr
i3Obe10knZGwkO0zO1jffk3UjcY7gzvpvvFUc0f6okC3yu/t+uMEMsKjXcmi
IHowqExdOdWrfO0DxkjmGlGqkUlxU5V/ja4vlHHEBpjsJ+JILGgC576z27D1
02LaF79un7SeQJuEHboRO+bjyJgeCqjcOa1U+v69VAFE2hAxnW3WWSCIXNzf
52DCm08Bv0mhq5ieYkq9RPYrvrl1tJbOTI+ynwEHMwDXeM9rbTNVDHR6ao7S
09lX/qHXLwhEZC3Lrpnp+WlBmkL53+9PiaiXmfXzAbQt5QGzwhMn5M/r34bV
8867dhh6Gj4Wj6YxAtFDL93Pxuy4iP0FwrromRuRXf5wirhrlaaIPejiREVp
oDzYMW+epcNjIWzJYecq26cbBDrN+Gy4Tzu+tcQxAtMs3x06eqUu5MxkFvn2
+Idog+2DOW0vjNxLTBExnpfSwPwXSysf0bhhvpQgnGCOHwMfzyCelzqLi79x
VK12MT9VASjyAsVCAxRSr0e1K86vqQs4NOyWDBhN6zxQnbXe+v7n7bhFEgwN
T8IJUUMsBnNs1iynmWd3kwpIKQ/5oD1ASn6G4e+6vFDJr1S73+kqT4BGAMFX
tdImNdJn723Dx+AVb4EJGUse+k1uIBldf9OiCAiXXOWKVxdJvlCzmaAGfdgW
IbtXv/VLjpMUdONL/1bpB9AvbrPP/9TAxujyoohRPDt7skaRC6hFEQlCfhjS
AkiSvvHkyNFEi/vtOgtgjQV4FTSjrL+2VWSUeZ72Ncusqsur11K81eKFFLJ3
ecz6aQAqvQROvd/K/wiK3w/LAU/npJMxL6NCMV3SkdglRfExK00AH8Ebo3z4
TmsGlvDaiIw71bRR109ayYTaA2NKPhrSxK+qvCq6RW0pj+nKnu2oCLo2GnKI
BGAOk5BkutSP3nMGoVre/08O6VCm/mF+4CDWa9chbOIgiqandPGkoPuMLQAl
ApBH/FY/gvV/S/jn8DYJqvtJYiEEaVlIRkEfDZ2KGNH3sZ2ht84s3glvxJ+J
48rYBeG56EkY/gOa+h4y/u6jSiPcu8PYhOoeKeIUm2milIDpmn9PIA6vXgOO
cqONSGQtIKpLXdwE4JcFfdCoNS2CreoPuBLDqbtFtvbRQKxCwCkaMkcNqEsC
0dP0IrvM9lBV46VAkFp2+6ph1fzmVNmpmfvg/+YbD4yloKZk0pT+vuVVK+Zm
/5HvGmwrZRz9Z0cNkYuVJyYQLZx/UFMT29Erxja8p1CjDhKJrex1yVomT+Ga
sio34gX7iJEOweSlMEuQQVXvxUMNsHRE3FwEJZpIUZfomRis3tDwuve80l83
WdbUaQxhPILcn/o5O6F48tiK8QT3Ub6zODQnhaoPYY4xBPK1B164l+yHl+Ib
60+zCl54NXX208zIA5G0ZqFkEsIUIg1+EI0F4PHZ0AVPnUPDpt4+pnSm8KIj
QGdEB5B5mLJWrlfxQ6DnhHhWZeufnU+2+TQVo9B9J/dUcKAuHrVKtBB76Wjb
sKjTQRL5SuuVUhdx9Mp2iU9FlFGCTzugcaRunPu7gm0Pg6Ma6Zok3DMh44qd
3TJgy6Qe3C2GP0wGbEHK97aDBd8588EWPfuZuxqXvumLTFtkIAfz3AaS

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3FlswwTRhNRpXJWPiTiOgBic8SPlPsYbf8IujKlV/2/0JpLQtHMAH+j/e+TpHtLFDy+Hv2h4J0CUMqtQCkK0eIdMbWaiSPh+iv9zrbCkjX2ojnrKW71EyKmAbZwtTpqwqP6tYWOdTsam6mFj1E3MFWJU55E1CT1+OpVYEZ61P6wyf79fLtXR5zNnDPIb5dab0M5CaZIuENxLwn12UDLkr0zJK1bM2Cmm79dG7eWKpNpgwrhFKT8wT3GP789RGqSC61UAgjbFxVyIfUjLIhc+ZuMNqPVBBexWKtWC8xYeYJN9zHfpYJkjGeqCnxujnOLjm9SPy/A0tl9NT/sDkyUxekOPvUvWrZTUV6smD1OSSYdXzX8YlbgRkTP3PcWnyWptHtr0xQbwxaemxGY6th90b3aTMRwsjLyUaHCkIBzywTfP3uQGkCs6HEjWysfgUqbwFSplc/6g0KkokPoURHY3APLQKQut0MvQ62wOVBQLM1y1upQwM8drQMGnk3ST7votASR2gXEtOPZ8LPgCNJcnENVZ3D0oZXkS+zs8njrgwP1UW75JYYO0NSbUTQJPwkm/jTXsGzxvVo87HIbI44i2KdmHm++Q0xm0lbFKltyKa+hThl4l9JjzWiu+xrkDSp90/TaWIsztPamzkrFVdmJfE0+j3TekE63eBuycGEBepaQMjRid+3n4xQWVCrLLRfYfNZwPLgxXGhKKu6gWG5bpn3NTXi8jgxLhA70ZB2x08LITbbwtvEyPofQDJh80Gequ5CCmObGQ59q9KMjHjGIaHNE"
`endif