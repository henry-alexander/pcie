// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
y6QGvV96D8qOj49hoh49Wt9mtKtGwvRk13Nho0rWWKCbaUsSyFgToyB1REzP
yyYlZchkL+27bRN7R55CBhMUKcR5ztulckGdO9OU5QDrQZtbv5d0cEHMvIbK
17tkQtaLyLZF8LmrkfvpBjbxetiyljbtiGhbspbG+HD79e/Kxp4kwVlHKFqE
zgZtUplu0ahDY5my3ctth33DwFE5IBRBGJqrkKTvUb5zlqhmdpo4Oa65k2Kd
3413+bkuGVXw9gXw1rtqAveeEfxomH/GWXZox3gVhSEWwP/Y4NwfL1QY5hCx
ZobZM+og99FdBIoXmZU1KsI8zLPUyTStGDmx1fYUyA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
oWnYSJq5aegfl8Td+qj/q8z+JCAwJA4Jdr9iLL0UJEkgANxp5eKE2DoipROd
fADQOQSPDyxFPqCSr4hqpFYFdrZIJbmp3ZUEex4ncEGLC/paQ/eKaze/71Xo
GQ6suaBzVZyQVheNd87J1bLXxSmYBNo8gD6xVn/IndHveYr6XfVKAvrrHNQm
Ig00UeC+mfKxnZ0Buu9dIxuhxqoE3zFoYFvQrANy1dxKW+55T8JHRp6sw94v
wNeqofzFeKu/Io3EF8kTNuiEL/ETkP0nSGVByesna+1BxpjYNS/AEDFvqzWF
p9kRLmzvfcUhv1kaSlWQxjdkCVZ8X/jrIKa9Zyg11Q==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
XXAUcLkQJUUxMg5rrFsqVSt3OrajMFOX4acUY50XKlqPs7ebzvoL9I1CuQ+R
RReL7YcqyMBesDrL3OCdeQAlcLy3wH10C784mJfBAAk7YNbP/MBnWV/uX57z
9uHu8Vk9CN+R6wl+dQUHt9yhiXRPxxSoRl2qqcXzS3s38xJ6LG4kOHyxqZS/
tRlDwuRdw6bhoLZpGHnIBWwyqxIN1KL+jFffz4MAP500nekoeFAhKt3uLiKK
PFJQ9a0CDNBAgyN7AWLBX9GdhjQwKui1+ZuBbDiB8C85GPakBA1PetZyZDWb
rXuugG1h3zbVUnSroVYYGga2HGqZ2SE+iwaT/jeiGQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LEuCQOLUVdh/6pGeUoahpYZqCrdY8PVooTP7ha7jG1G4Pt/FfeEQeghLTVHX
fu/eiXeLJQsr9F8rZOkKGBN8FPAfYe3wWAAiCQxLhbpuRfv7FfDIEYEk2H7u
SIPJqbNyLCPkSkP6Nc0gE6jDMK6N6xC+PmQFnT7J/q7veiy14tk=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
VZiVE2yGlGwxR5E9rIGlzB0uAWV0bq9k+o3a57VxiQpeTwJo2IfgXVVmkf6m
YNI4RKh2vdjcC4q5g3kYdA09DOcemFe0DQI1KsY5aPoR28fjI4u71F7sMFq7
KleVopwTENde0xuYIh0mSUzItVFY6TXnoMPIIzNLo4GkgncXncead3tl+4qN
oeld2f4oAgS2lGBCEB2w5hAgTcelwS4gUNWxBnecFRU08f2KPm5uyzOv0uFQ
ZzoqD+X2dVeWwAHSho+eghYIdir0MDbAs/TizUceGiFM15XJAiKemzkxmtoS
AemtCHizRWM1DXcrGL28pqXx1anodgWYIZAWijtFHS3YVCuHTtH5rflCxK5a
UQ3qK5IMf7xFGyvQjninNAWy5M8tOmQ1qAC6pX1/kjMXurdyEroziS0kKVtE
PJL+sf9Ge09iEv54cysoBXyTrbvBx8b18Ogg9CQPTId/EY4T9VERb65IXQfQ
5AqDFTeHfqqEEAE9YW8MYBpwGF+8rcjI


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
JQ1Liqzblsh13J0e+iNBWye3jEEBN88r8JgtUSNYqOH3K/8XTnLjbUyZuwP3
PGk8eeASVoguZkkkQha+hDF3j1eK/wmnrpHRsqWP3QVpyIgLNzOM0ZVIu+PS
tyoWb9ciVSwrLKFSWxJmzc68ukuUTAx0Z9LiATBxWlOI9e/blak=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
qJrUjgPZRK0rNwOFxB85SalWB0GjagPYSzSO/7oUlAshQE2HzxPnElYlF2m/
EbdqwD+yrmhV/4znun8IwUxBGmGd7sY5A1bnZiMNMv2OTshMgbOk7ydofXvg
qeYxmCndYJ1DniX/R5khPzyyHoef6YvdbVrqMi3b9jdfXKmL544=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 60256)
`pragma protect data_block
Uf2Q5HCP0PQd1ahKUnc1IRDTNf5AcsmqEGB9+/xWdGaV21bmGjKRkqZTzt1m
lakkUC0+Ldw7Dp8AmBN/B+Cq9HxW6LnzIT6xw3kqfhiyBHbVTqhNxxjb3r6/
JpM2TSs0YtZVjby9mFtsZFo1YWljD430dkD/Px2YpfjSl92YF6gsxK9KbGTm
XoUh4ffcE/v0VVU6JmV2lhkZQpSptTjt2tlATd/gIO5wUkF9YY88hguFEnni
2ZOWmQ/ty0keKXj9/0ChZLG7z0Amn623GHL+IZw7yyPtKpYiX3h6nGJIvpRE
+VZfUc52xva0ix7rqpZw0d+1dDLVgSnIVKrI8FcV4q/zzq+S7P47mXPKHMCL
XaMCX2ll5KrnhrP6kaE0rJGNc79ovohCAxuXTk1YoCHzQJa/7PGkcXzssjkQ
5APJX37JyVCocCZVBPTxVbL3+mRoQ6prsap4BjDk9kB9Hvk7EHwE983zpdxA
0/TjIKruRkQZGWm8YRWr5F0iE/d00UP2ZIjGE7pJJHYAkViXseaZMvdGjz6R
EVyIXnxpGndftkinl0Yv9omY419603isYa5AKatInUNzViF5sANQk+HKOIAv
NAveRHG7wxlOMWUmCUs3FoaTDoXobeAOE14b+32d2bim+jySmD4y1JjMNSMi
DI/K9UZFxp/gedLnozneQ/K/nwQQlqHjGDngE78X5ogTimd/gojeiCIVJjJy
RZJwacsUzJwLwKdDKiiD2oQQQhFoTRmCmcH5oKnjxAkjGs9ufvd84rgO6cJc
966418Rn9aOGb+Dbkja25ZlSeZIH1BUDgwg+bo8aU9zCsaRvF3SoVkWQhYNO
n9vlinuE+ZH7IXN1bNLAne4HyRLLup3KXi11Ih1fBLD6xM8W/d/KOmdqQPQ/
eWZ86BlKsTc2JUAaJZlvAU5LbgO4+a/YKYY64K1yxUSLbQxUKP4zZ72K2Vaa
pfS55hma0yIfWIsaXMxbaQwruXAYw6nb3mhA27ddXc2Yc1S4gte3/fDVkkqz
RJrIh8tOZ0gZxof34skjezpTPIkKnMLqM797RG26G/O/R0UdTd71BMfOSNIB
JjMSzK647TPlmUGTEov/mUKXCr1UQcU3k57LMR+eXDDHv/O8E4fWFYgUgeCj
zflEOeHxw4ZRGeVZDx8x9xLStV6euJY33dnZvBJMhpvJ4h+tOn7kVG4JvbY1
OeOif/kAPxECZSe4y4Ynj38gCZyLCgXRol3oKStEbCESiKSBPXZML60WklU3
DdXkoiptJL792jFCuFq5kOwx6aRbUJxMu+D+m37q3Jr+MCW6RLqFyGTygsiw
wQrzkIbXJbm3eFIaZj6/436X/FtMp+Nb3HfiSDLpzlB/wocMgpFX+E3k/IXr
LiD5m6oYOY4UgysrrhFWxqaWIF1WlKvK0trux1SzOPkPOJGYWC7Ceggja0im
OPEVUUIwExOOPDO3Dr/DTwLpRyOsuIm+KosAlriK0W7h3y+gyzXYofcgS6bs
a5vQ64e+h4hWj1/X1jWOj/FXzpCByj41+deVw9T/5jM+/2UTfWBI+w7nVoKq
RTGNchGxTDZrVPbDoCqhjo4nZmfvUhj9sUGaeooxHP2txf2OmIJtjXqi79N7
PSuCvu4Am0Gg3krJdoTk9RxrNwCCWZ1Z5EaEyeyVzX32yFsLN7nsCexSL6f0
BwcF8127EOxc6vZzynfZIKU9OTCyq6mnA0GqdXe0AmpbaMkhlX6z1QNwlscD
Lweg59tD7BU5l5lzq3rBsv5KnJCWxb0Of6UJk9mZY3Gm9YEsJo3zyX1HRQog
atia0kByORZbwgRlDFqasobHx5wp/gNpwsihneq/87sbfPGw0sz1QWidutRN
GVHGn72pOZn2zaO0tgE0+hlaOmKkVdBzRHdW8ya1KAPrip/CJpQXQNrb3Kp+
OE5Ic3lG2fjcu10kg0BuBtB/In9Fb1C8GLZr2TuqTeCQw+TVVWSqiD1hYgNN
/MdVL+5VcO2CXFQ3YlFrXwJkjZUU5T/N6dm/7flmqEIjj2+V4STuR8cv5ukE
yHP9qr7bgAuBaK0mQJTau/aYLSaXueunWEpUKJJMoVDVIclJ8NlzpmYpblPt
vCdRIJ9lg+CAOWEHXNJfZOiaGasNSSfavxCeDw+XXGBraYHXbpShmOxemLVB
kWCvuNI2w1vRC+JAy92y2rUQSyCW4auvEbuKEPv4x1tYc+9REsSQuHYgTf8i
bqrffpnx5n0x3wCr2YiiBpfplyQQq8rWerGBJ3HjlNUy7tNl3pl/oHD2diTI
lPzYZx0ETxwrKGmtNh1bY38kEGF/8faZLvKDD0vmQC54oHcV8Gb041KWISYc
GYgkPkpdsEWO4fKjiJnCJcNMF21YmYFWVSZxVH3LOnZMUGrYEJUu2hFC3PF/
W3lXGIrenL89iURPsyGc7I//uL3l0WpZHAxxZz0r+a0w9G6HdKcNtk89tDrE
5DhzIA7RhNph+UPfylg07P4H2BU9ZURJStmIVdfS2AUAfSbK9/taJ/h/xyd/
6JUgTjBms08c2kF+mDwCe6swPc5jVZ+yIC9GlA2L2gEp+dpk+nF5ep1QhgVZ
ErUtNZ5gPBgxUNvuyWWhmYgR2ZPUrDyS24cakI03zd2YXMY/DinQtnOJwq/o
R45oHQIFlTJfZOLwxrzj19UPHdRaQ73hpRcullQTFAW+NSEqUnL4OFIIk038
LbL535ORwNrVNQKikFMhbue7M0jBpqJiD9uLRiH7tabE5K+Qv9BOY7uJrRyi
WyGwhu6acyCQGTavza7xa6zZ/0KziICDMdylDYPaRwbpirfadYtbc7BMN/4f
zdnY+Oz4DVQztHsc402eWoN9slRE/L9ZIt1/4tzYQanXAI0sO1o8rvQJX10p
l0z96TQaC9T6tcAF683xSaSMDkUk+RYcn+Y/pEprmVHxHEQynF8w+dT2R8Ib
zFLyP986QQRa02XEE3kfabtrD5lj0xl0hx3oPsSXybpoN2at4rPXe0UWkJsm
hl9InemyCW7TwmjXXDrrrgbsmJW/iolvwcKRxvj/B5RhSMXoPQjkmXyhkTa0
i99UAkZSkNeL8m0ekHsXdMZPv4IQh0y7sWTkSdzQ+VHar43x4OCau3WFdUQP
GPfGCDCJI3a5/iLoFFhGlTMal0SvNvguzbdmBh02VYRmh/KQ4fAQ/5pXia+D
Cs8IbaOdJerhKCAPDGTd7T7qT+PL6OWo4cDn88LQy5SQ7rpuSjmTqzYvaeFc
buXoG13ofliNowgJub1TaKwOfbk39vNYeEYVAywIIiNRvdMnTwHdrA/uIA3h
cOImL/HxZQzL54o8HGVcYpTf00k+TvEDROuO03lVapC2SECy8aaKfvOSxG2f
fblzESCuIQzj6qi6u7iRNngzwU/X3plMilCsgY7e//j/1Lbj0XmkjHgQKgDe
q5LRFGDzkW4U5h1I2wwIwgcSu+ZG5HrqAZtA16/XEP1rGKOHtXrU2L3b4Kvg
GuP2QmjGQ6LIs1fD4p5ujuhYlcY6NGVIsWXGtDlBjn0urylI4Nk+Jk6kn9H8
nYOlYL619TjvfejKLRTO0kbcDBFSGF2buqfCQJ1TdWptjLTogNGnkVxciUt6
xauynzg1bNzWuYPRq4MM0KEsX2tmkHw6+XpZEC539rtcyqljuB9wh2pjL52p
nZ0Qs2yK4QknGdTX25RPmmXzZ+zffbuUvAAGG9y4/1G/NBvbLuMMnvcqBe4v
Bs4GuCITfkDee85qQWyrgA5UKC1MXXYNFQIo4gcMGPhF1T0bFSKDcrpY4CKl
46RkDUiaKT42pASegMGeQ8lRBTZVq5FsKgJuqUpcDxeSkZso8e2+pPvI7T0u
7yrxxDqVQk8Uwc/yQaA60Bi5IruYBQR6fPsTEY1T6tqbKRbxUa31AGOYqugG
EODnrmzOR0WVIs25D0WHq6H708ofgu+f/Heay5acdSq6NMCwyEI6OTxwcHIe
mDQKys4TkBQO/CzFDn9BObyhEWzsuO+qdgUT2Oho+qWkXpZ75NqZFjr0FzZ5
1vEU3maD2aljjtmnNtn4CggL9LEUgO8RVTdrVEKJhDuY48DenMbFYm7iX/hQ
mvnFEUZm7gZ/czsOFQxobRuo+U0tOm2R5rzAeVJQw5kDfUYVaoogYZMr9qlf
+uLqHBKvaKk8SXv+gLDciKu70mSJcBCyWwHS/3tLOrsDZQj8ffKW6rkS/5CF
YLgcAVbVEAqtqWjjr34LBwqKMgTAvnsSumA028Kt2qrxvekiXY+hO0clX0X+
RjuaQqGMUdHxleJm3jbf1E8bx2hFft1fBWi1JE0xQIdnsXTQ24thni3gZQLI
IDIlwgK4+6gTiB1Tpz4dyjG8/KHX7vBzyw7YGs144vvUebBP2c/s+D2CKATW
OAhy15F7TcAKGM+T4UxbKC9Ao/amPhoXEULzRYf2nn4Pe1mdP5v7ou8OtHyU
f9F0KWlfDDl8QQr/JTt9o8TkKIftED42imEkAFiVNxz0RPtz1plgZp2cnn7B
kMkL79y9uM8yeCQkuNq2tKRoFGSkXN6QMEsJvJp4L38hFIYLpK5aDafirEHk
IQZBH3uQXw+u4Cam+xS3XQexTVlf1hVlUOIkqVjkfQ1gRuVMEG2Ia//VNmsh
0o+EU7IlC6qeZiL+ft7bT10SfZp8asmqOaeYQ5BKHWj9fgU5JHXcrWcWC4O/
kBXqKJ3aDW+TOb4SrZqI9knpVjptD30yA2UCwFQbZ4mDNx5xg1UE66CRqJMD
5GjPlKl8q47wxM/7Pk6pnRsMqjtP/uak+5Bxqb3JguQbX1v3yJ//BjbKNIAv
X6yjjJZfoJObHb0f2ywokpHNj5uVXfDQyG7pjJzrC9e7pyrIA6zaK88btcSE
wJDyl868Zlu6A31A/fyFC+LDi7UrYs7dub3hWSZNZf0wtp3xT+BDXxpOkC4Q
AmBtoJLfUHk4bOle7/L8Yq5LF/2ubmZfcUOPxMI5Bul6h0yQjFVIQmEogRys
LIoXRyqimtRvRUoU2j/lUrkq1xJyTVTKMZvt/axYMe2N6fLgNv1xMoe32CCJ
/Ap4Kgy5YhXrhJMsrYp+rlocx8vfR3U23zF59bOOC6GcOZn2Sb1w6rsKUzjY
Y1IRBfQH/z3x90MtwKO7FeU4uQzCprSD31tgDsjUTDWcQ5yqZJItOi9YoTwv
gSX8FlrHN/BO+CDT5zQAm0NkdhIYpa6sdsxSXk0bYBGbc1tt55hJdPBIJbSu
Qt+4W5CUBbUK1a0Ta8LByx9C4wDifiUmpddTkCuafOI/YaZUVrU51447Nlzw
uyB+iuyJKfxp6AA2vvefsF/t8pfV3lde/Iv59wpPw1AjvyWR8J5mugfeYCdN
7QMkh0pE/ogCrXlrzhYg4ip8IEp8VcqZJ+bNwVrPIprZIb3eJ4CK5nsbvqpC
e4uwVHmI6AalhlM5wZVoLSqOGxmH61mguldIURH9FwwoS6yudfSXLKIVFcay
22T1razX6IQGD1nL08syIfn1UdFvGis6AvNlXw1jZZs3rPLqNOOC+x9OysPE
Kcht04n48W4+KKrmw11uaTmCe+mujR1dPJ+LgnnGcQF/78IPKfGrOOjWiX+M
qK4OJdkk/4HAiCGVm2HMOEwoinnMnqzMSs6Qu+H8Aml7YQZpOALGOW3JvwhW
6mtjrdAu+P0B9SoLm2QTlFfSsOCCnt7fdIjSW0etjyVsLlNC6jg7k2H0qISF
29HM1WOUViAMdK0P1aj/GLZXQYvaupX7DHC70kebjU2Sw8+hyPc+SxLLD1A3
QhOk7bcIAp8B1v0mmvkSTOu62QGJgH+Dm3L3GhycxT5RR/D8Bb/4JWwhxIqa
ctJSK7ynSuxJBofWaThPvkhZzy8O79SLDSWrX1GliV5+EzBlBgDovfSbeF5F
6P4laUQEJoMUo6AjfMVFbcJfEoG11Opqyo+Ux2JFxgQ9/kF3mQ5meikFLAJ+
sHiwV15sUzq5ZRYy0vpEIrbNGV34PqeX7H21lVcweO9cUfR1IAtGNZPsx2cz
wMZTET5rB5MDuTdGLjYStj4gE/037NC1TLt1GA91mhF+eXBFd72gt96JvZcJ
L3of1KAKw7SicixlsQyQAft18FGO/jeQzBU1x4aygUdTfCorUkn/dSIXjDqW
Ik7oIWM5Lj09NvuuBsWa5DkOGAcOr/U6MNejL7vcm7dqVsrqsqYbMDwWZ/1B
97C0wYoddY0M4M10UGxNU+vA6oMhN7n/565QOBJbje+O/QkVV8z2EL0WvX40
36/iKIFqIiy2xYAaAbqDTd8Zz1bTjTgvnEi0PblqXjz5P2iE7qPs6/nkywmz
0MiMm0EmTqvHQpun+TmnNFWRnvHbIKk5HTmV0CSILllR9/bLJ3DN+G+HWEIQ
GhhVrxKPG5b1OHnEX7WJla6cvDE41qsvuStYdrsx5t8nM4k/WrjDphW6hOdF
+5pRYUM/XOZHnYY4DbtqrDX0z+E2vE5+NOemL/LgGJ0sr/ictx3aU1A7WM93
v5b5O9jHGZ6unL4QsxVsObZmg4+VZvVJ7mw5KGmheH0QHl+6H5AdIwm4NLNn
R78S6bzJMjC9rcdlLxZyXr5XEuSrwAjfVuVJGjK1eX5twqIG+rqXAfDSb+8X
wDH8AoeSmbJgPV2ICJwTbPPq0zHtEZgIzmMAv39Y089mHQoDTHfYxcgP0tdH
ys5XM3/P4+d7KeMqZoU2bTFhqLs6jYJHAZ5NYBNmvT6PTke/vTZnlk0C1o5B
M36FyKIEZzBI4Yo9b4GApS3C+QXlgpcN0Cs3fEbqzbhSv/b6BO4BVXzHMrNp
jtrj0y5tozzXbMGOo7MaHY7UyKf447gkWRrYyl2DdYec9ac+HKcEv+p31I2p
pffbrL1+j2R+VAJPp3lti/o6uxsnnr8aOq5VOac0RWhIfzAlCXXTNUrX+CMF
CGhjRHWie4dkXTrQ+rmBe5nW+2kDbqFQfSI9E4+I6QTb51yUi5mcD9D8NGwz
xsue38QiDxPHTVtwylE69wxUuMVmY1mfBIXRiZWZasUcSnnAenQfW6tHETON
o5SVzFy8WacNbc5UXL2SpUfR1+eZ1Z7168MyyjCO5Isc74KGJP4XPJ1G0SvZ
4ZinYCxxsBryqyu4wLY8s6im+/irJcETspatKmMWwqwD6t2Cv5Tm4Bdho9UK
VbcykYAswoA6mG0F61Gcdi7W1rEW5RD7wJRlbEn743zcg9fiX80+3J4zVHEj
X0t7b6hhyb39Cj2E5AKsaQqSQvirbIqLQOGyAS5ufmpk2SShUNSlZvvutRZQ
RI5Qjlyct2H2Qg3H5xjZqBIU10u+4iHKXX0rOBsTIvb53X/y4SpUusXniYES
ZxTOGdENQL4yGDADRGBrDeRZCxy5EKWssBUo1xEeH0KciFe0Vleu+y5l9LNM
9rAv8l+1sqD/GqeRfjIqYYVoAdAjtfUHL1d/BHXKf5xPS7oZr0GSj7euD32j
O+oTHssPUgWeFrSS+hyfMgJlrjJ4maoJDSUpgZD9V7QOiym7MvksEL1IZdrE
mwtOyWwrHifodF1QlchxMiTs0E2M3mcijeARk58+4ubAV+xkgp4PvCVJecQx
e3pugutyvusKLjD4ju2yB1mCjYnJvmjOaZUIxPcqrHyTd1PuSvNXAob9zuGM
H2/dNRoSitvdQvxhBEo4rfhSyrsnQYTSCezjM2JAsIF7oVbEKSzGbOEQLQsv
UdESZMg1ZgVzgs4yr6h5z9XcWIluRTVLABWmm4eMof1kDFQ+TyiqbhQ4BjJj
1tFRi08KaW+Ee/pSO0KMOIcp/rWQDkqhJJhCuJtKe+kQxCgbMpMwHr4DKZLZ
tut1eT3MwsPFlmVILvKJ3UYzkbpXb/LF+27yVjA/xOdwHgzy1nwgwuKMriPd
HG/20Ddjj/u6NNXyO28UOHQFFLcNLjqC0zrbV9y3W/LY+Rq6eqE0kPQ9Qc2p
dW/YUCLU+saoAZ2EjweBscANtk62j3LNKDqZtLSQ+cuWE5w/X5/f0cyjwFlq
zpXQX1KXnGCI/xkaD+2oje1pT6MF9nE22fnAJInKIpr+gbYdcM9R1MwdyHOq
/4ODZGo7irb1CpB0Ym6/RVo8+GPsk02lheLMRVrk6Nwnmikgf+/Iu4hNOTae
HRz7U5mwHnnTnnN7lDIw6MsZdS8CMSd9hzbQ13bqtovm3t1+lF5KO9LrrSVl
RVHETr4XHVz+8kas9hzfRIF0JSD4qdpiEyf+eRksFurUK86LpFj9/H0+ZaCG
eXjuQV0ow9w8OgJJTDvaWDojK6zHRDkubnJMYH3ZIwwC81sZyIBwHREASRKH
/Uxg5WDvz7JxfLVUeRRgvRudOBzFAoIyaFYng97FL9t73YRlQ1PA61NYmzTC
+AxTWZO4fkbsz7bvvSLIgK4zQzG6AZJrXGpTDiHhpZrt4OqbloCBbkl4azQd
2kqmHHLAvYVJ2sADq+GaxBerEpXbAzIpUVC+v8aWsAagC9vMVU9rclIzWjO1
sl3cHdxxOIaiGPfS3j4XhXQLMr/YeD3Iech+m4F79py2KJw7GjUm72J3iJrj
YTCqam/bYyAtmVjKo3iDHU45OKHevaSDa/h7BIqbR/Zyt6DG5JRNzDcRb4u/
neL+RlXeFxy/W4reFM4WmInwmZV/b/imufA2GOnIpEklUH5/SlSL4rvuZMGZ
Njp+JZuoKLz4C3kBuO6nVgQlajbWHqwv3n1v3Sm9EEyJ9nos8tZVqWLc0Ttu
Qw1oU5QgA7FV1069aNL4RCXSIRkxso8FqXNgdUVCtTF80DWMrfsVsfNB5jXt
ppWcB+zrr9YGMsJZJzO0WAHRmZpRIoI/xntJg1ByiG2cPl7w0lTgMBha2ZpG
OiZfpUjDfS6bDnc1TA7tmu6sr6licSFrdOWRdVpjmQWDqm4JEoKmBBGEZhHF
W4eBCSkhE5ysaoViF2jPY/w067H+42PwJ1aqhAlGnqgMTU3z7XWkn9MxD36U
E/KuPizqcfW31uib3wuf6fl3Va0a+gXPGH0MUg+GqcuFTo1sGUYOIrWD4eEa
7DRcS3H0zb/gYZOZnDiHLfNQfwWQW+T/cr0Px2tElkJITxBbEIA6zVOfeAI5
37M9oq3f9OMnW07D0rt7JHuHU/YNMMnxMEjLEndFFdRL6rKo3RkR1jag7sOS
+cx82i8yO5TdiqX8HQJqV3BGYjbU8ZVWkkql/JtVGa1y2BFBx9FYSwn+IB9A
O1uEeuVAbl3EZ3SkEWL+k/z/9uKllWv18LFsBZ0YC2vULAbyD1ICo8aK5vS1
4TMe5W+FQmRTa3R3dxKtt264nAfNhLISVcRQMovlzTPoN3oAG+8a59ouCZh+
gZ7bzHZcyHfOO3998jhE2KUrqu/Hl4sSeNSaJbH8DBDyZ2FKPi1cwkgX64J0
WpS5pF8zt0TXtuswzpQokvLVwFLpjOjUX9HmfvjRz2M9kI4Cu1wOFXBx7Ph/
6oGb9YlCjSIM/X97JFX5fz/w3KUQ7GAPnGhH1/xjD5iGXRiVzLvM6WpJB/SY
CDj0EUn2jyBMy2yqb8dISJaXKNPAmAUq5Rc0qkEXCD4SGYCdvZazJV60UVuw
ub7qR7EwBoY0dFnrUUVEKuEq7Xjd+HfFlKKFT8palwrtJu2+VxYlEsW4kja/
e5xpySbZXjOW15Yb+CSVnB9bi3icqbloRlBxU87HyI4SIRL5cnEdMLUMT94N
yE13cnGGsfkhn7/nYgPnUbrk0HTuf4B4xHPk5g85k1n3EHqmrzoowDA350YK
ODkw+IJtkEm8l/y7UTml6T+hJPcEZOyuVhH6+QIECS50KuAf55/lPtAYG1UK
2IG+mvh1d/eqth0yPddtAG2pb3Kxc1tCAOT9Tw6wr1w0hLaQc8QzJasC1bu2
oLJZ//vM0yx9Od0Dit6tV7D93tuXBrX8dd1WcbfrKZvFlsfKnnSCHG43CFNU
MwNFlL5B71hZNS6o4VT1SYpQXu1zUcMVjUu8RMCevvcyFt4KfSxjAZ1amM0A
BW4Cs0c6R6VZieXPW/Pr2L9SLWEybUmI1/yPZk1BdbvS76n5i5ySwzQH6mkP
8X8TLkdeWs6F3jzIhKwRh7GGika1s3bJTs8dmQOV0ZdFTN5GXBxDWPPKp23z
LPVkG0pbo+Z1mLGtHC9G3jHpxG/a/3VcZ4rWC7SW/ftXxC0ssRjltd91FeYe
DR9tqi2xGj4DI6gE2wTPhAiIvX9Gx+AQmbcl31RtT/3R+QrrHZJqmPKfGzxI
DGGdwVRGYXhRqm4zKqJeekESV/ZUiQbBfZGBcbhGxB0llzJJrEPUzTBnzGIX
GdgM9MvR+InsHMF+UMEAMdf+lwWB2dOC1BdMLbji1pTkK4Zu/xoqj7t3oB7Y
HbS4uYdiGfTGWRr2VUyxUxaH1V9pH9qlloeFueN9Il8IxAP8pYlQNtwwfvyS
WDqFGxwijxslZIRkRx0/2Wz/9VK55/AepJDC8mJtcHK35BMNaYwNMxy7sHOx
JRjgIJTacdZD83SnyJvxCNacKXrBSDDErMAB7X26RP9x7Qq4aC7EWsBffW5j
RzjADwTKZXw3YbcqdVVqV9LzGtmN7tYpXYNbTyzMibNOT3WSCaUDKk7k7X+f
Epez5w10JQzoXy2epocHOU0mCROdP2ouPczuaVS/FFE4UUZSLsfz2QVrBE5z
S8EZoXmfGegVs317y8xLdq83CeTMcVtH/K9MooVZvHEw98KgHHerFu5n+IGt
XvIytIGDGcX0mBawmm5RSlrRgu6RS9nm8dWRhNTNWx9H/MfHokoyuF22FY5i
MiWj7MB0JaGCA3A5+S0HqpPXUS9n4NoM5MFMljguKbFxPAKFDvwPJQkzk5RU
P/d4L42YqRotDsMbEGwISfgFTez74GTTKKcSe9nqXCPhTsQzCnj4r6x8E2GR
GxGzIOA++wC0g8tCBb4N/oXWUNxvJsOWLd0SgZJW9YOhwsv4MJ2TFwYf2gXY
lksT8bnVmfC8XKgINigIounHfJcAPemrLWGmuMq2bMF/FgkURpPsLJeYKC/L
OAOkhtFlO96fv6FySt7g3au1cIYMimJqGgVi3mPAuOalUBcG1gvcOdfZC8k0
LEpI/6XKBko/WbEmaDMod/HTQ7J9ItNE/oitEIzDGrBMZnFn+zM/IMQCEtI5
vECxuMXPwvIv2t+56L+0gLnbG/2utDmZhnM+HwRWkQvIireOwhGtiqNFGz18
0X+oiDGfMjOVNQ2RmkxoVyPbhMJQIER+jBm9sVAXQFb9/MeCZ9X86GxLWtHO
KcHMSS7/BXQP1xORYV+pjV+VgMTefzoM4+cCUocEylTY/2huqTO25E2KZCHL
CgM6rz/F8RCnDsF0pFMDiD0L8nhMkFAz7QiTwrndA9FL9DTgxJIlukAg6Qub
t7QMlHlL7HrhHZ/M9mBR75pOwg+mHrccNIujRH1wQtCE4c3d/6rH0oJ0O4a0
Z8bdbUziH6lzqDfAxh+I0Q14HGJGOrajxtnxeZDyqars0gNgGvrNoQ+ovEI/
X+Lah1y/c8K+0YD3GgJHrxclIAG409dv2pr6NQ2wnyieLgznDV1rtybE3rnQ
7Tb6u8vnsIaUa5FGP2Bz+IamYUaXBfDI9qGNIiNAe3YxZ0OnoEBV7YzhUGAp
AznVbmM9Dw4Kbe2O0LD/MWN6XXrTK5E/zgBn421ogXI/adCTUzdKzjLUCSv2
8MhRB+ItdLo9iee03+YeV77RpZs/HYjt4TAonjuPFHrljnX86rN/iP8giWL6
q1CsecBxLpRZS8bkXQTVh1d3XzNRydB2Pz7yDT3sdjUzT6qIl9yUuxNW60wl
ER3xW/JMrysqIJNHXhF1u4ajCQWHhusFQlBHX03GKCbCItf0zH+xRKdK/Ffh
h2AJz3OYVQyD5fmsAptqLi9SRzKweiEQuTpkunLKBq5YmFzLzS4ubz8i8yjM
g/4vLP8EmRIv73cxg0y6J0iD7RP8mT/9FFe+nGWhzsFTiHjB9xLa1w/ZZCdT
/C/Hfk/E3dOzD3b7BdVPq24ddv6GwZpNUWaf9oo/S+CHgGcxg+wnHoj29usw
v3vttvMeIMtia5cqkPUyDk2V3+UZexLCyrkA0MPPUC1LxRYsvDmpU9Xbcbs7
uuS+Erm2AxPftluyhneIcjkYXXQASrq+CBOkHPgnDUQRsGQaZyYdwBj5kW8v
c2cLK9TCGQCkFF+pRstb8T1gd9mgPVdsjjZ09X029QDxEH9FiEVTe3/Htoce
Yr2d+MKr3UUsmzNB5Jqt7OAG4SEUmsL0lXEhoWmMRLvgUe4GpvPQsKlK0gPQ
cnVETIIzMZargpQkiM6R102TNUh6Bp4yuOQYOmpElRh8O3RsWVLYqCDuuWvK
DOtkZmuVTB7dmzhBhTdfbIBTi7ZepvTiAvVuiNyr75iHcXpXx71DFA2ZsSm2
rV87o0TvQivEeSQeK6j7E4jn+5AAMrVxZrytVvxJWsSmPHCscqjPYgLG6sQ7
/jt9yGMi3CDnUIy3JFqfolt4e7HEo16LqLLNaGjPlNQ4O6B+7DikGExyNliL
qlw+hmhusABIsDtU+dM4vYlg+vUIQgjZwaXK19kd5tZ4M89pw8OfyXH/Zrk8
Zdg52CyOtHdJ4hlNtZ6U4ul5I8Th1hhbmK+H2FESSQWgFpdbdt3NTRavoV/r
lyAL7Fx1158S+n08piJtqtP45eDhjCObWMgPSuCv4v/FQawY0iXRaa3597gW
kAqofsN3GalEZkcn5HYt+vUHcBEEU29eoqGZIsqcqa1Zw50Qlv12Dk5X1KH8
cVb/MNrms02yObU298M7gmAQZSWcLhjuRJMJgb3v8/77hmUlvegMqryiXvIR
FPoi9NU5zPQO2wfLKKch84RD0hUDcvflCEJ6MyHzWspqh4FfxeuOohmu5vmx
3tacob7vRZeZAlHb4hiVFjBuIbIHKTH9v8DGi/A4+KOSDBfehPMwtnz8ha01
ZxQuy6XtCtN+OPT9ufzGfDS90gKftSPkbvSRwdH4ko9sK1qY2duLxpTCyuFv
whj1dtjHJWfTfL5Slc113ucNnG6bZVseVtYQZoKe2Z+iST07SBMx6UBbqPmI
X6AuohkmVNwfgl8HS7USMtr/LVVHsRmyrcXixYulB1K9mY0YyLturkKyrs+y
vxoKeEBTxZXRYZgZ/nfgwT3syOFyhzik4t0vYr5Gzqa71zwi6RvkZAO6YkfI
2+gNz6Cf/jVWVtpEGQErQWEaLq0CtbmJQKzaERZvUTcs56HUOBbmBW/dRtRK
VKWZUnsIQie6c8Z0nptjVTHeKz4/il4LjjS5Axel75j3hyCoDZY/7BYhmRi7
k9qa7Xs9QhwM2Qsgrcv08ZPTLu63Ce2v/EblTbHMq6+sPvVFSzD5DYPkfJQc
fm1mY45GN8VRRog9TJ7KDPYIN0lp9agB7fpFORoAhw4WcB0U3jqVK9H9iHoB
1YLEUInt5fiQBRA1w+aUOL1VaPmWUS/8GJ/07d9KitK1cyGcSU9jRXQdd6oH
BwiLxqhoC/gZ1KRUbnxOInWZmKm1g40ZYGCqmbu+89a76qn5kITGts9S5wDr
K/Zvkv+Wb22AIE+90yT3zLNaeiqthmUBml2Xs9GzPe0Ijk0IJkIkPCiaX4/v
F2cjUnrz4GTYa1K7R6mSRkqJuO5frgWWPdxLVLwDzizAUpM2wSA/Z4+tTLJ/
VWzIqWVMph7qyEACQCl5dURtNG9pq96DIxyt7N3gNq+zIt+QCkLyeDPFqyO9
sWs+kIo9+Nx3r8BSuEac7qpLLuEOEQEPlQRgSRa1uI0LHf0jiaj+VdCPdWik
dEfs0Beyl48f1XVS3iXCZl6pmedWpnw6u/rqI5QhuI8sr5TvpstRoFzkAELl
iVLnTVSJs02qOaE2YYdVIrL4QThcy3VlJuYfPtJGsHllwRltmEzdDFGey/Km
tpz2tRAu3eCFLD4ZZBN/Za61kG+UpAWiwHUk0cck2BSsiHnRbZ2GLYkfHLzE
GaY8wPKd9eq2XdIdPfHkOR80CmQmdBJYqQlzcfvZ2xZDtX127KfboIkuHlR0
1YKZFBnVuMLifeH7bSEXIZZJ1Gi6W3y1QbTX7Zch8B/qq4gjqbkNKtcC17Cw
dGB3diMJb9GS6BOGOUQ5I9fB7cyJaVc7XFWQR1Xg2wPgtgi4lAiG9eIfDZuz
ROsRCW+5Nl+niX02cfNJMDCO3PBV39BtC2rH9uihSD89CSUNqzSrTL2etVvS
yOoFuJD6rDalLEdLX66CRpIanUN1JuLrDGwAVG6dWehYYrxMxcjZ7cWcie+I
Km5wam2HxYDHyd4bU5mfn8hSkCQ90tgrUgIN/3FSHjI8TWl+yLFqn1zelQok
JPohj6ZsjgbJNsY/8O7JLeClPJPJoguTHyXbep8QAfNDaxQ1thHwZtvuI8qu
1Z7gQ1aV9J/i8YFmNTw/Hfo5AXVKjS0WGRRRP0l6Qm39HxIDX/J9MSy1Nwf/
gHKBfxhSrjjB6RbKgHCdrVO5IjbfYYmHFnfsPBqZlxtMnG4t6vKjIHwzN08Q
pOXEy7g2dl1aemvcC+OdQReXEt9jpdGC9vvowK1qJ0lsLTl20RWsGjUIxC5Q
cOZDYPYZpBa9izgvtfA7hb3xaiBu1jilftELp0S3GPzoAm7TiiNImbfdBags
bOr2pbbzI799/Ce49o/DxKxFo+t7eUyZwApKP7mY5AMEvEbIMo2TE4imTzyA
ML/kgFm+tSDWpmflw/GKZ76aF1PKtl1qP0eIW80sKrgzdRnlgQ3WNr7DT4ip
ncA4o5ybOM3SFCND6OG7MKhafjAKPqytsMtzk0jRyc7gO7aYnErbsAFP6R6r
IGYX2cbXH2SlNT5NbD8MY0jJQd8m6MX4pU3gawsE1uivOwpvNhY6NbwlOTPJ
ieQ/uGC2JNiROAn4dx/wC1xX5oy3aZf7xi/IsEDyZPmbcJNRf0CRS10fOsQ2
4NREE7WSM+43zdPBN+tgSqMsGqaR1LUgY7CkQMU//+AnRTJPOsgv+6Cb/Upd
pXDbmI56zAGV11I+snOniK6WjkY00Kl+0M4QTds9Z3sNa1U6Giq+qyR/aCoI
vsCs26GhHRVn2Ocfcf/kGDYweUHdcrTs+K2nLJ2zMzB6H3HbnuuEcjfEheaS
mnrck1vYIcZOCjoX+ZMMttHTpE46B33zAzMXLLuCQ8siPi1juwGf7vohf3Ra
3Yjk12Z9n1tWuBAK4m6E4Ui8zMRk4+s2zLLItYQJpixvU9rUQJ8yUM02RswZ
UzA5XS3tizghy0mt4i/2xJYA2wAmQvvkwAWSULD0hGhgnK5ivPXURqX5D3cm
76e3vMFcmSPdfS9r3AJiqgOrDF0m7FYE57ewVANZe5HDy7DxCsEOLYDZnv3R
AjuV5bwZuwW2amLyhqRCbjuFdAbrg7WPq1imOQ2E9PsFl8xb1L/eKAaBbxHO
mzL12/SAmZsBxoBY8Lc5BLjA8Wsk2ZN6MI3KRIE64V1LoyN6pg1ZKZjJ6I2T
MmKzLV8WJtrWagGLIVTq7s33+3Mh6R4IZQpWacNvY5QBhLEJMYLhWkBgROjJ
E21RFmdO/3+Lbaq4yKDA0ZIfhG+1rbrjFTnRxeq5hGn8cpfJCDpOLguTBkyq
hOQje2Iwu0qAcfue4glRC/2DW9hy0+rRl24Sz9M1v+AjR5e80vo/Tzlt2ZVs
4MEmEumM9MvaDLYWT8TYXG17MdBDVZ71vysEcgGNEwhHQVl3vavKuX2vTxWp
QCR59eiaANjX0fVsLXzlLOJkjk+3GSYD6t5B0LPmfsoBbqi+B7HuWeNJjX8/
Vs9cKL9Dh3R1OHHvaIAq5IGgOX3BbaI5NJCc3FhVOWFWfbQQ+433fHtDxWxz
EOZKQtGuIXy9+TB/r43/yrc+FdDgNll7JmhGSmaR3KplZLTr/evYCKdHTY5t
cxvpkcBToei/b1Xy0V5sW9qmrNwaWykPXgh9MJ4Ny7Az72EQBFZX4hAV8+AN
/TPGbggT0Chhzd9PM41bXeXVcxLLq4W0ii5X+KOu+eK0VM1ltzZjP+Jg2ZYC
a8YGduRzvXYyoIgdnHxzGUoUTW9VttIckDLEFVO5Y1VvnSuPizhlEe93U424
wGvRfhprzng88A89mlN/rvvyo8UMo1MEMGnx195DToRvW4+qRKb/f6QEIPgK
2c0aF1BiRj/qLm6l458dlIfmyrKGYuShgwyc/PUptwzOw1Rj36p+XRccZNNl
uwMwXLUsUkNVnEn4jj4i3jztcZo324FAEUoAAK5hJjRcTjAP3i9vGOQAVmWO
+hFY8OWIaCiss6+8CRH5JHrAtJG8kqcelQ3fS+DGxJrtib3qeWrPfkmK0oNv
HzMz2FOr3skClPRxO48R/3CIocvSKi6ROTQC4Srlg8w9tf6S4JFKCF34m8Cp
nlrD42FHyivmzTievgk4AUjaSxloHta4nWVfW2mK/qWyKTSbct/BhhbIl2Hk
VkePr8J3FSiZfwVvCfx+DN8uP0hXdq/LPObFJhA2KAGB+ff/hHG1UhXTfS0H
Q0EJnEmYZUP/u+hqIzov8mlsSsi4RxaltEIr3468iApMpr0fxGEWL5b6AAou
GARbbT6NzRuHfSr4bnGuoLfFr4YsCcUVJ0nOw7IskKeSwQL1LaUWXcCLNpeE
x1Fm+cVETvqDanoVhXdrX5zsFjJLyvByagsbIKhmXeKbvG2oLbrJaMgKEgpb
z5sRF3rxLwS78FcBGyjVjBfJwOVt3GV+zUD8qG5YHdaYu4DR2BUTitKAqGNP
SRjvK4OLJHPP9Nr94Xj7aVF61t6iPJh8AN/EihjjSG9w34iIEKgouSf+3Jz5
spiJCOfEdiVCXE9FT+be/jah+sDRINgVmDFU13BVbi80XCTvZ7i6rjh6aJs0
w4nQTKos1KNSwGbTiMAjkUTlNCiYgzBqG89D9s3eiL9OPk0OjQDzVuE2SONQ
XvrP4DNSoOE++SOpzWaajooXrlF0YD3Bt3qXzs/YY2XM2kXS1fmObR18lhpA
DAIlcJwrXF18xu+SfzXHjpUKJJzgvnKgDyXYE/CwfTRrUZ+sDc1PT+k52c8V
K0O3G41T6axWwz/xwSTC89mwJg4jFh85W/W6RIyA65wzKp5MJXwCsbLCW02t
N0lBo+QYLAmZ5otFSy0nhs4meINu7t4MbsVsRf4kbMe4qoWNAzLFH+e2ifST
h/lyhAbjQ4dt28Iwcu2w8/iMRKcZ/dyZ7ukpqdA+xsT/x3o6cvtPQ3DMoNb0
cYsIAkqzFhV94NkFTQJ726uRS/4jMPLZIZdy+bvgTsfdFjnfColLMPEoYgCD
sbfX3ybl6Nfn+/hoOJErgUO0vjKebYJIJyGoK4rF2Mc/RtCDAAL6KXGJQE5T
GteqWSJWuMtB4vQiGH/soqMKx+e9pqaXRiWVvR+4J3TV/NHFpbtiavUakjqN
MgbIjJhmfvdqOKlbPTut/OuvAW/3eBIuNQ03N1Cf1/wuYj18M6PzkLJvBGEe
cW2LBDrZIsVp0seIH0+JjHMx/u2zvJ17yriUorNyNPLqQQbG5+L8GMWFUU9w
7dcfhRkj+VCbTxmPVCK/nwHvVDJsJw/COE4UWHk0UVZgGP87UNAIlSukQ4IZ
S++8Mm1CIza4GFyBAW5UQCS54rux4SK1yK5kl1Zze3RTsYnGJ1WMOEGfP4ca
Q8Y+QAXHWOuRUDe/QcOvgTk8HiDmAyScxotAGMRF6WCruH6Z98JVDuZjKwCl
iDQJRws4e98bcfVoHajfHQ4O7t64QTA8y6N3UMiUAycAI/BCeWKFEGa+30G4
sU/YiAUD59JM02EHAklmfgv2vVuPZZ11JBfUYdAB5oRioNKdO2mfKC6TXAaM
VXXlHDCNLUrdIOKG3hsK1JUYXevRrs13T2tK5Dm4JOTlfg7ZxMMmMiBBvzFn
LNPagk1Tm+aIDCY5X+sJPO9Is/bU+LhMgTZYgJi/qRV9X8NWmIgeq44G2vx6
UPQJQlzBAOytrNR3591BVu/VV9oAMcrOsA2zPe4ftBpbx8xNIj8yzTeu0mwz
vccdv5VgYPJYr/iUetfxQrKrFRxtjhSqgx1uHAjrrHcv06skMsuTyEomMyOw
xhx3JWubPRxRA5/ZNdb413vYw58b+ctit7832V1xluEKw9MUeaM9sRvRgCfb
47a+VUUciQjzJvdlVovzJ+5jYWpzh5a0gvvejVj+3CxMgjpHT94JLo5it1JV
GYU1XGHtLcZ2MJLBbjY7ExuNxmNsm3ZmPqDF3Xdyf8284wfPQlRaomFoP2ox
8bgbdaeJuKXX8oZ66snsO3gbxEBjCsp3pV/kvyHAAhRMzzaZ9xs/Iw8icSWm
H+epYWFZqoeTdCNYCDMljBvD8qjuKrQ/rRMMMAplZXKI8SUfeSo/4earD+/T
DlkbewmaxcSM0har5rgdKi0KAFcwggaJubVFG+DJdytlLuSisD+SUE02RPsf
R00+SbB3jD1rQ2aRscejWdBk3saERPvXgoYlGyyMVEdxtrt63KzY5FqSnu16
XbJnKO8ZTUBbjHoFCrjVcE+RH/PGjCtQ+Nsi5T3wZL/w5yBdKFbUZTNZxNo0
TbR+fClJYcgHoCBC6T5FnObhGpfGZuWhb2oRtFnasIOisUiV/OSstBzvu3Jf
Y7FF4RneuBBRv5DUAF4EWUpSAlQ7+gGYbScbMiLaSvrYTE6tKwZo4jQtaALu
L/f8eKrSjva84PHvWfZ2uS2BC8hGJ1UNxxl5z4TtgTiBqwSG0sk70T5IY0rq
DFgjsBdWhVWvR0g7qecTNO3IISqHJ3VwOQHvRR3X67vPCaMRC/F9+2wHKAri
mRtoDTaWgv18BggPPYz+SfEss6PP8L+8kZeOsoivoGKzdcEERa6xQ/vLUImI
j76D/Uaz7JMzRi2c1DY9qml10kBrdmaHSacV6vISRw8/dis8riJ3UvhE8BEL
pqvezqDVsXPDu1oAYjJri7ME1kSnEiAfvyRMZC1D0KGitotA8sGXp+Fl3Kzs
AgpPDBb4dtUGsm1Q+TPi1LdEKb55o25vuK90+onCHs8+MxTh67FhHzjJATVh
0VRdSmXBPN3gRzsdW3fYzDQYhcdVH4Mz+bH4DYEAtXLew/6pOL03+c+XRuen
pJhhI3q2uLliawYYZFqnmzcLgL3xH1pnZqlexlQGwJ87TBYZq3qmUPLQa15N
yh/gWQber8jrX1lRn2BqOcgmaFOeZvQ84fBnulVLn12NnlAaRMKKfQp5PhDw
7xz8qbom8oXUyowD3N9P9OL8FjxM01f/zkLSjt1FRyebZFbB0VQ+sV6eejkr
eEjeb5p6py47U5RAsAuCW6O7U9B+pMxNRGfzBb0oqJXT+7n3kMGJCYTZHcom
BiXc6aoPW1MN7kOBQKRA4SdqqXrL2Cg8y99rp9lsMlfIZv2dRcBFPi2hvspJ
2GsMZOZikWLKWcPnt6HOmR1d1P2YIjXiPXY8o6tnjyFxCarChezEbvOjIYXi
6oadBQZjpycH6rMcBBCcNLZFEbad0C0E3ibhx+hDJ0qMyDh6s//yRHo+9dJZ
HO1wkDAUbcrQY+zlI80cKRNOOO3BNVPfQ4y1YNGN7EnswJfTyNRiTdNm58Cf
NzXIfhKrEq2TECc1v5ipZOztsMYey29pr+/0dJENUoznfJBHHtQabQXXjxzz
sAvadVhTSKTTtKBssNhCREk7d349kaZNi9ope/h0RouSTkRm3jSc3U2QYp4R
GX8KMN9OiW8VoH6setbXkQ7wAVNayOl0gsNRdmTyBcQ+v1U5Vzhlz4xdUVdn
YsW2PtnGjj2BJoFtJ+KQbeSOgpy9BpF1rQ3W16cqQQdJ6fgoe266FGlxHNN/
W9WPRsdNg8DeQ0eZqeN2IqZQbPoz8SC3r3zfzFprIZ1FLo21Rl9OejZziDUM
3dvW5Qj+JTbUiKwdgUXDCNjmnfZsqAsrumYQSzMdHBsdFAIKAhdLPF3laqg6
bWLzFd5sk4pMXYVdm4mOIizR03Kc1OkJ4eS0i+oSIXQDoqy3cL8OlOTMXuax
h77wvnYFYqH5GerWhqyFxCmIbSQm0cjHR57Nil9v0HlBJu9JXevhS81Hxu5S
EGlp/HYnQ5Z5zg1Pzj7E/AkGOCsnMpJrXMY8p4x2n0y5DfGy+8IGa4muUdj3
PqPWk2+ICWFLD45PcwXmYQu4D22cf9j/miLpr/Vp1Sb3IjXIeUoG+xsppRaJ
5QE4O9bFf8By5Ywv6dUI03xVYrSwxSlBici235nCg9UF9epv2WZ4p5jUHFMJ
oYnnt1T7Vx1tr4U04L0doauN54AHblQ/E0VILOa1pXINcCwsqcvwZ69/dBsg
AsaC9SDa5iDv7s7hYXetipYtVL1G5C89eNjZB8OF8dBqE3XNchZDqOSMdcDt
JhhNFcbCLa8F78gJWH5Umqj4hqsUtw7/mes7imKv4joklSRZWC9iuWADeqCR
urp5VoRR9S0SluxgeRevJvR2ig55UFD4qxHgGP+AAkYELssc/V4n7M2UBB/g
R4EIVBAyG7q+lTc/QDUfqS5SSTUH+FCbtGt405yV54DSiWGmHvblbiWt3W1m
LlqPPWNkJC0UXAQ9Lk5zqx5P5O+bxFtY/7YbDtQzvNO/H1YyeGlE2mFTTSly
2oCgK592vcgzNYuHRP5mDmcewJP6Fq9esJOaV/gXaqvuYI0V4J8ejxhY6avj
kd6oI+RGcVgjW/Gxt2QuYjB4gJefv5mWI1veHI+M0RSeAfDyChb3ubpTZOtO
dz6X4TVp4cE0zmdtjjwRPlbnFv1I/epy9aSfNQQQkstK4PO229TJQMCKMYzp
mT+FvpEpxqgjYVQBUsu6GSOHpaMtBIb5NZ8tI1uneAIiv2umQpTU+lDnhXW7
Cw4BE/iyo/qxb8pXlvgSMB/EnhleSE9Hz64TQw6k91pUSoinUzjY2X/NIhHV
tgJDLvxAHn5FH6yHz1vUmZLar3gZDaOEmWguoCV+vUxhohHQdipTRziLW43s
EQ1B3Cu8ePL3R5zOBb1EzeXZFL8nqix7d+uITM8Q8Bwx3NKthZWvJjvi5uCQ
6ROGugYo02EGSV7Zhpgfau+fCQV0VR4PnS0eVu8iaKhy01uK4K3tvvEsoz+2
Ao78Rw6n7Rqoii4spwz3kCQQOqr7ZXlUllSN4pZAx6Bh9T4+fe/v8jncwmML
S3gCuOkzTIVcYkwFBV291/OesVAGiu3J1OUdpYM9/gE1IZ9WdhdJeD7W4dVm
NeGB+vB1G5jhNQwkHObBaQGIFM6Q4u+jhxcvTD0ZK/Hxg1U+Ny9XQWuc+79d
ZBIz46OkpWPiG9UG9MI9ntWksfFEo1RmafRA6ko8pvwE3gZ2A1UKTyJTGK71
UIvYo/9/qz82Uklar3djlKCkqN/a/64qaTfLyi0RAPOBW0M7497AFpf6JLj0
G+dI7nGTjAfynWtzgj6Mi6vHO5CPH501UqEUcuu+hYAJpDyjTliaaBkyF9SE
RiK/pQgfpCKXpoE8Oq6Wp3rHn4W2H6MS0IHdTAz0Ky94zje6CeNn3r8AsAOf
9rAPR0N+ra+CvpMc75PcIjKOESa4HLHb3Zhf1xKIcrB9ty9/jW7Zj9Yac3DA
++OUzZ5Lb2RHoTMM4rzW+UO9g45YGfbktQWxCwzFSWHLfjgqIK9hkbn4KZ9X
jycAMSeyTZDiUU70j1gUL0a6eiH0L13ahNukQfNHZVu+u5l4DkCXVdVazCs/
e5kjo/zQeIcZWJRr7DruXexpz+FO9LvafDCvG0ignPrtuLtnNARrBujIO1Vx
WPiHQVmjeyFBA21UxyDadkQfT/N00lg2qISGSXzuw2OJmM0Ex6RYn8pSF8LW
JZ7VpDbqKA6jhS3ZMPsOzdIjSfxr7hRMpO6jZJchglO/UKUDtfUlXSI1WIi5
ojH+nhiPMIQsxNCUsDa9e78g0RtXrS+/JO0bxAX8SnrQs6a7AO0ayrs2/ezx
FQVyQROc/5bkUn75LiTqbxH65JRBeyVVHuTNKRzUZQwvfDQiPfi1nqpRhqRW
fnEjYk/fWRnm1M41BNsH/0+WXLsTH0bAPRRePBofiTYfLkTzfwmv/TbcFtwi
rTtNPKLrgQFmmd9KNN47tu5asUu/2nSr/aGWpitDWBh732quKlRWFoysLxDZ
zbbzTNXRyeCdCjNSyyMc4JbQ7McpzG06fjya4/2XVHN6TgLc0+ze1Q9PjGMj
INZHzFD3YpceyZ1MO+wPcn0bXDFZ5AfPzqrOJ63MmDxHdnjkU0Fim22cIDbO
C/2HmaYpcSiVrrmniXmTiWUVZcEKhrgvJi5jaf1//Ixgv8WsHuUr1Y2oKJXJ
yLwUjPdb8B5AKL7+Q7nUuvEDdNzPitVlTGZth8CK6GNX/Sm+YhAA+F7ezptT
nbyYyhcGMWew0QiiUhzqHHkYXYW6hGho/fV+XSo3oxLiuhQF4z8vklbgU39z
1DUadleBSzbni/rBMxH8V/BqISZAcrkOLr6F0pfRkOQzC6YWzugrVj0gSHJz
1/8Eiu6aKirDFY2OHf4rqoApc6WcM+wFPMm6NE0VPtvWCwDThNNl8R5ESZgb
yjlEHY0NZXpYY42HyNRdTG39h1wsEM8/N9HdBF52mcyO1lvx0LGsgUKW5Xnt
nymSkxblJqjVUf6KnWlKshsu8NuTCxNvUFBUZzDUaSNExsfea6Dzw9+WqUYb
WOjMg5LZHKc8xuqWWf0FJKBs35id/CzVr9KRSFng6CMUueAHew8GLpNJduNG
5T09R76j/smL5Y++r4qJhsgarHIc3y7O5KMhdct6jF0He6l+Q1GD04HVzYKz
AYtcQ2YMELOI3kagdDZ+9CTwZup4mCyPFG3EO4QwtihU9ry8uDc96i/9o81w
kHcBzTaRXYyogSAHdhNauRlLQJCHsWIdlEWeBAwFca9YWUobPCUVBkyU8UBX
awi/QATGT1ocjR3jrrHSYGwEtf5v0cCnmIvTHMy/qf1wZiIkMPauCPTPGRgf
XnUTAPQNBODSIHREpU3W6b4cutzBbp+F0s3obBssg7JBJClc3xaUNqfXytbh
EZQq6D2CO59y/LIK/g3SDR6sIkJTuol6QxygSY0dfIUGQoecY+HaMlMgDqFn
73rOcNUB4QvL2zUwcCZlzjf5aB9gdAQmV+fUCdtqVz4uRSv8iBkjTSWUUOa1
c7EhnUJybIoqIL/IFJPl7+FznFG5h+qaoi8YaAutN31pk7RVs4ViqjJMEolj
whQYiUMDFUC8phiVTnyln9zfaV5ZuXtmLJB9KLWXfdGpI7jJobCcKegqrBZr
BYKsodi6quO7c4x/qJ9pD+uxYtn6jmexoAMc9qkf5PiODx4H20rbrEBdrUxH
Jo553lTEdL+5axDeaQEZuPtrxt0fm3ti23L6/MF7klG5FKJVWUKGJ4PLIvYf
9vhcWAuW7p9w50M6wm5d1tqHpLqm9iG4HOGrV0d8atEB70t8Ut6jVpuznJ7l
oNu9Kj5LKHzkT+MtmO8BsH4V3JGnjYE7N3ZQQ0ZECylbgkoKfdxuWRhJVIb7
bk/yzoD6IvmcbPruFImuDDmrnNl/hWiGttX7BJl5VFMiQifftFZkQ0k7ECtd
RvHzukiHM4QiYClRS/M0LWeKeWBurXImJpBgKrCLTJqYtUkz4ME1s0Vlx+lL
MqUXvDhnK2Ova+oHMFnMHRynQgEwMQBe7ZPHY+zsC95p//XcN633FhTxAArA
GZT7rRhXKN/Q7sctsCVerlgzxgTsykYIiL7B1EVbdSuo09VjTkcKJjBQ/hi5
O0EkirIz8wV5E3juMzBI7MNRBDrCqonKKjI5m8hBG1RaIXccZXD1eIiLfAFP
pHICTqkIKZpSd44ndeJeKW4mS80Q7C3YOGPyyEU+Tn3IH9JTXtR5esEdsqgQ
UllXXrmZAx2J+bk17MXaYiACE3sTfg8O/+hcFpxDkSjCYiS4yKnkGruHW11b
dyeC2RHErIrDnHEg1eEjJyvMTYKnMmA+QzK1M9kQwjgM7B/tkhZe1cO6PaGt
T1TxjJ+X2anB1A/zmz6Nf2hiXgM0AQzS48OcgGthqvvcB52oSN+F2Gb4SzFc
Tf6OauZEpEJP8mSwpMOPEfanYIG2Vl8Ud9AcKkiTGQrbFLUfhaYnPkIy6uyc
Q4fjhfWlw0ApiIGVQxql7dpm2Egj+7bPCWzkPw5/CWqAhSC1PxftK/+cYvQw
4vU1mNA5m/vGaqPucIVtvAaG9Fn/OozyOsb08N+h75rQy9JLkfR6/uWdtKIr
j0s9V5wAQ7XQomXaelRYYjsgQOdttbvugB5gFC6p75HfaIyRMtnBVUz5FIiR
oXspOKhcNKL0bKsrCFFtLf57vB16pI/p83VXOfNGonhTlbGip8Bu9EvlReYT
xj0czrs9SzztIiAugnPRdFSKT2dr1sZRDgIGna0ZDutgdmynRvLuIDCclODy
l4/4i5NPkFL1N01pM1Uzr4CePJOEWoNyzOPtpGDCRj+66OGIwq9W4r0QaaYZ
Wj+tiF8mLYPfA631HNKjielkYgBwaFEuwBCVKpnZOlL4ErG1jDDkyOMvHhLc
YV2pfd5kvltY6QmbMpFPhUKWV5bDbtL615Rwm70DG+rxZkFbrgWit0WMjbzV
l816/TKTsj+7zYAmK2Kv2i3cLz5+UK2kCHSAoO2UAWGMkmF4qiIMFSohM7u9
o2Bb9eonjQqtlNtP933/Km8uY5GK4CGR3IvO2dmXnnlQPoqm+Cjdy/FfQWRl
B7ZU59jEwetS3vHS8mHnZ/aPckrffUhBhigu/GSMt0h3oyrl+QXDAVJv29gm
vSWpfn6ZBFs2wB8fbLOovDcxffBWcfM+QgLUXM/MXPeoXjXDMcxNaBYb1Abz
uik61QNhhDZ11wbaC0gWXcFqozAvHGk7mcttSgwUKfceMHpmgql8UMsdhiVv
IfwfxlpW/zHqaBHbz35lQDEKEv5er1sVHvk73fBOk0s/TsUfh2dJ0FMm7+q6
hhZaPQ+JWJd72EX4APxSi+z0pvMQWtOFyhSwqpngL2hG7t6NA/8EICbSJ8Mj
r8MGmVhkhY4VXpLQdYKIg/XVF70Q77IclpCUelHpKBZWjLpTNZPCOCU/sXKf
42hUmkLE4OXiVqdEn+goAe5oZC6MwJFv6IkRL7xcpbhFK3+ia+e67LSaENCW
ch+o/cm0Q3ZBupu8RuGmNzDTwz1V4UkB0WVqSRFi2x3El9zOYiagQL6xNttx
hHZE9emJ2u9TsSHEeU2nywJ0Vn7urZq595LwHYRCTNf18+GnWwrQScyRJx4x
ImaJPzh99Tg8P03PnBxO/+WST+XL1nasStVp03sIiGevQwTpkQopm/hVy2yf
3DLKmeZQN8tGVzKBsOV9fP8POJWv4uCWIZ10j10yzsLyHLsVfJjpDnTfgqy9
NlM1eiB6LOG3ZurbB+7YnNfWkNySKg9YIZD5MIcft6Kmu1+qm93BormpDeRA
DvTe/Q6okNTAhrcspXpW4PwSRD3SA6l0nlrlpkIibgHJRyGDVb99iwRjRttX
bZx0svh9+YfYM9GEeV1r2LDb8e5orlmhho5H+ZLAYBI3fqGwseqcI02ELXs9
HDymyiBoiltMx21WhMK0dOHuWty6bvulDlXDD3rMuZiRY37SrfZFPRjLhHf/
YNqKbf+uqwYulGEYGBw4O9Vfd4FuY7q8qq/XHWiWOpKKyhS8ac9gtC5+hwd3
4mZv1TWU5CHzk9kJcECSi1OxPvZKKjrTL3yPt9x74ViX43uXEMoyZB3iMu/d
CSLcvTo6t1IJOGTu/GjXg5ReDUIUFz2z2nk0lx5/W35pMmX6N/blXi/lZUGN
e+hKcNBcyU5Co7QizBU6/V5mhIfbAJbEFgfg3k8id5YFLqNntRRSyzvEf0jy
Qjr7wNpgO2KHeZMZkuCvYXiwhOCPqJlXQQ7/5WtIUJcFi1YAIE9GUFG4n5kH
7mVMKAWhs8nDa8gly4i/rUTxq5bTWYqoLjOCEq3refGd56O/a3wNa0LBUTYh
ivTDPPEAcvRJgXGclzlNy3JWSEipjHcGPIBEQoWYS8A2PFWzmkzJGroWplaZ
w10niHbZb6wppbeTKvgIZGavBcEGSZy/tD5P7A6HUbBCSctBL5A9vu9xqttp
pzYaFczkY4MzNigsi7+lh1yDRqJA2l4CHfGgMS6hIMMojZXPq3fs4wMYDwTJ
VIGx0X8DITcwPO2GHEdr26ajdGWyMQx4RP5zWeC0yfgliGJNWL02ztrz3F03
pYPkZSJjdw6XpORl2KzXw/p+40dSrCENuU7Dpvlfa9QRGbf6lNWenjB6Kywk
hy7iUV1dn/Welj5KUagvzSanYryYFHr6DCDkjfPDX01IGpM0ipL4Pn7LxMJd
oYbukdw+qojBhfO2rBkYFrto11YBqo8i+0L3kuRCt+lxtbgXKWSylqyPF/st
jGrbxBzr73FGpylNI43SKAPIFP9ZIqto63dU7cnsitYT11hHi/etUBwS2nzp
EFYl0gD+lt6aMBa99E72eavCHPIa9qrNfHp4aQLjZlmSMb4VbrPMAKKAvI9b
jfQR10cQWIjfufUMDau6T5WkWWAz9PwSq6H848+kBNmMfeEJOxY++lSntwyy
/zDh4kc9TZZQ4jX9EfYyLUFwyk6kAfkNqniwNJL19ruLMUVPDyek6SmLfW9i
KlGh5r5dYlIyFYThGiqGIp8Rg49lkp0AHq/CpnIV0yy04ebHgkOOT1RqAnok
Y7zOsKFLNWLqq9O3hrkPiuS9O7PdZ1O360P1L/1V+vyuJ1dnwjUeC+Ti+bGU
wB0h1uMx+RPtIWrEFrhQwITYLNyws3CK7WKJvc/6v5SwJxcHDvsff/HWFN6Q
+xkG83YdLYs+e0CHVS0UThaD9Rnwh1qQo9v4AH6jSSMrGWP5xsBnHACF3uHc
kNgnF+S9QjpHQnCrM/pqRgo2G+g+aBb0XpLzoT6gH1Kr32wEnVOSriEMioqP
19XnaQL8GfbRvNyigooUmBmQ0Y68NkLdfcoeOAmCe8cqrkfAHiKaWX0m1MAG
bHdhAEJqXZwkID3wefNpciL68FIa8tvOx8AeFKloDgDnadUdDiiTtE/d6NC7
fxbbQoYDnJ8aj008EIeWp59aNmA93WRfypXyhohniQ+9w+QTNtkKdpB75Zk+
aPsVqW8cD4gzlqC1YgBYhbw6FscMkgVOVzHifYvYsqmG+Q2kKtUlizpvns2I
AEQOvEQGLdg44HdujIDMdcG8d2LL5/VnLuakIC+shr6P7nP9GaUAZ1hHWugV
blYvBuqCpY80C2hahPeut78SodL1HEmDx1oh9zRC2gpf4+pzgewIC93AEW2D
IUo0ORDo4IyPRNsl1FTBvhjIYqucExwV0weCFbart1yBocYTA57wDDQaVI+a
fbvVvFLN+FJ5Re/8wh64/wL8n/6TbCghmMRGB6xInp94tpdIitgscAGzHuIv
IaXa0i93GGMQSIMihA1Im7WDMfkJqvcRd4Kkey25drwBr7pbIGRL0W/D3FbL
LWzDdsVHaVAawBhXt0He8diNr9HKozB+1BuDOQYAmcItNKIOLHCzmkyzixmy
dYET1mhal4jZtZ6ZhGollZovQNxh+6x0SLt5wFQlUg9bvWNCM/tJxL0qTaVe
Z4T4jFMUY0qNDW5q4oCHYeoEEATp2FPr4nl2jv5yALp+8Q6bZnHo5xJictK1
x8AylYzOG15NWhWwHjCN8mlJd1ofMRjJxOJgawWzkIxy48NOLZBRjUQv+r27
2c8h5OuKW805TnHih1C22fP+CiyDHZNk72YKLHSk3TaRvZkeprGMaK4fmGCY
J0FvTMmX2J98CQgtBU67E3X3GUp21Q/rVNxL/uOjxHhu2lC6uQLbPr7y40/C
fu0wnPtlXENyFdtXt2me0J1hNIZ0cCKaFVP3VMfdvOGUozHasgcn8Zg1sWl0
zboR9l74CiZJ5p+zs1NOT2ONHb4Aq2c7BAfGIkw7ugArTFiUits+uE6q1h3h
d7l3fGXI+Mz0YX19xk4OA/AsGx6MTg2D+PHM/ezcIdXFGK8PFk7uhb3Y5V9f
iQc5QbgBlekSZ8hbl2YOYtbUXDNnsvRhY2LQaJBG+ius/wWB9F/riJseNp03
6ZeazqulSQRix1jpngRL6rEO3aAYx/alBu8dy61dAVv424TFtaYQIpNAhmcG
LaWB2gK2jP+A2Q1lHm0CxTMGDXJy1N+X0YK7tLV4c5ih8cz4ygzxN2mzc4VP
NL/4l19FRkDQ9aI1SRMcVEGlj9vIcQeD72jNuWibK+VOksyxFSHGGRkHSJ4N
EmfbALegal/vLwmsiQDO9fob4H/N9KUFwVy3Sr9j4M/GoVG/MY6tKWJeysMy
5JIn/Uju0L5syOufzmUh/a1h55swQ33DBfYgYOUCf1pb+7ypMOW8ddOPAb7v
jWLqxO63RymIwa9AE7VRxOlAJMTELlIzH/3mw/8VyZ6GeSUfLwF+o8mqaMkj
olfXBi6+PkX6Mn6r51gBYQcFIiwe3su/iyJtzSEvHk0mQnXSRwPF5fn4+fpG
kRwHS8uQcHra2mlOG4cBFE4fbeWVocxPPQn17frhMWRi3L0a+q3VmQor2lAp
0zU9vPyI0C4xqPRIqVwLYAXrNuk5wCUI9rY4MQBhBwy9sSgKbleJJoetDCcM
6J5jn9aRoTstqVbQdWHwEZl1O6E2F0hY7FSomz+LxY1RxKpa03jpN+vdCuIX
Xtr3jrxRYIx+mKquKyc3FRRaguhvXTYrb0aHlAPKLIgltcZqACTaWyIuNSq6
o57Jk9UeFDo33/8mHNXBh/5MfJovLMYG0QzTLKPsHCOZX3sfwQosXckbekOg
j3eHyVJSlL76e5bzN+L56tHL0I5aCwcdX8r4Kuqa6N3Rrx3vdSHma3y2i30b
f1Rb22Do/UDRF/pShG5tyhi2jlALz/ImtEJePb0Bj1OutaXGyyyDpoEjkEzC
ct582HdznnD+ragQ5tyrbrVaOWz9HNWS8Pl0r/Ob3ojD3RTMJfoyscWq1yvf
CqI22EMAclINuueWH2B0FT8kkgQgnsEKJbmyFbeNsU7tUOO/RvgTBOVq6/FH
eUtEwzXapkLWbLn90gfHWG76OWODrrqy12sqYy4Wz9LE/dEq+8qAPSWLBFDZ
Na7BL9CY88Cs4XWpadruVfpJIxXwPlOrG85V9xfN6uHY2SWX8IFyN6g1Y1yk
RfFHEk3ITrgFX+j7PDzfu6gKursO4KqDzpcROLWQSGoeqIRd+jMTD0GKpbag
poaqzibX19c3mzpmBH8WnKwpH8zhmHWgSfNZx1vF5rJaBW8a6gzXIPA8znc0
jDLwZLQHaat2RYUgemcBKr/6afERHYN88SIBeIzfhmOPajy1wRrYBweS+rHr
Sn6bTjPY6WrMKk7+79S9zVN1Z2Nw+mqPdwQ5W0lyJ7c4EEyEXed93k4BZTdf
dRd3X2jJvxS7/S64Nyy1gSEOJpguSAL+NQzjZZUHA3cOee9jHLlO14+Wy8o5
/i6k0RHljWS2bRLhtE4A+1iXfsItnXyrZiu4geEFdsnFv1UnCKvtRT0t6V8V
O+9pGNy9WJY7iZuX78m1G4K5oUwRK2iuIVh/IKoNMkYxnMHRuLPFnCALX4yJ
DSWnHswme19ILWdRhrkDp4w8LP4WHD+KP750h9DU0BfAhxpL52yAfuZsPZby
8at9NHBA8I2yqmh4iBTqqEkzZ1w6gHuEyNjBqwrXQFPhg0V5w2PKeQzMqoHz
QxOEyqet/7Lc9Spg/H6AXFlVnS/kyFWJS7IR3DFSObCnf4b0xDKZyjHfzZ8D
xeTW1Rklk6jsx9rc1v4UHLhS6AykA/SayXWvnspSehH5OvdyIopu2GW0qjZS
zo/l0AqCS0j8DBqCknrYwzDQInH4vBb6Zv08MlYA7jnwR3lO+KUh5ZRoBsUb
JryDOjFN/REhML1hyfoKcNM4FNWOXCiTjgtNJCl7vycT93e7cOq39OIXDx43
24TtfrduF9RCyYybsTzje0X/dvbtVpZRj+awmoUv4AxxY0awYg1tERt28nDY
nPpblK6JNYcZbZ7Q9iihmcUUmkLsqzTXFrWG4kcTxnzxiqy65aedahX+YwyE
fWwZJM/7pemS35tI0d/cw+sD5m4g2FyLZ44lqR9vi41277RwOJfJFovb1eCu
0JhEowqmG27eIO5sXA+O+pb36BVeMs1AaNbMmkxtVCBXnz8sKqozIL6zvyrO
d9Y1kAcnqycwjOp4z6saXijgJUnWxleTATzJoJ89hFEDX6Q3RSfdw8V/0f30
Q34aD0pGPMaIJBlIdFXhLVpfXJmwKP8RD0wjMAIWgg1GEXmufdrxGXbICS5c
Vz7t16reCTwpxlsZqcg+bXIo1rKBuBKf1Ferflit/BDsyWhHdfQ+9GBHgEBF
fx26u6G01X4tku70hfwSMpfko1VKi2qZ6p8VLzzk8yGD9oUsvNxk2lzNHRce
yaaocaxAf3E6sV1UKTm+0lti6ad4dZNUeiQ0sbCclxYjWr53gSvnzNXdUUS7
/S0gv6Xc2vHcbEjqXPvk6u6AiVgb7V3bpDlR4ILJbdq0RkKymf0QwRJyywhf
wKzUDleh9xACLsfCaBkZd8R26bkD+mU9d8rFmWF497DmhMtBxMUmvvWHNvij
R/GvB4B1MNOrZyCW7cTNPEjWWDR3ckPj6jcI3ebv+fooVSxfZUAAIeH8eHmJ
7z097pCBNz/mO9s1hY8Ji+JEpf4/FdyemFd1gsbupXD+8+O+HGiKIOLt1tv9
EU5mCmKlG+LltHisegpGbayVK+GX6HsFawQLtv/O/eJWmFExoChmpmqji4HZ
BRjKvf/qx8h9HoySAqq6Gzc7BUUDjHqmh767bUAksfF+lyaO9+PVLikEvAMB
79zRL+qER4vzpH+BMK8WoLabqcGNvV5DwG4AjRSrJ9NZcXTYCDr2mVkawKjo
DGe1nzfEhoHPL0MOGiaG5K0oceQHijliwxYBz9m0CxV/zLCq7Ns0fglwj7Xi
h25L84fYXX5vWoo2+xAUfu64lhhk+GY+E9tLuFIcol/0EVD0aiPJ/ut87duW
aGD4sWv+Mjpw9Chd5fJEUyatB/MtTw6M86NBlFcel339y4XJ7beczOJypbuf
ZBvJfKC74hVBgqUyjG4qUNJVAwPHUbliNNebcc7ly0RsFWheHGX1+wZA/NbS
skz61yhAzQF1Q+Xhza1WrkAja1PK/RNwlWJOjGXZLFO10VK9C5n62jzeaGJX
NK/xUc9/hv4T7flVMp8UTIfqkj3ju46c4/z0k0f2gjB0vJbAdcVo7Khf5EXu
oAylf5ZvmL1AuxXSU4O0/8AE9/dkpv3e6HITEO8KIRzL+1e8Vx9LwBO2ue3V
lmfDuWtyJOA3IN8VQW/MByRmg1SelHH1VgxwP7PvJtyvCeAd7tRi/GX1EiX6
0VE76WMdXTeT6XFbfVRjFyxRIxDjKg0Mg/PdS4khi3/XrjiWAnFkXGvNHVjU
ixN7ej36hdjnA0cDa5MfLVxWgw9y+qMWiYtP0yo18ZEVMPpPE1nb2kRTBDe0
ttTRjkbZYhn7t01jp3kZ0Bl/s2BmYgXxS9nn+vHwzIKi4be2IbiG/+ntQw9t
iJ/6R3akPiQnjTfppi5FWe0tHYopCq5ytSsaAqHUPTgi/XJehXfN3epUBW0K
0FOG+r5H1SoZr4VAQD9fglGnF+Vbz8Xw0Qv4DBtvUWMxe3lCLXsRYRZlTeUy
wzIxqzD0GOAj5VA7i0B3DNWKf22ArGJ7jbUpaHDYFkcJ1Z8dBJiOgI/d0wSX
P/tZbadPQBkrQNwizE6Ad8w+qN4YxIJbD2snI2zub3okxyt7k8VU4/WWodf7
YbPkrjle81gbo3cyCR10p/75qnvxtIpPpReeaUA489XvHRuBA02SBGBf4bfr
ucpRFJiViDCb+r+n7J41YpfUe2X+A13Fx4s66Pzu8m1yWUtd7TdNGwOKvW/u
lhLTiq06tj7OX3PMF4q2Ogum2cuPlIdqPXgdbIZQkYq3S570aW5Gl1tUhzOf
UsX1YnAmX7EBqTuqtM9BoQmioIMpmp2q6TzM3NK3IUpPM5LLFCZAmIzTWeQU
2YFfBQv5DvFdSgBurskUk1YNgHpOvIRLho2vm165d7a9Dog3AHHCW1QXjDpb
pXLStWHYPLcaEI2WICJ+dSYuh3E57IfEaPD68/m+8n5UI/65j4nVdTZ7tc2p
3HD4PO8p8FogBimjvIRi6Ny+w0W8GDckVfiaECs44I35yu6wmbX7JrbNu9/K
hB8nsDv3+LKMvrK3wCaYo3gKp/jmPFj1cQAAGJcU7/gP2yi2sB6GjVLRcf4J
NSOauq8OFC7aNPlWaMS6dnNqG/GPm+jqjhegNjuEm7ubLdOk/KzXtIgml/Fc
MlefTpxt0aFlyEohmCybX0zdlFm+C6EprCtLc58zZN44JcapfNnFWpJlZkTL
fdnoGcAsVliGuZ+KW747gxNfZhRLz0aE/Gcf1n1xwjtV9gkQaRwy2uK7cIpj
yTNwzQp0t2Zz7NWZAbEPAcRoWR2HcCxyF0VnxcqCOQ4VXpeCB7jGNxx4rp0j
PqXYu2x8aVeEjvr+XcBMrrvhWh3+kqJakT9q/7lEV8gQ3xxt5a0PmBRX1Wqi
tButuwaicRTYgsAwtFAbdQPyr7P22v1kSrOIaqG3idPC4AsikXEzoZNyMX4p
3ER6veFaEhWcRXzULwcQZwL4LuixFyVdroHQpZQUJUPYtkV72+CCDN95Ywsn
VNfjqMx4YPirquh0aaJNuRzNGDJIfl5SLuJp2jNaqI050pHygfPcApw/RPhV
ftjnPxjB6CBhBK5aGFsaeuXY9AI+ETsxzS1wNeF4nE7Dj4iuHNO09Zc6HCrm
uDUBjKjmvCGwYU6cTjFqV2pY0f8Nd4CF9hm4UVJjMTL5k+q1me2FFd29f0Na
2VIZW2DDmigT6BjYQzgRscG+6JxoMmgjDJ0702y7qnZoQrF6N5H2DAvkY88p
NLp4MPu24jaGWCO4IhtyGpV9xXSXSticDMJ2l1WF7SP1TZGnDGOSNvgMiHs3
gD/XbAKy/KWwewwDQi9UaMldI7+8gys9sQQhb7N7DH7+RJgn0KqZceUufGj8
1pDS/nuh2q0bzNThB7GyoPd8oWhMHJoYJOSKkgDI35qdL6b7a0J8GZ12FeE8
lyFmVsPWhVxHyrK2mt6uJOGzyXyDV35D3mi7cQ0pk0Hioy7UCDOYtQYbuJQT
cNHNcc8UrxTLjhSe8wtZREv/0g//ziy69O13qMBYwLdmKEZlpQOW9iOjfo0y
u0uW67lmhf6FPHqczPT48Zx63blgt6qN7LjzYr860Polz88Y36Vc7ls8jPdM
pORjxs5C3kiS6nd+WUc1KQsVbwvr6Djc3hWN8xMtIPFxsPBzwnYOgn+FfsqT
JTmodbeAy8/eYAsd37EWxIZZVMuhey63CTfMtwXcZdtFNfDdvxclISr//X+7
yHBt8Ej6g3eX6lggqwGmj1IEkMEwkwXi4trYKbE0zLA4hBRP5oMRW3uC55jQ
AG+nthRuN6+V7I6l69wV5UfqhUAotveliWUOphN88ll5DZVVTXfLAq/1ftp8
+51/yK8uOWOfgRHsco7shReHEI3z2dbAquL2gA/f9QkmW3UZh9vr+ZX2dhPD
31RMMKAy49v1PS7p2RHFRC24ZmwR/FCdxGmms7ptqN26UF7KfDJHdqYYAOnz
bkbx3ZfigadaeHP/HkRDFuyYQEi/Qv9P1QyGnSZ65A5ulSwGlxzMnJp3luaL
7xnrsqS0W+I12/zPNadqt7X0/O45da9J45iJh/JGXEmFeMzE6iJSShNf3iyi
jkeAPB9l7qxvN5Z+hRNgEP5xl8BijWjxQSANyBvXwGpibQhs5DS2eQEpo99A
fn0oD2RR3NEnEd4JJJ6gnM2/tTb2OWRDj05OALlCQ/8hfeunhpSexSl+uhw3
z+QyP+cjiSnJnpvp35eSQbqTN7FgAr31cS9aI4R/VCAgfaJ7+7qW7kXodnna
l7lNSN6bq/X5FAQNWdolOvtBwCZp3vyyXAk2qmuf2Xpu2lL7H8pjTTZ0D39a
JJMqkQDs+Vi2b4cQdMxkIWmJoPEeqWg1tfo4HvXwizrR9fIVgZBojh1p5/nP
pxN1VbcbntWd0kMmk3AY4UCSCXzNUhaxS4VxfZqGzdBfhHiU8CTa8MtH10nc
L0ZFN9xowGnUpX/GSG+UR7uQSOR3bKGHuUZU/Mjj1uLKAgnhEY5le2xmRKVK
IdIJHHTCH61ibqudb73Z9QarT+FL9LqwP1guuynAZQuZf63KxVlRB2LlBHNy
g4mfY4jJO3m5m5mQhE37DbScwLY40hCTQ8c51LyuTTzhaXqX3XFfoh1VM7pE
c8CIe5bQGzIQ28RRD1zxISc71D2FwiECRlHM3tdWpwOk77/a0jx3/L9ADgPo
QLqAQLO0Wq7ZyxwZik7MwOHYeFAKU4Ha6eyZTvvp13x1j5EHEQpQ/DgXQzZ+
sMwcIeQIUTFOa8GR8xDEzG5cQNHbqUclIImk0ZfBzAQ7xT48JzteKDBgpyWA
+UR75nhicy8tgtv2+PSC2HXYZ1D+5X4m+TtdFX+fNQ/57r6RY3d55dDKuCwX
lisbLghO/kIbYKZ6zkB9DX18Qlh1bHiZQ8tbydsUlypwrfugtkViy0Gq/PES
D5OqGXZL1GvK1bBdQvWK/jJ/ToB1y/d0qTnPyaK/DjZkZVMY5guASza05Pw5
ZhStlDc45WVvmAcoWLKIEI0QodQefDti22Db4EEIMF66FW+nOrFjq/Xpy1GK
ScvyyPMaJ4o/yDQFr27T8WVdDpLDxUe87kcRBjsJlR3TRkYqzNeir2hilViE
aKcoXnsLq/7hjZL5W9NzoUZa793n6Lu2Li18N3idBTUzA7KqLrDY29bYq85b
2IVNiyIPxlTWyVd/hbT9c2VrnyRlh7+NWWG/EAQ86CplYBZiisMDbJTZi9Wr
0BIhCwgypdQT+a6rT5w4ePNCAEX4qHwcuUvlGjy5cevu58R5J51CRm+CT4nH
+dux7usCygy7P/S4cC/vUgpN8xqp4SEoPdSDZOPIKhTMq4AoBMY/g0COo722
tA9n0WavQNn4qyg9ToDwAaOyY4be5nao5Zqq2K3JVXXxc6QDmH6TjcrmsTCM
2IbUful6Wdg9wESt40l/4+kAu8+z/2RcMA7ZugQhFGoIwQg3iSP9JzosMDiU
JipD6WDOkA+u3OXErydXbm5TMMhY9M703Vfw/GMGbYo06a4mb0QkOvZpWGVt
n/8i6/Mx3qkw2OwUhvwuZd1PvMaa0wfae9bjDBpBarfq0ckwDwBP9dZLXnVn
CPSRZ4l0QJ3ccR587JytOok6ZUPJzJfbpJbWhAze35jtA7xc+029n0C5ypHI
F5fmIgzLfsbY4qg1ig2Qr3eZ2ePRAgssenZ5e0lZUpEKRo2i9ob5/BCFXMO2
qXXQsd5raNFIbWbVfl9bqZcv1XpYUdLYxx8GBVZyy/ecfcVYfOZde8mk+caB
cs88IDeDSdhfg6P1UNaWNAeohn+KJFCghzN/3Kz3u2UlvMKx4LDgfn+0C+IO
gBsyQ+JW3kcEiBLb+KrtwCKnFKulvZHdbk9VCjZm5b6eVZY9c2NNBCDLxtNh
sSc8Yw2KofE6B6XS5xlVSsBy+9Shvno9zqqO8BhI707ri0wXDLcVAC1dFo8/
YfQ/1kCD+rNcfgJX2n263cpt86nB9rlzPykWxytRD9l6WbbzfCHrAwHYCTkX
JwF+l6zWBpiFCSxdbA1l0M0nwHGev3oDFlxV/xBQums3Q/ACP8wPoa0TSpFO
A7/vzIRT9w1ci0HliKpeJuAEjO/Kern1SB7xHy3UR/1ZkkomeCPfdKydzcCJ
iJhGcd6eJhCc0mMR0c7Fn0wtupc0KvYHxoc8gwcyMqcPgiJB12Iq++VUT6Za
KiNPYAbVYxDKZ3KiWEaUCnJ9KxohifaopOVr0vIF5y0PBhoN87XroJR42bwo
tFJjkbmjPvcHh2xmHkCcrWg4XxSw2TNubRJeVyOOj6SFPoMu29AtRNTiDrts
WbwAY9tpKbqU366U3uQFdPAVa8qhnmIhOWES2yJ9+t3mlrsaontEHvJsYE1Z
gqRzvC5vYvEIRP5CM+j+CRExy6pAxQLJBNPaEfPg8o/+EkAEU/3baCZ1ogBk
sR7AEEmvAIp5ELlK0Ov8If/baTbiV6ubVuRJ19JEmJMjZuylwBis6TSzcPn2
khethhXMWpRdDDoLz8nFDjh07wSF6s62FqSQpgydh88C4w9DVREtDlQ4cPZV
qczHi/ZHAsdtSwmBqcZnj3cQUMxrUhVVWoA7nQJ+VONpzCJ8zPIA8f1IlZTe
w185BJQ4tr/vaIdKwQMV+Jxi7oXT9747KHHRq23PrqWTieVjD7eVeCfxkQKY
9oY3JzkpqWiiO8UC5JpcaV5cLB+cqPCX8/JGItosRKK5VfqPYcz/HslWxbXY
NnOIrRnD+79fLZkYmIvGthCWuXWau0ZkPLN8yCVel/2MTrU91PwvIzCg0dgn
sCwhdkj+AIzP+vtIafqhdriy/4GC3SqtDqYB+b0NeuodaMan5Ug2TysfreDH
G4MpkIMgeWzownExrDOdQSo0pF/tgvup/RHKyxo5cAeMOFnnvI5TjfgdYymL
C7vn8r9c/ZWoYwB1a1oI44JUqKUJ+rtHFvQEQ+59hdT21yFhRIJufc0B8bIn
aj7OhCp0TktgZhgAeXpoMgr280bDLTZ+RqwGGowifB2xl4K/kSh7+7Ek6ZhC
xzPr/0nDLYAbClnaHq1CVEHeuzKSBs/In18Ea5ozlYJbxsQ/VowWrc/jvIYM
E+gew9Py4y/ovYRPnErSZSmmYo5e/I0HGu4b+zXY+T1oGOcy40m7bmCwQtK2
PGUhpv+BtuF/ShKdygDwhwS6KM68aB+g5gUM3kqdmijgnr3hwhzPDfhVBTZJ
Pa2tNcxxUo6FJg5BRANSlQQ4s88F8I55F3axEmspOGAYCM8J42wrzfut63nJ
8G2BGD2obL1wnb9o96SRoThZbZNuwNnfd+kINVXfKfxxt7nauS8lmUy/mMiz
R8ZNFoISsYTisBDDGE4rJCBbhorRYyERZ4itigmMm8HUh9QM8oVuo/ZYwogC
KsBsPhfnOj4zuHsTLO29cXZDiogGXDZwn5IzQQskP+qsf8Va4ihpnBrzda6F
OVyMyAw1npzpvYjmg+p2lTDMeJClnz1CG92GoxKZDU8Wf20GHL0HUEDuYOzd
nn0yUojogRTSV8Gvpbbkp22HMbpvT//CduuDM4HelpyOE2Tl5WTUXpbmAJKT
SYKwcvhInnjHBjVJRs2Tci+ozD5R5FkVP89zbofno5O6slpMXVlpMAeQOosX
acVzrfljDFnUBwuLa+cnR0ZetqlcNz8fT/8bdRglA1DOMOdMYDKqC4BjRrJk
R3Bx+HuBHe4RXqjiKSIkZtjHXBspRcE6akHylabBmpy6ojYn0ikWRSvIQDv5
1H3yRURMEPUGCcfJf6kow+tgE86G/ucfaElr5eqbB6z3TWtpaxUASM3BWLBc
+Sum1mfkGg/b5lwe3H/TZAD9gddojr/WdR8lQldYQqr37873K5hSf/zZa6C8
5VHAkpFPEn6G26Tq1/sLgcdjfS7tIOyElSg8opG1fGVI5HLmNgaZ+aXFgwt8
5ZI8pLptpXN5OlsOnuTbj8DmUWpPSNE7o7CfsxXzJbpkSlaurmFlPwq/dOYV
aQ6W5AWc/x/2/U8epUUQc9efi2K5lMFSXkAxA9SaEbXNDdTOFiC1jiemk7KZ
h3/pUEupTQGd53Ss8dgSo89SOZ20mMswZhaJLyZITLIUgXEVwc9h9n40jx3M
tQ/Xcl3qvpQ2hFtIGj2Mowyl4Juo+n1KSmAwBvAZasB8ZCyZHoY1aBr+7EbN
OIhS3D7K3DqItPDdiL9rjZkmOUKp64O8AOndXEJRnR1lAl9X9ABTLkaUkt72
lkRnprCF/edX74nD6/ZZMYhgBm2ElZsjuB5mVFA0drZ8D76lciJj/Agwcj9K
+Gi8u0KBi0sjP604e4ZJRDqpvrCcVho/XyMFeHEX6kBc6iqonfCPSkZS1wjG
clexd7r1Z52XjgfnjAFORkZYuSben1M/1Wt1XVYqAuzV8CYBe6SKiI9MUaOO
pVSXGEewyJ9lsnoB8qraI55346nyoWgobNezoOHUmRX2YNU+pNNSg+x82gJC
GG/QiXAQ2IAAwJA9xEUclPNlywnaqlLrBV7hmHn9TQ08tsR29aFvjBlfUEiO
nhsGVgGzm2i7XC0k9EoKNzJGiFKwbpY+6kQV3v6Gzn8fn3/PYL2kvqq3YH6a
4XItZByMYUjHAJtMKsrGbYFofMb2tKVQeFeya3HjYGC9u7nW425E2TfUnV8x
qY0tGT82zDjB0cOO1BoSyS90Gx2LQHbirDewiND8VnkIqVTpjIMkHKUSVu9e
8l4YbeWKVAQ6I3i1EtBsElhJxfSFDoijPcNIrDWWZyIwT3eaKJOLxs9OPlZD
9ElylEYSru2kNtaoasvY9+eV3yS79s3+93Xr054BB8x0XM/YIBQVELnF/J1X
Kn0y83VsBK2XbK1mLyrkiEWb1UZCRUyM7wwFhxfDVqUAKRPZuLpOCmxLfU7m
hCq3xC3TOIIyUX9tz2qsybfSlM+x+2MSsuY951/3PoEZPPfiY+Ezs/Gpi4j2
ySE1l/9vmv+Ea4u1rlpix8blvIh1KW9lW6NNLajAukFeQ6x6dWlBuN/j9zvv
PiAEzoiv3NcjLbz9we5E1PQ156wRnXgEwg0SJnlku0Ps5xfbCgfs+Qb2f7ex
k8dlrqDqcs24zXZqKKtN9V/8+tS9qfAWOPTsL2oNP2fN41jT99NbeNtSk+5S
n14CpSzURqu/tHi5e1Rvc9mJjps0qYIyj213LhdJD0RQUxOc18a0822uFO3T
fveeI2CEeL2kBvpNTitXu3wysNMVDf8z5GfcswpkXnSSZLT2fOMIZGqo+kcY
P3rmgZMlA1mkzZAWgz1q6IbfqIGyjHOzVZbzzNO1Bvuv2qU9y/HiaSKJKw9C
yjdYmQVLExxl57p6L5xHUSs3hI+SsnqXIPPn5THFK5sZl85w0pF55cgPyHAw
HCd8tophThO4YEzURf6n1iwFqihlfFi3RrvfY+ND98HqFaofNtYtwrvaDJSi
5JXelj+O5+LH5Ala0PI8roJi5tPKHHRXwj9W4ZkkXm4EruuITvhjhibNE2Ah
QhvFwCasK71Vygq6rmF98T+2FrXhQfwaZTC9+6V+JZwWYbstPdu64lk5Eho9
dxoHh9QVaRE4zR/e3uE4i4G35We2kAF+LI2lmDPxZ7okLmAB0McfTlm9WCGz
Ee8hjBMqD29rCRgJw+w12tg/ue3PrBDl+515YHwLzPiygPkSetmzo5+hbSQz
CyvFalrx9iPSsrLZ+kgWkYcXyxVkS7FCQGrsddy3TcrkmAoXUBviTW/FlaR6
gpyemRed+XcCEExW9fgChfssNRnu+TJeQfByVGXjI2ldu8rS0Hbm9OliLQrY
93/+6seLuUCohZDPyQznDd3JL3MbzwmlsqhFyYcgemmq1xThwNqi0o+BEGXf
RASJ7OA0753fnw54RFLmoLmIlD0hxunQfnksJO/2z4wT9QOL9323qrOwBS26
AUHCm63P40KdCOnzuRLbQOld4WVRrbrszAHAa1/CfEI3DMDNye/nYGn6hZK0
L1L4qLTIyL+dg+y8IqPgkyolcB0FL4TB/oq38T/m9Tm8GeXrisYkTQhTI6gx
fCSXCnmKZh2Xlh9LW+aOnbO6hjdf3wTAfxoSZpGxagomEGlj53KbxWNSx0Ex
MZJ9+PwI8StrTsddTWIWwmrTiHUxtbst/yT+lLKPRWwu3ufv0T2Ksn0lwH8R
RduzBumIDp0PEYKvZjri9w5g5ETq+BPL5b2jkF4/Ou+TLy5xb3Fbjgs4EvK4
JwuT/EOtlbjSTkLwxw7HwTcVMhJa9soQnBPRXpRtf2ttxqLjFV/oG/U6xzvG
GAPw8ACjmCFJrp+UOruFkEVuW0180GEUV6FdI1gkkAh8lNOIxsFw+kbVEko0
YaD3a8TVs/Zfr/zUxwF7Y9QIBu13xbF+ItGjeFEX62+4NKm35Saz0BhQj6h2
e59Al1tEAqqJ0yceItm0ps9/ojDbkwVaLXcXVl9d7aHz05iY3cvQ/DlBFsPA
R2dT6iE0xwgjdLTr+Gl1Xapbf9cmriTUnENTDY/Cu2GJwW+Ij6Sx3NpzEs3U
Z5holYd2vUuBc4t1KQqlS9HN8Hz+hUjVnnC75K4Qpc7Ycvx+nw8jdjazGfWw
FludkxFq9MUUlxBLqveTNhVICMBH8moMxKbzDgzK9Pr1b69KpOoS4uFeA9Hc
6fDIrVJKFfWaGpVBIyE201ll+Bsz/ghGvYCD/T4TYxm3ur+fqFOTWykcFY3j
84sD9KkAZjw9Mjp8/5szjN4ScwtKBxh8Vdt4fnjbpUD8sKjVOBsTDI5+5/jz
MUvDdTGpU8NLGM2nnZ6rG1H8TtUXYXP3eg1EpXh0vWOWjPauY9FAs+F/pT5a
rhrexVYCtFy1j//+jsVbi71h8AlvQ98DDCP0jhP6OFOXuc6VivWhR1oNxjdR
/i0qqgX0P3G4m0Z8XgXNMjOKssUVoJPl3cAPaelnj0ZO4ANycZW4noKA/VS1
1SNPMj+5ceVaR6MInI7e+sBWxuM6M22UtP3q/AFkwSJAXgY3OifDxw954vtu
aLv58VWXUzv0CmkzXgKx17vyFI+TjicN7Cnu8oL0e79M6qR7n6bqk3zhH0o7
O/8A3a21iB4QGh2Z94caDVnFDcCs/BC38A9XQ70FDCkUBFB/7ewMtezv67I1
wXq62jU0RDByxxob6e6ltIDJO09jOFNs6bLiynaWhUqXrpyOL/JSV4GJM+IX
4X4BZCx2uFXr5XgI2L8WgXfc4n6U37tp9u4ngk5g1NNnB+sKe6qxL15V65Ua
egYtB4iaz9kTWVBzy34VZ3S3ahDPgJm1OqOi5RgfTX1SyNK4zhhy8Xvh7W5V
q1sFwvhKQq91Pp57bg8xL5JK5xXOUWXVGqMw8DVWxbvri4hB3xVgs0FR53ks
H4Cf1KAWcpwFGEC55Eef20O5q8StZB0BppdC7M0kz0qmWIMZv22Ze7/3p8vM
hpYJNiSHwDAsU/Elgh7u7uzFtTk4DBB2cWiOGJ/dCKd/9d0D7MO3NpCDGbTe
O5mcbHCV8GeAJLqlCZL9Sg33SBymhse225j36VhRy+hX0iVApFrUUF8ZSsio
TgRBwSEhgGjhLNrFHNYToy4Q/mbYSD2ie7sE1Z7sLLRphJvocyxnypB35UGf
kj1mcuLiOb3b8QnhgnZP/wriwxEEw9VSpv8rs4ALq9fVs2AfZlXzNX2Wmtv/
0YND5rCsxBSnEzlvDmzFV2muahM4vKJqPL3UYQxFI2ds+f7V3ZxuB9YWZ98h
lZoufzzthvoX2caywyZasLcuaNOZ5WqiUZDyHM9rauSmP1a1uXqW+LXv/iwr
wBuuZJffDiWxyShBCC3Ph6007OcryG5XZ4rOME9SBfFS9QD+Tfz8/ZeCG28n
pdmw+3vs6Icswd8Xm5HKKHpgwdbPHQCN6ADOhAKAvQcKyKuiRjQsptQaoaIw
qFdIOdiY16sMff/zSLnqsoGNT6OyLNTHK4o2KlmlGvZAUgtNj/veu+MGFP5e
4fL5H8qLaJJqSxfAki9yNHPdtN/PP5DPruCuqrOkZ9EJUp0pDI4S8RfrQ6Lo
/5g9Cvg8SrAj67dHA/iAznUw3IciZKg1YpQQPxOVt6QGHB2ToifiUPV+oNK5
M+NmemKtV3HX2CUHH2GYTlHMPvr0ptrkkdZCplk9dGUtYlyifgkr82jjTbRT
t+BFYBCCAtYpkx43kKijXN4J63yUzdkkSdZas+lQhpBM0/rH7XdyMjz8XFPl
MNghD0WUEW0cjAEqvnM10mdiyQUu/R6ofQiOSnPXePsZEr9/gqaDhBDBlVuA
5BeRz/pjQk0lfbH++QJhljts04q0OxKyqLoKGDYVJ/BxwAhkCfJ+6h20BV3t
YyFhq8DYXTNTJjP43aFyMd30fA7SbqRc+JSeqn2we9+K45YT1UfT7Sud1DyT
DRyGGceGDYigvgGICUCAzGC5+ofaSV65JszKaHvZfLSsm0H++xim7ZGjw57l
2swxkRRYOC1se1j9M6owi+FIK50TU3wo9h7NE9NAqgwO0/esCJMsTTbAXhpD
j7AtOXIAfSekpbYzx0iL4NI3dUHVh5VscmG5PBvMCrCT4tOJaBikin5GKwXP
pneGVuqgHzvURH2527zCgMrl8qAwbDU1gXXBerDJKK7+orEvCR/6wREMvYAF
6sWfG+4LqgJFv8bayo6uIJtM9PSXVpWNiA9puGMD99Qt1dpBLEmMQWz2sJZH
flzlG/cPBeGLOBcxvglG1ktzunWfuvV2zUWkslEpkBGehkL86FBrEX27Ryfm
pCdRu8wp/aCvwHJxhZ38ZOFGMTA9uxFj8hTjk4UbkKudTLSYwDsY0Ob1/a3N
IhugrgzoA9G58whxBwvWRHCVsdNkg+p+52j3UyGxCjTARx2XEJFieahDV8gy
w60uFSv/sLfKOVI3h/FX1U2RpcF+2wHOWjTqcgLaaTvZfiTHC3RNQ6KGtjOZ
LOgD86Y8qrwep8K7LM6EMBkeqXL39xEqb7o3kDLLKmPdj7wiSJDXOz2O7eps
IX16hpX1J/cvzs/fDg+b5Q0+RcyxP/mpoxSXz3Qn7OtUEowXjTuHFy5hL0fT
OAeWHjSBwGWHVXpd/Ud8Q8QRik0+/DY5Uo0I11OwuockF+f6GV+rDLs2Jq3E
yGZqUqUVhDRZOhWQMSX3jml6n7scpKxC/1VV/1YifOBYrR5g0Lcgjyx1xzeZ
8W/mlDsDVjQS45W9HsKEK653V+6dqxjZgtyBy0NVpGGv20JJuz6zHyiT8vE1
0uXyWCRCPt0n/JdD7WjgYRVxykSEJHRGR5sJAZjC6dPsv33+QvrtoYZwwMI5
qSRBVBH2AWCv2DyzvAMEZ8Tzy7ZOu0S+gsSwiwYhvr8APNSuSg/Pgo0I0iz8
EayqG6CpgvR0+A4oOiuBOm3OYwcRE2UiktFpwXYwP2nVQLQAJfu/kkVNorvm
3HN2IwhSjmeK4WAWPueLJXMpJ+kNYD0srXcjoHcyMHlgS43s7HesJoLi/upf
gC7AbVupdA47OW9yqjCvQ677GGWR6MFhmctOBEW/Pqyi1TZX3VUwUlPpesex
ureOMX2e/Lagfghpfd6CZL/mxOGRNL0NnAYH49LdSpIU/Ccv14qhJO8/qaZa
He1ZzFkiNfYE9BYj9oEKa6fdboEJJ33tNt2GmLOj2igUh9nJ2Sc6qvqizc3z
hLY/0YHvNLcIgGLS7mxYnGiiBrmS0fckgVxgCoY0f4Bx+xNjAN3xdYxf8WOm
/Pm0cASnCxHOZJn/kAD4VLzNqZQN/3TohzLaiNG6Ola39znpNPqO2okoWAHy
Uzz1SKY6WgkLI694dIsme1Y0lSHSibU34eVWLNFD1CQpu47wBprKESwEjPdm
MryUXAxAQ5uylT5IO2Plzj1uCor0keBl6/HAmsJ88W56AcdGGw8zvgX/fgK9
4r/sgKnc+/RDCAwTveQEadvP6gO/TEW744lLctinH1TmMBTseOcfMKmeffhg
/rgsm9K7hxc7L3ZNi46iUHXWVVesnHQAcRA2FfM4M3R47Uhe4gXt6UOXGMl3
d52oe3G3hoi1iYscPKUWq8KWKJ2DfB/bp1QdsyRKMOlGQKrjaewpljSX1hl7
ib1mbb1pe0EosvoAStTZ5OCu5+bKRAZ6MeXf9VngAr3LZfdu7bENCoL5JVef
lZnlQxVLsCcjYPYdlkIsg+j8OIhwCWpC8YP5q6Vd47YCeX7Du0Vks+O/p/4n
qHqo/safSGFZOmyUlki+TpJPFER4P6sZsUR01lHITnKHgiE91vFnx7cz5jDB
/yU4bJB2jBOb3PVyAg0zjVPizxZlZP/8Vl3VgU+HioCWRHeQPff0L5HdODGt
NMhtWRgoguCr/n+ZpE5u9f0CGsWjpnPCeZ5CTv/zW6G/PKZ+1RSNRWP3wwRP
ou0kzT5avQSrbeeXFqM7p6tSnfwGiU8nMpUNiSkCfNFJAVMgZeuhC/2VdQw4
G8pSszUIqyM/BOlk9fwYqxlDZIQihBmo+HQCcoIaoeeVX1yPtRihrK3WF16h
l7fwZ75lN3ojnxvhuKkI76xzCO4kSTn+Pn2JRDAXv5B3w0ySV9q+QLtjuyO/
gfWTllxmWg1Ku3HM8V6VfuY78lPPfm7Ce1+A7BVG+oiig8gmom18SaDxRvi6
sIKv+R9i4D5J5sf4ZNEJQ7RigwnzdsFJmvcZBf3IxxYZf/HzT4t6eevdgM7x
j5ny+pzQ2XQVuqVhXhw8cXedi4WPcxRKV6p2tg7lvGzwd0qU43AakmxJCUYA
gmFOx3YkKXYo3uHJL41AG/+/VeOKhgXDyrjw2ENDMNdBB2qwjhtISaTF1C/f
e9s7AlBK8yXL3p1hDTIuEOwJr/owuvBTEUphP2ThFly1UardbncOOv2yCepg
kXZoqK83aOvDGKwtTxz1y8nVPJn856JvKY2RfEc7cO4QaLukKvXHmjprJhnF
4KL05WW7C6o8d6mZ9NcY5PN3Fiv7SezmV9Mzu0SC7RQL72wgZC/BWvRq/l1X
HQpzcmV5iqrMQ0zYbMD9zxGokjvK0CqGVkqMzZzcikgPENhPzyxEw9P5rKaY
3zkccYT7yx5exMxrGHX3atM+ijWtpG5y17uXbQuIXewnDAIENebboY2MsJXw
1I+NbODc3zq4ahhyFWgtrZbhyeDv0Ab4NvsjAmvH0XzVJwyCmPTHhVHDSgrW
7VyC1rrHRFa25OXFo/4Q2ih+hXWwSyj7wI+JyF/Upwa9LQn6FHwEbP1wezlJ
V7HgK5uK5Ft54f+adSmb9UGo0vYgSUlkw5gIfIixxO+VV0sI5VeH/eRV46BU
E3G8RyikbuY2yhHdkescYXRvgtmYhPgcaerNPRJQnLI7I3S26zARIIoJvAUg
I7v+40e9hD/tp9B3//6j5GkxyjZG1EGUVX1TovjPdE/EyZAgpYxD2oOkxu+B
itItxQ6NhkWxQT8e96t9D5lI9Nr6/izNaETEtfb6uAYy0Jt42ThYCgw6r+80
2kUTza3PiYRhwfSMBUK/VDt+mFGImPrluHV0vVXE1GXI+vA7Z7rylWdlUVIb
w3mx2tYAr/gAl4/qKlmvt86ouYDQPzpJaXYkeltejDo81hqKGyDgVeAwcsu2
r0WTZYMBQ4zcR8pOlfDdqWZGZDipUrxs/adrXbvMbCpz3/abtXvAhf0Br7yJ
Z97FZ/vcJ0gYY6a+79Z8AukxsAHxnbII5T5/Dm3h0oD+ooEt4dqQrruTbDJJ
CpRGOQiBXmzRntjCy6njpfbG+RoebvzHimVZsL2QcKrLpQPF/Bi+8I+crXK7
G3HwjWsrvTiSx/xg9quMBaFn10L5iaBv0VJE8u8dOcKbPipYjMZxiUi2go9m
uy3RnTb0W/N3/Z4XX9d8iU8rq2nPLWIyqSgYijFIcMv/+O0K/h83cNGclMLY
ABcZvX31Yxn9qRYubqRc+rgFU/VQRRrv4lBCooKBHe8xTwMuIVMgw/jS2+7H
ctGQIk5g3FhHfq0OHatPWyNEloQDReTtI6OnY8hmOcZnilWw/ED7Fw0MfBG9
GSQ6pWXLthL8vCC6tbjU1xIixe6MyhVb66rWl+MUn1km64Eqb9rayMEyk5W6
1yThTOlR1NtKRmo2vL49YjCns0tkL2FjARmSWrEpml01++NUtZe6vZA5lkZq
3l0giQ3YLSGja3KA+uuaDwVkfFyswk4mRUf7F5FQqm2SyKFviInFlZfy25de
N0l1VI5NR/klr8OgOs/rnYv3qUU1iYajpIr/o9rboHxMKPd1KVNpXkZ3SQua
jLTTvXQAmkVHwUKn5lc3AsN5InV2m5DhocdfR6iW50wbVGXbyv6c60sp0hmw
yab8xcuaHvytLL9YSG0SNlOykfhrWjQxVUWZzDxPVHJbvY0dz6qzXD/sHnX+
it+dEm5sjUb9B1GK374ZB2UbeybItxkl2VpoafTyLoU56BU6kg97/9wapfmj
UYP8CFTzFDp6/4savirjDlqMrP78pdgLPJzsc06fBz0X4FBJCu8YHZcfYDv7
USogJOPJT0ix1rD3nbO8KsepHqPsQqvkG58kaU4Nlv++6kx9Su+WpwsiSqUa
rIaEMamoY8nufJBGyVvv4fnvzIJ5Es6cYQ6PIOM/bcgBx8vOyMut3ypbQGLS
ZazvMnz7P8BuJB/AJKTqbnR5bB4gJFy2iNDWw3ROvIb15u7iwHf43/OsWhXR
PcK65880FousvJoGYB03phgGKz2agnURMdkqZKCEb4O79TC75WBRb4MhCiIN
d3dq6+2OzjkVdXRRmfJLvEXcuHt1JjbnKp5Pf6e/8MQe+WpS3XO1ZQ8DZYbF
lcjThCe3cQVOblQw+HNEK2pLER8DP75VwUC9PgrpDodHjEjCvoQ4WZboy9CJ
aaMVttHrTduMtN80igrvvgKfkD7P3y3mM/donLroSmqrl94FDTnKPOHUB8C0
K28Km3tE1rIHWh0DdZ1jFr8dSFSVKsKOBHOturcYSeJnceVahCJjLUt4skoS
i0UE1R+hrDkcAW3dJfDLyVHmW3PfybXLeg8k8vwNzNy0B/xFtcHEcPU0RhuE
1fjmWAEPc+0YLYaF0DHd5Dwi4YUZQMW2idBBiMZUvbubcclKIODTd2GlwsKv
kvpM3TDOVL+VJwp2aLWdW6w3AEECNZ/HAYbe2BOZh1PiZEzTiBgBuFnKD0Wo
0tJhnjoWcsFlJizAHaiKkJr/RfKSwI/0QFc4vRYVUqYwzxaBilsICOQVXrl6
Oyr377sJV6d5h0EVNxyUkHS1AEogEoqkDmY0PK7VKDWPg1aTc/81nETTNJdz
FwBlLajWmSgDdxilHzVVxokMQE5xWcWPCygNfYVe41Pjp2gSw21CEqfN8mAU
SDxf+rIpc+pLYM98TuCriGu+i7dnHSH0iASki9F/znjMtHufT6BCZDCumWyt
wdrOsz7I39G9wPkq9vYwiiLln092VV4FgdFnzZKvE7VXB9eaUeWjPsqdCd+o
/+kaQm3DRvGXP6YPX9JwYwYMeaGBZzf/3EHBCsBa9Htqy96muCQaAB4WUkLJ
z4FEz7OgtinZbLknXcJHTSsDDdD9kyDhH+1buASXgnHMuImz7+4EmRGiK7t7
5QhSS7ClimWgYEBqsgJWhtNHRGgQYVSRHf6P9OXF7vxVjpjoiFTjovFs9TKM
om5QcS1I4M1vx/PsR/P9bJOMVQv1yeoYbcGFpF1SpNy/ZWBNOz0YesreV4cJ
OIRjqN1L4BhX3ecOr14Ic6OaWisFh8xKk6WSA57R7GvGxxPqExKiq5SB8X3m
5n5RtvHGJZI9DYzu3upFWzC+5ZUwasL3X9W5TMtHIrkYAo99CWVIFnFPJ9Ma
GWi/wzZPO3jqJVb1rjNjIM2vUlQXMwFxeHTLjjRZf7q6Psf9h7zR6pq82hW1
AmiYvDrUO2k2sbPgMO/T3dm1bx4s/yEILjYZR21+Nain+9IiqEY3hj7nbHLC
LGZctwPD41q2o1PnbsCYfzJYq47lrlDur6SqRiUlGRus3nxXybaN5+3BVsgr
kSZeVz7F+TTzsnDGMT6s6wdOh4WsCLrYC6rdZjkpG5Ch5uczLnA2vxSoqfK8
W/3jwJWV78RNG3Ie7Su1XbI4iWQGRaCYVlJghKo78Uq+Ofqdfw+0LROCP8kG
4zCKFzR0d218N/8Rut/YMvuLR/ylpERm44Ez5BvsJ3CBCpHcR8YQsU2T0iWm
IzBY1NcGXEVedOu7JWIeFm50Ijo3Gs8Zv1QlYJFA4d2TdbcOMHXQBpR4zU5E
fIeK6pHl+q1gUJQoSs1zhZvih44pqTtC5wOGBADiQ7v2hHXpt7wNmOmzkRoA
i/Lal5a2FQfoQpWir2RQ4D6NRCR0vXsdMG1kaDLoEuGkfkgJntCvbU5zNJ9T
2LF2r+u5TmTOpmn1sThnMSdmi99FJWY4zbX/1vvYFuGiVQJLY0+M9U5tIY+u
FurP+Po7ed3SAENqbUKwK4W1ky8otWv6jnZ016QuBKfKls908HZS4yGy7aiN
/qvOjCIxfcALQJSn5Yk3eH0OMAjJ946BZBrwaDRZkU2UBgyzHDK2QAsivAnK
WfePPS8IiVCdbx/qKZN9gfA1wMWZrtDcczRuHt3P5cIhypFKSg/nM0KIj+NS
T8pso4C7Jc6c8jp1CP7FBEw8pW2Vh6kyth8z9Hr3SIS2aWyA7N0Gt/RIvhru
y2wMU2ZrVgTrFELVDi0o4OaNtR6okztjfnR74bYSN1bN1AurOF9yj2WNVXWH
1IfBov9WLqik/Q69WIwqkjXGoScVzjqtBprM1809RTcThjvrBBoPEOmcyRoH
2lenLPq19Z0BoRNEeUkvUW+o4oKuEF7Ujshnvel1uz/A6VMmkDd7Mp7MH/Gt
i353AUBpeC8WmacllN3OIAD60X3Lk7aFMFsccttkel3Glsu7gP2JQqwlV3Oz
iuXEnauihMhgVyj7DvenrtcJu+WjJ3z+WUOmBnehAvySDceqhHAruJ1c5CYY
NMKHvMQFCxEJ+8u6rLn2MOvL366Z3wxeHaTRWBauhM6oq1cii/PMlZFrkTjY
YSyknVRZjTv/tKe5u6ntUFzvSbiStuuMrewjoQDwFbddsocuV40QNb4Kk10v
/xA0+fvuxWTyJNZe6i2uMRz16x5hd9WMJ+fFfOy14Tl1/wGClirMFzqmznG8
2PwhOHPWgIApyDqMBrkXkrMz+bTQtCyfzugAjY610LPPnBMFVefn+hN46ev0
Em1MLs3SdhlLMi5VdhAP0WV9Q3QnpuhbdymIz6beijcdnP8m4W6yQd3ajQWB
tUHI5UbMC0viTHFJ7T9fSLEY1l6l9uZmFWnBazhRJOYrlRtZaGG9HzDo8jWv
Qe+1u80MhanVja/xTD9PQFpB/d6mlPdUJFCrbymbvOSSqRkwhS3psswySx5v
IucxToHm+32gxRp/u4b+uTkYuC0vktzwZK+GUULSsNh/57BeO7C7DLMlkJ7P
FNIH9tCQW3EjULlZC9FqSnfr4fpgMK4W2fQfgpC8yXHY5reorWARW0Ytngki
f2gITGye7ioUKeqB0wLo0M8MUEoIYdEuMlwIY2yyGUrhE9jmnjdRjjrZdHsg
SoYugWkZkZ64l7/uHNhhLFsm5Ik4m1NveDF2+ZdzZDbYSVFY9WnK0UwmjVSZ
rgwc5zwqPXW7nTh5mA1o35QcY+D1g/8iRkjxERzHkFqtmsjiTGc4oERMKq7M
rcF0Nc90M5uBJKAF7UGoom0ROVXdUC92ZlYpYCzJpJsow5XOKp8TbuJaULEp
WrxjF3Gh/rr2jUytqCio4Xlc5cYB5BpdvdT/7Zs7rPQmC0kFm8w2/fIv9G+J
Z3nyFOoKcOCQ4bHULg3vP+rqdwb279tnst5XTueayxmTAcEV4QtS5wB7D8Z0
txKw5wuQI+5tdTTUUFLsuxg3dn/a2s/kkw3JHOLtrFBacfWVdrwUiu2yoazt
1gapiFU09vqWorjSYdoAbjaR9ik7D42nEq5iKo8IOMK14tU40xZCl8fQqFAH
rn7R00o1Y3g5O87ipgVTsIFRlichzJ8BV3cLTDGGShPPr2fsmUF2ytTPPWqa
goey3FQBbcwsrfkjMxENKuCQcJm1w8KiR6DKxJpP14peF90NmD9I8ICxPc0k
LXgDn2mLt5Os2NEQEHtB/8ZBWGOKt6lkhPOuIdyuqtpnwBd5oGAAF1b3L9xS
vq2TMR+bcdcFgPEXZKjvKlbRGS5WXJHmp44q1srEjTbb+PMNSQpbx6DjBjO8
FWHftRI9pLHeJJmBnjhqbi68jnWIM9SolhVYfOavkYi5O5Y5oIbkN7suRJ1g
zfJOe9NaAcMKSi15Il+zf9phvsph4BE7CWBhWnQTNiApTginHwaj1s0y9/Vg
l85BcB57HuI+VM0kfA5b9YPpVnS1DKt3ycD0Ff41CZ0mhs9J3m7dPHRNSWTQ
y7lyPpnFcPNhvZlquZpte1Po4qZKe7o3kAr+ZVS2dihn/eCoC+zaX+pihiz3
/PcUf/6/u4bpO0fvwVDPR8PJNjI/vmH7BHQ87Q7F6AXED5AONxa506cmbsQG
WqBkUM7RomfjT//Ni/4cegRCR6sHcM8nY46BnTRK9EDCp5FglaNUxb+aQDUn
zMrtlN2fGo6CKwoNAXg8LJ77cExQQBgI8u7dg/pBK63AV0w144DtYo5JX1pe
WMt5otK0++us2TSz3A84BeV/G+4DJa1Jpix4vcSZzkvK9fBJ5sG410z7vT0X
gz6yGy5kesqw/EzqPO+JBHlP9wKx2S3UHSyeLUYN1GK4I1NBBHNu6wENMDO5
32ltlhn6q0SULfSi2i55lFswZ8TOq6H9C4CvNfcDG9zSeZc/FE/LwqL6DJ00
rahqRtNV/M0eic9F1oZ+8YDNkW9DsFAFgPx95x/a1MKks0iOjvAf0AGfVu0w
VlZS1oXdvS+wzZ79KGzhfdq7p/iddj2YYNItAHIOjYTa9BRcpuOSpY8yyQ5T
0uyxoPG7De90dJGvSHg1BJmn4me9PXvJE/X2+tPXyYnJY5xSlOdjDxvX59Qc
zapC/lqEQvxeWOj0AgUXuPC8vqtDkPuLQAEXrZiOMJibtcOefIkhi7oKZBpJ
ZsgZ87C67QbHmTKX28xySQnmT8h+i1JZRiEfVHnzTlOOb6i5oGHTKasTzryB
nmMsY2+iXhccNM9G6T5Cdqb2ThZg0vpI6Kk8kVpkSzlFJCLUGOg1WbVLoEI9
G4wPYF/4DpC+xjtTdSo1WxKiwgbDwzu9GegJ9seRANVsdZQkAe1oAXTZOSkI
yfTktxwPrleRqxjBRT6+pWZe5ODMbMJe1kR9BRSSr4dPnxddFyJziwgK5TZY
pUJ+qLW34vgmfYnickUTwh7e9KECxGF/4PQVKL6J0NTb29fMPU7E8LapUTvO
lmwi6bYtyvojzfXHzQM9oKWQlcz9f+2efSU9I+Blqs6pRhwU4JjW6g6o51q8
tSdRheOVA/gfBIGKvBter7mSF1HcMkXoqpqVHe26cjlfMk+QwfwMNFCD+cBE
TWhGLn1La+JbRLxKp4TVL25I07I5Pi2rj+Vnpk2MRXK5I3nhwJqAzSLMcKIt
J0aIArqMvbW00+Pz40k2sFjTmsC1a2IEovmiwpEwNkAUJ6PsYV5n4CQvdL2z
vBDz1Pq+ljcV7tsQrz7g8UaymWOqK0sD3e19Jas0pqIBLS1PzOp9uzhk3OJw
AvjGIxCibSLXWcP7+UL6gPA6ui1KMOMpvRHg17nGu7SH8lY0f5lEcTPYvOMg
ix5yYXJwE1UHS9jSFrgQFKhFGPbs07IF2PT+2NIisggldRuxAEr20rhthoNp
sYCRiwOE2a7IUHVvrD2L2lK9Gafv+LFfL1ZGAcHX9VbhvZcqPfy5UMkn5dfx
qvBoMA2LUh1Bux2yP9B4IYN+GpDL+BpdJlRfFlJqZ3Arc/JsBEstAbgElb0h
Y/Kf8B3Mw5BXxIi1AD76i2L7Vu3fxtSYVv10914JqZwIMFM3Fsj+i0xc9wfQ
Pu9js973yVF4eVCeWXZ1ltc1SbWgu56v69dw2iE/QSSfGjYyUu76cKobelZz
m7r3MKy8Y2wZnqhnYNy5Yl6sxc0zwRQFqUPPZxDlue9XavL8k76hRXtkguOr
lNmku2LoRkOmVM+uMWfGGwy7UFPrpno1ruIx4ajErgd0Dch48HeJRPo/hJb/
+0IjEvl6NHme/dFWrB3SQgKVNB/AfFWlXnAAhQ22PbRvnXeqy6cj+slt51L0
3++Bjj4cnTO8MvyTOx0cYv3mTrHMXyX+dHFgllt6UDu9533UbcySJTTd2/U+
GE9fslhQrrDKCW5HuYCJvS4ZJZLlszInU9AyAcmRO58FgBveVgHerTzl+tEf
1wfooaaWSs2lSVCM/PpSYOKDk/6TejrZXjW4Mu8QoqfAjOVyC6TwhwVFw778
yPVjXEGrrdl4U3Dour7mFKR+7CmB55WvgLJTzvD6DKhHAhjFx7RWn6r1NTC1
AmMeoy+cINm7ag4/T3Tb5XbCXOJTdCRRVW2h6SRn2lPjm1bNJSBFhyrm1JjD
uTJ4mj9iyjcHuoyOjbEaN8u8jsE9TxNBeWq+HQaMgV5D9o6Ow70RbQgfkVQe
NiQoZDigVjCr/6KPJv5Yy+28lvF1r6gROhePn+RhxDTK4P3Kaz7ZRnktE4MI
qPAT9rMsENc29MV3CDO3htdeo6WSZngny6Exk/QvQSxRsOq1Wi1bOKLzG58r
Wn9adJWPhvQyZiExxZxkrVHjIBDsViP5HkzE+B1X8WXcyQoBrxuX0hceXb7P
FllmMk363LOItGcnqsVOBkrqomQt/1BDg1FQEDvTj1MPS6XnU6ZVYGzcwPKE
FF+J7ord+7X1psueFTbcr1GOefAoZuDMqla6UCPdwzoAtF8bAloUlSzRwl/d
en3IO4JR73njHUDu+4dqTAmLcTaA/Q+V+xEYoWKt1MHTFQuqAjM2ea/MxF/d
zvMIjfAAgppxHxKD0EtxrsrJ1lj+gfWGfPWRRgHbpIPO3/LeO8qMz58n6hbt
1rR6v8SR9G4RtIiabPaPQHRKLj/qDMoexBzogmUkqBQ8FKzFYPodLK+gsYug
FEccgOC7YcMFPkNgVE3vxf9exjXSFIPSUanRcl0Zz5gLdnODC0NJ+HSTqgbb
H46drSUkII82QuS//hD+ZwehGKnDcrT7kKzB0STGcFe3LZ11ZdwA3qpUyUvw
Ri6WxQmC0jrWpd0hmQU/12ubU44YIn0+Ooj90nTVl44WYN8bWnQTBYMwh+ZO
pCam0AgrlnfB2u0qBiHWRnzp6Vx/MJcHneJO5nCVUSMNn5BKRGz/CdaYqx6z
ItHur32fbcF8xk4623qEtSmzmegiovRJZCZK/k4ljjKTrz84BqEDXGY3qE/w
P2iKgBd8NoBz5PBbOdrp6GU18rusOcEqCZSJcLj6bHc87uiBTlTJlZ/8sVKe
tLU6yBLLCn8EncUAFYhYJTwGSeKF1uv4UU50FoGei0W1oN4odAVOmtnc84vR
2n7dI4Wo0d92KvaZSuyfvOc6wwSkavaFq1C2AlcSdwLkyW7vuW081dPoAvO7
ASvSR48Bl6qtZASoCDCaUVO+k2/09JsAVbpf8qnNeydewWF8rpsjlXnGWW/r
H4CGHsNQ0WfUY7YCYenENvwXAjogXnIWwXn8aNZl9gR6m31NXtnWEIVpMfTw
gzaeO5Hp/3sJnPBWvJ2PEzThCQvwUGdQEQTFc0JLwMeWR9UMZKXWM4c+XN/0
b5GcreuWIyShHpnXJeeK9TiyZbxd+Xn+pkgRAHOQQg+pDJhV7yxb/xg30uBi
hjNFgwF7XDn3dA6KvQn0BLrYPMDBL54TzfJbl+Wh8K/S6Z+0AlOSdAlvXM1J
srPdpPjwszamhNg6hb2ExLDMbKmjEysuI6Kwn4bO79AcQ75qUGcmUoZu6/a0
A8AlidyPesRKrtQRxhOqAQE154kT5oq4QNgXh7inbr6Hwb30qkIFYU+t9RZ9
l2giCPhH/MvAeIMt2Sk9bxafX3NlPUSQV6ijWUoQpCMUSIReG/pSHYnBX4pr
1B2RjH+DgP8aLsumBKUOeez0iIlo683MX+JImdISpbesoEQochRTn4l3+T8V
tHwVtwa7EjhXu4uMWwaFFVzSJ9gmgjkJLeZkpMCn04yPyjRC3qHsqA4hL2kN
/0cbbIosJSwSuTRsAV0ZEEGDR4ctclqJpR+2zSY4BMnjnr+eY07ALcyfbHFX
xF/ElwqlekjEXEMfQarOoM6uUEOxMhwWzuqnDw6Jsp+fV7/ImkmjqvIdfUjB
V4cTJRlx8EdUb5yk6AF40l3T7neeyAcVdIOkLqm3CH5aKzVifejyPVZW/bVw
/r4FKhmqYXyyvJlV/LIQIGBvvBfqaIUGtMyf6UMm1bi9qsm2cnTFVLnqvOFf
58u23qnyE1Sufg5sVUpjULAwTmJBLx2/2BSObipKXlPnu2XF577vrz0XP/56
XTd8ZbuaD871BRywHbKTpeS4QYWcdvc1cFFONHIa+/utMW2AXUXk9F1MFNhA
VRAusM2ryWlodZItFj/yPHqsJ0NUgKUiLbKqaoCplZYoqVanGTNAIUjU0RxH
D+YHn4RP1aHWi7QIDOSU7xLprmFTO/eFnPSH1YP35ouXqoE1mGZ7dzDprPrf
dGxWrXYeKeHz5NB4+HYVP7KJlOXK6NJ7ObKVK+8mF6CpJTk3J9m7NKwxW81d
QHg4co7drqkNF2n2BFlex/4XhrHIshZvqS2Gr0r5HPGX7QwK5/EsBIUry2kc
XYltbn0WyjID2gc7Ik+OoHQwteJgx3hAAAMG1jv7W81PUff6bNxpJn7+v2ML
hBiLbnHg56XP2MPiaHfBu0RDEFgqCSlKbbOgeInbwRnv6c7k2YMshCA0vfko
wfYFjuxZUPDJOFufYOml8q2u/cTYN7sxAYWqCf3Rxg0Od2Nndd2ONsMWQWs8
qxommD0iJdHWiNKoMfXtQ6HTUC3Wuo1pFG964gt2qij1tpd1HrJ8tLVEVxmr
lYqUjy2F5IT8kGeJbb8d9gEu33zXNP5S42NlHdoZGJj6tj5tBANssp8o2v7X
cC23TeiDKAl4GGFJIV4CJfp+sl2QBg1cRxG2zxKJ5EA3t7NExUN86OkRHupD
PJ6RoCEJNbHMpDgV25WK5gEZjaIw9mqBIlp2gPRoloRhCSEbaNHLrdPHARE2
Fls30tIqaThEnHlDDwyhNSXqwwz86AnJXI7Kw9ox7dqeZ9bEvx5pcu+X89Dz
rHDDrL1QJByP2/JVCG7Vg8F7vVn/DA8gexxuxs6JMNP2l7X2a6ORkX8TkQlt
jdl2YPpBn2e9sCRiaTyhKpTCRp5GvFVxYDcQPjw9LDPz/unysoNk+BPYoE2s
Sqn+aO/Bk6eNmoKvaq30qoqJbFITwyb7dLxCQfN5lLt0B1KqW/U0eW0C84sQ
T2vT1ziQgM4GPfhBTdlSZU4Uio8xRSiESdqhDDD66tDFqhni0nh/NlELkSXT
c6VRAKdzyod5kTQIlH1XHIRX+SEIigNafvGbGcMO6EskzIusj3x0smEC42rc
5XGrjmzlti4lYL9QMCNZ7TZ2lZPyHxMiD+E+4rqfrkNbqgx01JVxly327t3C
lO6wHnuUBoiY+RIv6/gAbFvr5cDHDVMkI48hclFujwp1C4Di4DyVS7/33zQQ
0gnf65VDDLsMxuxgn4sur5DshcmlBZ8mEnqNfKk3QKpwRmpqergStwEcCv9P
t2h9Bzre+EdVuluPfBuw1SD8cR/qwfh+vIZ0cg4PdgkiYsQHMNQZ3rA1RVTE
Dn6lFXzIxEdgvWdaas/0rhxXp3RxcMFi/3KEcqfgGlwdikZshuhpheQYyFHS
9ovG++fquVCuRJjWKIljkDNXoY32HzW/4x0Y+TxOQUZnabLTaZced4SRokW/
ZP2kiCUe7vmOJYxIpoz9sTKNPhcGtCuqrcEVxCzZI5YUEOQqpg0QnqyMzYcR
HQ46u9M8CMgu0rBrf9wE3DbbGJq5FmSjh94Zp8H25e8YF4UnOFRagBb3oda2
Rxqeh4XWzXjEpBUw9KrdiyDrz4zMLKvE3IYX3ZOMhZxGaJ7asS/kQLYiRwP3
6uLSVRv0BBMAOv+lBrvgm94vAEPU5wFN459H5f+Y47ouPgilY3tejuLMKpej
GXeVXf2jxrr3oNJtDQMEEWOmMWRI+07Arz5GXOVY++NYPJtFnVU1PdXOIL9z
iNitFKMpWN2xe2FSMBgqHPa01V82r98nB0uN8s8YXC0HZvrWkrQscYVOKqEr
JPTZzwdnsJyZsNzndlKz6pw/ui0xJBN5BVuO+eZujjsXF8FSPE7QyWtyYsSt
t24l/9YTDIp6VaYnm2ipx7bf1J/+heZUFFGni+YopVN3g/NDGzM9vw/KoeK/
Z5cRoFqK5MrleacqivRicUucXvTJta69dcFGuCCmsQ7UoYqGIN6ojrvavABT
44jV22MBjD3YvfsyabcdYOm3MjAoXYAE1LJSE0XQhBP1ORR3Fuf0PXB5xD1K
egKvRHb1o+5e64fWtywhUz4fjyiDI03Qk26cyMzTSFuH7hhhgTmnsNGMXUl8
80OGEeSzhW75V+uVZXvgt6lYbEqbV5NPpJ/vni6vcIBu5f3ZMY2uyQNzA6P+
PuZpCatLAYQsWzVdvhVX8v2iLwQq9JIcW/SloyqXaJ+c3K7IpBSH2NM3mheY
LBYdcC6yiTdggd81qTh1+bJnkD/+ziRaQXPTM30LruBzAn72fSLcopJ0KY0P
/Cewtg1dQBuhmrNWM04ip1ezCxMWJirRUypMDjvywzD6Qq26BazrkDd2EezY
2TykacS9GEzNV4CBxpW1NvLImQbgiAmJix5+2HuJ1xoXTuldHEjgwQbUwrQ9
8OnQRfQncj1mXSZZBJeEy28u0jslwj69Rpg0VUKC0CGyB7HWAwTDws0MWjKx
EHb6WxNPb9qLYNZQLjFemmHqaEMPVzvmmdW2yveTRQ7QzcUyC3gE4+QdEsxa
IC3P6ZvucP6qF5qe5RZBHPX76/VnvYuEnD/VCvYTtNSrUFzKb6cImrcmW5aJ
ER2qy/uy9Hx1Z8Hjy2M00LSZCs2O0yKvZa2Zfsa6A67M0xhGMRne+9GFr4lQ
O9FdkAny5UDamIKJkWnbLn5MzQdMIapazEa+W4xTwtko4PM7/WSjGyJ/yoCG
OJlqcSgL7dHvNJfz8kbxBx8UEHF01tXqZWvaQSdk24jtUAuwd3V6Om1m6LHn
3P8SuPYkiRsb97Nueidy/V7qlF7zp6M0UX40fVLXVG8Vma8AeO8B3809eEIc
9pOm71tKnDP8KzEpXCcgikbOkcPo5Zy3NUtbEDjImuokcwyiXZzz7QIFJkT8
hI4Y5QDaFeCBY7vRgeJxbm4BsiceaVVL3zw/Ii24kwMxr2wlXNQDAEw2n5Ju
4KzLZvYvGshwczLc+3xPnztY7dzQ11z0AxVD82GtnaS1sPAqY1amjq6ZTksh
rQF9sFs4p88Bu3U8x8J7klxzvz6VXebCF4/nNWeRAh1O9/YALNet7onYxTVA
QDBKY4/doHuncWF5b67g6F+eLQrBtdm7QIOAtzxVdrUumbHCm6MHN8FuxzFf
zSjUPpUCn8vaCvRXfrQ7v0ODofwI/SXXEgbZUyMuES5BdkVebDF3N7snTV3S
wWZLURzZV3KTMaFEMkzrBrR0uECClq0cWrvgnJNGntao9VWP7BPnmQoARsJ5
WEv8JDNRJq23X9TPaiY4fsMnW/zVT0TcIwjnUocXscV/mLFWoB9YqiQs8wEd
TJ6Dqodd/U4JvXCOm37+MapiTb0uEJWwWzfhRwRAaco/VzB2T+ACSLJEQ/PC
Qp5g6+CKlwOvPHVr9wckhpPx3pfd9XI9rteriwlG1KcmJVhRowmoOwvb9ZXI
FJ3t8FPt4Q8MmaBjl5Q8FarHkomKWP5Ec3fwse6e32Fm+NlMEMqZsesY9fpY
vHMCY6v0sO5UMHQ2LqxnYBq9cHDKjzZJH61nQ0xySlco6SlVJNeWaxiHuXgh
UmI9WYPuj2ZyeuyW4gRaQcSNxUxClSvft6fx5gQdVTuvSgCAmV/gXd6hGk4q
LxpqsJVZb2RFw69NXVa+VSfE3NN1887yq0dRJnuM9eIShJBRz9ZrX70N0DKM
TH5JvitlhQ+qbDD1/tE4FoNOmH0EkBnLrkjnJPAI6DKLUHZRbmFrAYma0WlX
2KSbh25/n5OLQu2cngomQy2C+54ILC/e9TBUF+TzrtScv78fPa/+H1Gd65ru
OZZGe0iz+vs8wdPwouVe5Qu9Dtm80MJ3qYD43ipje9niu//RYLHmT+9uyF8j
NrKdNtnEL+6R1dPJGu9XwjjYtDyi8e2tvTaneyAO+n7vEGyvWXGKvu0AdpIK
5zHWHDVbC/1PZe2mbi92ydsRb3wNFj9K5mFsD3FUaoeacFZI0CUTyPqq9KE1
JDc29hDqUNYMRvMdPTTwIjg/hAWSzJRNxuwVS+FZrkGIzAvQNnGU2mCEqMUR
3Fw08kzj5xlB5nxk315WPWgYaN5ttDXwPu9aiF7DSQSluRR/P5stXykYo1Yi
f+D+Py9Tiw+pvx/WVoiADOyiRljS/6A9ZZmv5LG7EZ2REVHa+x6RR1OYKMQW
Q+QGtVir0m7e0Bp/sP6GXZsPcKAUripXnMZifnraj3OdTfRy8N3fOofWRMiR
wdBpF7lelqzWNdFzv+Cn/dz/a+78pkIV746R9M7I9ZlVcahHabRQWmFyZAcd
k/fD0BFQuozwBT97ZQlxqV4xYRnzBEaTFVB0mkNLQLDosUkNE7C423I5E9yp
KqXIdQM7BlulGzaFshP6uiRr7a5CV7fCVBnByed3NAXUoNAPQxH5aDOc/sBJ
nYEtV4GIR+lp6Ygs8E1ZF1fLi4pcUojuzjYXkjjBJ7/UZWRvgA1QMq6RcooQ
2fS+HvhHId0JZnVeQd2rxGXa1hAN28rRUneXzbMKIyfD3xcrqReJuJ4eyD6s
6WEBShcw9tXCOjjJJwl2fqZ0iFVu8B6y9S+Z5lbOmwECeaUxFkWB2BFynYzu
n7uVftaFHguHhEzeiHp7WUH10Ib6bUeHwNz+jdzzRqjV5ErYWpaEl2m1V4yP
Q8PibQKEeLh+PLzf+nPQMBbL9cjrOI53ZwMkCW/ppFi05ieK8D6VKuuXu7Wx
3S4L0tZQoxqe4jfTl8iLbw4gM0XgMeaxc9HDmYSTCe64gSVNQq3a7LDOCt0/
lDiDzY6Z5yu5wC8ajblFfZzuFZjtv0yWnXYv1Qu6fgmMF7DXRCu71v231EFu
p3r0PVGQsInNlTnrqBDZ7grjByoVVwnEqUV48ZR+SS85+QOjj4Ya+fzSUXtS
OscHV33Z28lI9O7ToXbNhuIZP+6tgpKm7Vymrw1LMu6J9OUW564socxdl5Xt
s7vUEiOapuQC2cqgp5i9bRZTgCZmqIzTiMgDCVrXtwJ3yuflQHMI4A/JoLBn
KbxaLePQwiEBov3+gS0cjark+/bPqVL1LkOgBNP7LFgaukT6EEj5sc4INh5d
mBeDhMQ6WALs0Pw55cCb7qwlPXV82fpopYfjK6/7ejnBdThErO1M1yFs6lah
szAVaarfK/w7sL6KHLZAp4aJM/XJDMTqJA+MEP7R0O5LXTr4hVbFYbxEVxU7
mlIJAWI5rVC31ae1IsgpijCRcKbHrwgOVp6IYPQPq+00Z/14IK7yuWRY4H8v
IGYRRNq1rln+haszx0zUu/i5iAQ4/DSZ0rbGS3BomopVDrgiE5su5lszhP+z
6AZu5EigUDIWspZPohszcBzwHlOMJ+RB38k4yelEg+Edv0KvQp7BF/e6JQvA
bLgnToz4SfWXzOodFKoxW2eiO+5dRG9/+JKxvOQdGNBn7UDyuRp1BgYSqvEP
NmScpdOEhBResI0k/eiIKiTms3BoI5bo1VrWC5ZbfiKWULjqXtNz3KIVBwYw
2keYQzlQNQ/tabP7gykuAYGP3w3m4EcIfAKrOmLWLW5hukm0eEvrCtpQAlrR
vbgy8OGbRd4YmUSvBdMEoyHH0MUBVJKmw10LAjSfHkKrsTAxWp+Knuf2vNRG
VNrzGbGBHtCF1tVSyrGjVz27pmQ73Nv43MPqe6B8JcNI0LedyTyqXaNq4YoY
n6R1tfVRsP/CSNe8c2xUp+TqAfaG0nbk6EnqlHQkkft8vsbSFAcGmv2Fv7OW
H0x9ouz9A+nDLqGgoZa26TK3oSLZlhEpgF6zcak/vxSbDTquYsRXIw7d43G+
/QyMdK+yr5lxIwRKZRbEWOhJfyHhu888JR0cJ6EwV0pI81WoV/bxuSOkWaNQ
QCjAUN8KZlmd/MVSngpM+xwlf8AvTk85bVHwKui/EqtcC0SBK3sWQ5iJgBjL
04I9sXaHFt6yr/cVwIXTBeTS8ADUNTVITVFfd7dt0neKzkv8dkVP+Tsez3VL
7CxncZNxRt3Hcyduv8m1thf8bKk47E7FSe8Qv+lYS86Hhtf0ukGqvM7TGmR6
tc/2T2XxzZT1I+L6YUUHp4+yZJixKuProKugPDF/sfBNCaBvYIz5EnWzMlL4
95xak2cE7EZKe//bTSl09FCVx0zF4/XcFplZeUD++RBSRiEnTb5lRgI3veDM
vU8PuDissGb2RP0MmyqMviDuF7viV8FIS8UO206xN2HrxMJmQ+S9ZzV6ehc5
6+sI1a5q9hdRaM7nbZw2xEGlMDX+2X38SJ46s7hGuQXZQ2G/EfW9LPPMwwhW
Ug1shxqWQyNxNtQqx0pzLSb09ffhzuzjCa7YA8wS+1BJ7O1mikvdxgnE4DcP
aRNQ9MlXf6TRI8LjQadzg0THX4nbSmWxPJ3AnMkc+hYUg884RCUYw65hUyvv
oom0IQ8vaXh0D7jpqfciC+x1dluKrhBY4I991e8552tcDMURYV5J0KEcSV8W
6lLffKuD1HGy9HAPTcCt4LQIwlhLESTPiGuWa3ECQ1v9wN8yNg4pVfHKBhR2
t31vQPILTnuEm4P6WaltGj/+SMHTlPb0lAvxZCS4ZwiY40x002xMFyeYrGUe
ghDLIGiID+aKojb5NChI2T9evIRhdJjNnQCnWtIiKXyD70GQycfes6wnhyyq
UOghljIRnlPaWsuEtUPAjEPMlZ3qhlCyjzc+W7wZwi57BKJMAc/d7pWabfls
Hj4uUiP5oo2GejrJbHVLmu8F5pfdwe01jdZ9CyhVhffSonmpl+tZkIJOKkoE
Ft2W3TlYMoKQKti8RVM8+upoXiFQdBneTDGnZDfJHb+VaxJVMzLWop1P+JOc
o1QeokH4pl2ckLYBhbwsiY7mnf47+hA9bZmxDLNwj22rUNTQ6RjecGMrJxCf
AhvVYKfp6jL4t+GTF0x/PChGnSQl3i/1v83qQDqeN4PLxKOOUHcU/Etu8NtT
oAaPooqNEmkste2UnGnexpcLh7hfadkSgJuQRqQVPJyy+ND7Br+V0NQYa2V4
fAKddtncSn4Vu9ImlI7D4aqtfIwcYu9XbbhybaLYpCOeu+JBQvdD2PKK+a53
ImlfTOKPD2/zXqJj9dZ4MZr0JJz/jsiJzuz3HagVxJWhO5Z2q9uH4HugY3j7
gTW8DflKu1fHwyuS5eTqSwdgNU2doylXHubDVEssQrIs8pO9Mh20n2mVzFG/
2GJMs/U4bDHVvqB+fIy2FfjJD75U9fxE6WFqSdszNW+J4eGPI4qi62N+2+oj
NONBeNua7h0ZODu1mR1Pxyt0vwO6yN1fpm65/u1aqK43uJ6Q3CUEN787y8SD
4I3n2S5qFrFQqJqsHCuZw7Q3CT/Ss+o5vzblDrr5nYDR19eeGbO7fQO1xgrp
dPbOuJpLC8jlAi/eqhGacoHKekAQO7tIlVXqusgFSiqU/+djoIZYLu4GtgL9
M4nepvumFAty/AlvwlULj9JBYlD5ndjB1HmstAcRU2/m2YrKvfJVFKwkmRHS
EaAUcfdfZGx776rl1LjZ6aXx2NTWESSz4EnBVLcbQ4V2TaeIvSUWJqjdootg
h8vcgpnFFqYY7b5bjNpk6ZDpIkALoYHt0clOeJ9izkzAsisQI0H704K8h1ry
5BAlHWpzVNqwyqf1m2BwtOyJeXa4RG3fTZJUaKR7E5MpKn3Wj/JFeeUVdUBM
vVFG8Km07tnrc7v/Hnr/0F9HXrrt3MXJNkw9DxPLFlZpSl/9qCJhWvWxeH1U
SqZzrqzwBTOaz2J9yqg2w0FzBpYq1yWAE3Iur7kvKkiI6OUGVtMH4SVpJtVK
Rw9fdYzvJHjf8Mm31As8PUwCXoXG8FYQrBnOnFp9Vp37ix9ucjPHCHFvvAnK
Y8vwpfU45x157zl1wDtKXKBDahCfX+2wP1qnV/QcyA69Qvx4Yirn5HVmnmjs
72u2eWgJR8Kv7qtuuc4dLAUb0tGSTvzmvQgRlSfHeFtjUcQ6ahgJ1iMqAHps
8IHhZUQd6GFedDFU2WMBy9fU/4SGjTThgzvvi+a3d3OWK/M8u7I3EZWfV8mh
1YUlu3JYfQpHgPwc/741pgciTxd4ZuZjuKcV7bp3Qoe8fesZRJv5vvJh1eoN
GO8t43Sdp0HE80Gbgoe8GSAFJMc7ymhaSdk6oqvE5c2S2jMIxieEMH3QiEk3
j57Rb4svHH0o4pHknMvyvLIbvMg+ptD0gGbcpAbBXLjs5qykb9rAj002ZEzU
W8gF1Xa25BMUicDc+lMA48BaEKrM3nx2+DSkbXfv0WSj8MEpRtHTenVrNXDx
uuJoS6zNv5kEoycAWbzHn4Id/OzmoEp5OpeYKtgoglXV9P+4ykeWCJbgRUwI
WjVLdNcejh9xo7kJiupdEPdB+KJVTsu0O34JYnUYPOgApJ5a+Ul61VxgQis/
EBtyb4cBJDK7/u3La8ML/Q9Iz3f9oB0kMGxhPe8exszeIBGNnPeBVcq/stPI
ht176ErraMZ1TA45OfHercmTBeQqZXa2weYW9d3kQvOBpYYf5BoSXt2amKSS
MkRDLVLdulK7XLr2O2XXtlJk7mrjrNzN8Mx8LzN1ZlBjN7pxHOsXA1oPt6f6
Qgwb5M9q2Vs6EBqe0ineZylyipRDziaAJPsMA3lzWdunzZGDCdZAQXbj/3Fj
LRkdUd4lvo7pZwz1AXXjdew0lprgcGJiYZlX5+fmf4xN3/3ZWrQZ+e2IFoOH
TxQl4R4C40MPE6hgNWk9hHB24vU1vn5oA5nWGOw7QbL1NzXXW9jCHnL30sDf
xcU/fjrWbD2qcGIcaGGwb+rzWQUSH0QsZJjJgwO9eepeT8do23e1w+kVAGIR
5T49rqD6bq2RCmHxGjloiylIHPvz6GRdN+jC7wXNUKoYlQ8urmwRlwCU+Nfg
nb3hvuIByMGgTkdp+pdBa1Hg/eEARHwWX2c2qcqZQ0/uCEOviRXXicxej2EX
zaVgaRrsjmQRJ+uGmIFNlL7nJWdml+UxOKtGkIlA1wO3WCaPXePZd6cAjjZ6
LDPvkdcRCyIL5JBMKiIqVP/BYawzXdj/A3vz/Urx7KaP91LQmn8xE+BmGfEl
BhvtJuKdaBbBgYpwyV5Qdty2wt5e8hpDap/fd8CxNZElWeWVYTFAAhjgPUBM
Tx4pzek85g5niSbUTBNzZFSiJWOVFhDwhN4Yp7axha7fpq4GSQQWt+kZ/LDI
RLuRf6hWBmCXKppI8e8aAOv9JqXg1e4IE1aOYSLWravx9RlHZ5LQYRTUk1uj
6cWYwKwas4a8GH1VTjjBvPG5G87BKiBTKySZo+nzeGMrvHUptb95LfQ/qg4L
fom5OOJWYleTcUIpr278XNIOdHes5hG2ADNZ+vji/Uws24+TDrrLI47v1HUz
XzvCbqRGn21+eMmAT8CpRBO20XbGXOwziGUt5JNfc+JTvhVeSL5f0a8TQuS/
8FcVLphxKMHhWMUi4mav4UkVF6QmRQZFzLAAd//tyhnweH92ZMjTeLjwT87u
DkXWrJY01DLwW4mWNWBEoU2a1XDiAB3BtgLAVs0m783J71W7IO0cgQ8rmMG+
OFi4BM6CP2vJ7XI153vatPUbGWZMdCFqvrobx2i/ixQ8+A9xiRwP50QSIK+Q
ujwCyi0Gt9P3sw85eZMLn7csOwhgYkGKhLOf07/s5OOfdovA4Y8+oyBXs4fB
+4bn+c/otB+WNk/rIw/7RkXEB5yrC2YNZlaXURsXh2Nku0wap62BA+bWWYhb
s8O1uD6n+utB9QHovUYuoGQa53q9p/B0N8uFNZE8tEx9cpHICaXgzGdugrAE
XwWt/wsCsTifTwkLtBsgtiWJQR6WNuxWJvMXZ/BGCnJm+A0Q79P5bipmz2Rh
iQePs46dhlVxAnuq7AOx8R9fvBRupWD068rM6TWqJUs4kdlIVp684X5gj4Y6
rskOY+wcc5XE0qYAjcJTSFBieLIySOLX/lGcKpIM7faC4GgXtYXjUj6jq59/
lAii9aOvULQocUBr9rRCIPstqFnRmlHRiM3grnzO49HRvzDZhOneN3INUUQg
ku+82l6msJ6cZcUimJaKKoHZwTITMKswmDMRDXewfu1IRMiVYgVOZIuD7i5h
CyiYDS29EcKkCOjhabMkjx80c/gjwSqbtkb7AmlQ4Q/03I4y6m+8LrEx5YCH
blqKA+XtoXgCvXk9xVSnf36kuu9lA80fBzsqfdFBFyv5qr6GLgq1dEhvtaDf
+vcl5PwfqKSwcw6J9rssJjFveZ5rk9peCMJ46gBw4xvnLz7NBoQb4fv3kyY1
TsXGjSRmRayw+toU2B/D6ucu56j44pmsxwy1J7HeHxgEMTA5YzkpTuSCmQ7z
PHZyGSOHeLJD0bqgxZ2UXcz1ywc7f4HG5uIcwIYPPZfcy0sh90ug326vOVl8
6bHZoAjPb5fA9JTfiBsBRi0Se0vZ7TzSgPuwJvwrOAPjCMhZTrNd/hFrzutX
fsuJjDZUPTwi3ccvYjvENIFmGTvfZ3iaqSlZW/hRoAI46fY0SBsJk52xfgSi
JnY3AtoBkDH25PgFQ2wPuf6sQIisVG8gC59NHjat8oJx0gAbo1Mt+OXJwmad
9ugfV9YQmWFA3DnWNtIkmvjUz3nJS4qJ5yP7m3KUfUkpCLxw5OpF3o3ANhEf
/RZZFq6aX55LUnrfMJODC/JpfoqZKm6PAKbAqAwOKzAy7WwhTdbcKPGjGH3l
5A5y6LG9kyxfOmtF8fhl4AfmFs/9bTG6SGMQzY/REKaQ8L7g7rQecySUUFac
DyaJGnE4CN/BnWSFAN+E0n0XYLqQnRbzG+So4LQPD9s5sJIxHmoxqR5gX6jY
rxkZmrbUa0BvJ52Nlbo9P33quUQo2n8RE0OGLETJU+XyH54CP3+xuIec3Z58
WWHcAi+evv/lWfNw0pypK119SYmTvcMUK3CD6ptU0j84WgaVtRnjJnkDtwfc
Fxvt23rucbA7hQLXE/GdsDyfPF2PzFZdiX164eWJ24wi5O2I2XL9Oz7OK6yq
sz8xw4YsoA3okl+jCjbgwFzK0Ms4Cxzf9zHzZX0H8KTI3xapfFWdbuOqHF6D
bWd4h2WsNpS7qFRwRr1oe/xKv/svJKNSoIMK/+3vOcEScQ3lRqxnL6Iq8EuX
6so9d116+5dvWlGWfMftQKdx95gePn8ut/FzX6gQA/FemxpkMb3OpXuW23Z5
HT4hzejQh5Ijm8DHUAZii/gW0mR+WHfqnvTrivEDvpQkJ4p8SLArfdDnHeuZ
/pbbcdgO3GcDHcTBZMEkV9m441pkngoepWc6xHiH4WjkyUB0akPBnOQFd6wv
44a2FAGkCpiSf1eJI0CjYB/QHI6OgQu4qryl6aYb8oYhZGHJTwcTixIOYe0w
reSifieqBbr58g7kW16y09Y2I8684QBODCM/M41FtsHzKkZjS7SgGXkknt2V
QSXV7hwZ3EKn2c/FGVRgJE8sWqKKjVKjshGHz/ItttliaEQ2ytw9TeUjcc11
LxB9sC0Q3ibPzOJjpmPynp3tMR68X6lYP7FA9mZKmP6/ZAS/7wthitMMvZcH
1h56TcWljmagyIQWhfL8yDpEb+UiqINVwkZJikvMgZTzqT/eXB53zUi65ZNL
574L5HmapwsAoEGRUZUy0rcP/a2tcoP0zaR+rMZxFuN8uAfMrHLEs9qwlUmb
jKwN4vgXmEcTEQAUbGuC7ry/p8y13TXB4A8iM06jgs2HGhvLJikKAP3tLNay
CrJz1RN7ZRQyQNmROxLmeoaMuKyZq/CrTvyz8eeEMv2PUrxlyG+YseiWP/pg
NDvRBT0W7plILwvh0QaKz99UMgHikWZnLOAfceJkhe5oDVz9Ffca0ZBjoxrB
uIprRmH08s2goE/3fUCp9o5pyfQbJHGiDUgtPI9BQT8iOQrOB9VkuffPgoB7
J9bRNW5mdcec4BmNdTykLZmxJiVRs2t8NCLDdOgYOohA2P9jgByABd1n92U3
8Y2GmXqhigTC7mBjMD0JqMBapkjq/vTVTIKeCybpO/rvDvn/QPiQn+7i8o8s
gcqUrJaK8X0bD0YpTh5vyWEe8dNMub1zNJnMngnskFsDxopyhTQjpSixh3Js
8bPOyg5lCTWx1uV0t2IJ/K/3KCNAMo0HU0pqeSxTi6gTTjQjt+zd7lLkGu8q
fPA0UJXBKgZSovwHNfZRaeWD4ljwpAFf92iT3D/4Mj93avgaaJoPmiDaU0S6
KVuTo3b5JanbGaXXxkLmLspX2B4pJpUwwlwd6UGvzZcZ/JUDnDZYaqurqLz7
cK2HzGZe+n6TvTO8EMsUU72UIpVpDGQOrz6oEBz9PJlRCg8srseiCmBvrg1I
VXWRWdzKlP2ljBnA4cWwRF5J774ILg+7IC5mFCQDnGPykE3c2FuosVBWlRqJ
dqilrGuG0xrY4NG+5vSUmt91sgxxkAEWXTHNsLUTOMUMfihDyFepz4gWUDd5
CWu4qdlPM2LW8dujesIopODPOkiLE6OXO4CbVZDsMDmjEtv8zFOUAoWlySbj
z1t81cBqnEiN7A0rcHVIRea7mQlyqs/alQV89sJh6FrVY40d2eY9sKTNAOZr
Wq53HOQR0P4mNfdEYFXpAfUbtUJHJGQkycFikVc8hXw3RC0og9Cc6oMV4Fr8
PXXuno9Yqo0KhWHC6jrvbf+BrNKX6kQthCDx3wtfqmYnWzTp58eVjNIvuhuJ
GSewPwsyuviWjw220AU285oN5dTzOn2Ue0mtA9uxm3mRExewWiHgB5xvIU9I
gfvgnt+jPC/OR0rH4MhXlwhywtWnULsJL7XOXE5bfVzlsikqlEVJ2JzyqHPP
D8qxwH9OfsTVGwNLX3Ry0nAI8p4N7Jjo/7cCoAPE83E7rch5QnL96Ul47T/G
//58IcqtxYng0fR7D0dDbpnF8D7U571FcaUzoT9iRgoljPU7ZzZsKCJgrJK8
uJHE6LgR5LUq6fhsHgQMadhlSR5cyfqqD+QzCMmEIL3fr1liqpbj1vNsYDjb
hLjOZkNypZTkeHhKvnUwUHU3jtNnXeqHkV+Gd7IEoEx8T1G0TXzz3GfULxn0
nsHpAOXQjJ1AF52hFoX+7A8wPApatUpUn7dCm3bA6RQSlcncnkYvLaHehuXm
C3NRgIueodF6C0P+la4ZklioOTQNjEPT+I27QGwboBNlSIXXng2ehHwRRHMI
9mJO4NY2H7Z0BFi6rqCsJqu3fFBDxiLhBjEbdnyMGjVWpZw0iMdd5EBucBQt
sY1cVKVimSlHk06FGsRGFZSibR4S2JvjmlkzK4hAAvyHT0erj8emYQmCTCd8
FVZAo2iOns++FRTo66JF2qPSfZPAC+hhfNIoqz1PFE01RfeOqpziWaDvnf3r
wAe8YyYKDpa4+i3viJzIGvZQM260aODEtbuyLcYO3AVkODIwBldMrsUROsVm
1pVrqr6j7AjolNruTX/lzE1RbNecwM7DqTaPD6fKadzqhN2lk2+Uk1K1a2Fk
sFMoLcHJMROg+n7xfQVfGHKkCPTNmiV2omn+j3h0eRKo9X0V2xYERKd2kzKO
ooOQT0EMjmmgOySt7sGqqn2HYiPIQzrJdbl3fOYK+83OEk5d1YYm0G/Dewie
4xIuYkBJSHslHXs+Iiv/jdCVAZImpx+EsFV6cIH7FSxHbPTbgv4ee4wC7yDU
lcnRwZymcX3qQWa5XHRzinDe7Qwos9ckfEBlD4HSgH+GtABkjWJdYczAVCTk
eaUPq9jjQ/vY4am9QOZZFoXajx7jNhj99PeBEkXsxz+BYLNs3ZIcEoBtkP+r
tgNnbOFcHJ39YAFHSf2jdANHAKtW09JY3nnv7Da+TeIYW5ZhFNMeclQjnqCP
DydKFxlgpNuilpiuPAXIZZzMHWc5q1Y7YkJf7XxoqJA1gllzOeSIJT8UPR8w
f8GpYITdDivCKwGE95qZ+Hzutv1Ux9gT2Jy0V2JPgW/9yYrymm7L0ZD7MRKC
GTYQhjM5f6C84WX2LH8bZLn+0qdy6JNKVVkKQL0eejs3F/h40eU77f05pCOE
J4FEaQwMOKUddCf2OGgMt54KffFykt41kPuXItwVn1djQGj7hK1JfZPqYEca
XAThMcHZHdl/M46iJCZs/NqIUns0Beud+OvTK1Q9JLVaodvOkWg5AFGbCnkO
skcYux5Fk5eiIQd50c379ZP1EUMNRnAMsEl9IvPKcq+7nNvi8jJ45gYl75n7
jX+XhrmN3nV36F1sHZ2dpadUjn/580U5WgcluuRckU1k99C/hcSNPNYlEbqB
+8Xnv+7opBe15j5IHp+1P31BfV1FgM7l7iTIRK5egPvgSyUmNKN2VXm7X3I8
5uEVhkpbjW4wLTjkCBtYgFtIjSr6gb9vslxXDVxMA01SE+mNlCg78eH1+G0d
8BrN1KKFUl8vOYJwayc92/nLxVA3rSGiTh5raacYBdiM/eNACErphnoIPQjn
i9sSlbuusw1ocSXvzPSZnoiO62Tl4laq53oQ7fof52Tkjl5naB1/x53fsATe
crfcpaPHKdqHTLshi9gWg8ITk7zMgvQVX+y9OQ14Go93s8t4UCKcVKc87jSo
BZNA/6eYWoU4Xaq2loRR6digvj53xUihObd/pImzXi/LXdqAOzKWY8sdMLNT
wMxfIzlqKgEjN/9JjeRc8AXKWRup+U9H1SwvnU/olOGKAL4nEjvtCrzvi0Mp
oqcYj1QHZ9UCQS63FH3NgekkJ5o1AWIH3/7vBU/j/ibt8y3qKMB+GhFHkQ9S
+aDGEAszn/7172TASGChcmFPPzUYEyS49rkOQn8QsFbNOzSvtghT+IfmyEpN
qcTv0J0iXF5HjBBMZxaTgrIOaAJBde2JtMBy+Mv5H5ig8CpqdqOZKL/pULpq
5Orj8U4fw6I9ulohuw+QqWabQj6GTi6FCTnC7yX0Xs8ycQRZy1o1fLESVU5o
kHq8nDF3BrZ1t7l1AcdBpOzCl3JFGBc3WuK1tgkSyr1FNajYUdICHrBraBl4
ukR4RRiw5A6QXA2wt31VsShxnre6YmO0uitnqX1xth9anwy+VwzTnvSUYEml
EgkgX9qjibpFjPa832slAv5e0JX3nm9G7fo2icFr0oKr2pNYsUk6qkhhAUcP
dzu5CuF8swnaU0nkK7/nF+kC/mQ0rZOGvTTVeU+IwOO1Zb2UwJvJKMUNkJw3
pzBQJRjfJ8sQR3xqgtkpnSJn+igxML+n2nzArmMxsOZv52d/aqxmiewC/8GV
T8qdvmN2cgi94CP/ZJeRb6sg2NAacARsIIo3XWp6DTs2tJ/s43A3yrtBIUzu
Xlveb0CZ5JtuU1OSz7iSyTRbzLn1F7s05Avh1XfmqijlnhmJe8WgV1xiDpQF
oDCxI6WJr0NuhXKyx/W/rKEIoRei6byvuKAJSQC8TBgnBXS257rhZf3lwmRP
yfsfbGtfTTDgSM7h7WbvvpxKS2Q0lMJGiL9eIHvGawj2+3Dw24Ck/o1Hblqm
Sw0T6yX0IxHZwchOuP1c4wgmsq0/N37iwpsJcjikZkAuJ3i0YT9G1X5r7z1n
Ki4KTKvSL3AmyCh7H6b+WE4wTUdZlJ1sSEHjTqaMVhweahfBpc2lcRHPvpPf
iQUrwI7LwzQdFFiZDFCg8AfbxhKBHwHuZ/eV1rBUNvlQoMQfI0DHZh/7orDZ
TW1E0KOM9VsGz9SixfBiD4bl3Mttt7zS/Wpnqp4ghjjsGDolhLv2luy7zAxX
Zr+7q7zxgeHO5thEazwUgfC9+hOE2VNExZ0bBUDF812xTrIw3xyMu8Gp7Wak
slVobVXI/grawAxzozXLQ6amaSgvqfpz4jzr6EywzK1Fh4nqlGpCndZ4Q3ON
4/kNQYcQ8D6q5NzOTXRKKamRuobcVJwx1YhjUKUfOMNezD1Ed+5x+puzMg7Y
pGfmH6cg5Q5rJqMPQYtX1HN9kAMeEwLEOoQvF1rSuJykXkQQSmrJ5ND5Flfe
eFEZJ7TFwiCHopxIKIP/X6xT9xRvUKH/MGgkHaamDssAFxgVsXhnfMp+IEXN
je6du/pYtuQsOV84LOCiyr609Qfe2d4uRsgbyZS8X1i62GPLqYTM9yHM3ESJ
8m/bFGr5UDc7kaNvl9WiBDMwZCKKpT8nzep5+ZyYAR3gNzwWuDXp9Y5KN0W6
E1BpiYlyZdgLtqLwd++mncKgIXztZg6YiOyXY46tp+DhVrBI577Cf+0KsupX
Xie/18FlrlVZTBunUqIPM2SUfcG43lKr1lfEGzuENYLubh9l+FMaePPsE3KF
Zr8rFCcmSBkMWbi6yeHGNsB0qAZYcaCjwSzCe5/Vr6agYPJqo5bvHB2ZTCgK
R6l+w1m86Am+0SfyV8/jKuXh4ejei1OUr26X+Q1qNWtVgBHdNrYQbeoPAMEV
8+E/M4PB95Malhw4nt/MneyQixxTYrHYimrISFClEX4nEYh+o/Je4B+nNRRe
2Jfmw0+dKqa/UZ3TfNKHCuLNo/33JiuLQvvKjBWAswyWUCvgkx1VxjW5DKod
epG+eEH7Br5qS6/FlGW/bX/U1rKNrDTciBJz2qTUr0JOjEWO/h4U3+LC3agv
MFOsLqNBK6GsDHRqllEplraYqZYcoM3o1b/331kcslBBkaDrMPl6DJWSR6ah
CQR7skR/7d2w1IRrgAhJOLTnUNphwZ0OCVpx0+SkjDmzUvAFlBYmAwfo2bZD
2UfSjwwQSY6raJDaczutjdIPw2mclrYw6F0h2XfvIuQnZfqCcT9nFXBo7SEo
tOgB0VyDHlpd3j6ki+dxUfOzdQ2Ju2tfiKXDRSr5eT5qrF5WUsL3C3Fgj8l+
GSSEDZUg/7awtZSPLOErrRwlwcJLn8hcPS3bBdQoQpCbPO8d0PFNglbE4eXI
DGecYhSgUP1YiIx3EcrRdRH6BFNz3BOnINlSA60gA+2NGRG1NXTAmfdbq0y0
Wxoswn/IoLOyGQDyXNLbGYJnuTnptPl6Oy7CGemHEwnBDxmCQ52zB8o7Mwgs
InyG+oemap5KmId8yzH19u8i3xJCQ3d4WMEArLd7Lou2tpTCmfpiC2wX6nt/
cvNfvkIA7zdwyN0H08tHCW8LlvA4CnAyO03J97vO/f1wG/KGCY26wTaj9sv/
+PyRT2lPNf4PtGk3AJukqbIYj3IjEa16dnv7FOGLnWO7DnxcmOeKW4lxF20H
+I7Y7N9N4fhZYQgAjvxVJSABmivtVtap0i5NXQEtqG++hunkvjPxvEVtCl4r
ciU7pK/erq0HddxfZIurUIKFAjeMT0HMAytgDZ4a5ZN0MxqSMUrMp2lq5aod
VQsBNRZQPCQeshkVU1WsRs2mzokYa/2q7FZkxIKE5XcQdtSJPBtuFB66nB3R
8U7qiXKK12P1mDJJG8HoP1B4PpsB+Aacn+LrVfC/80uhAnLyzrqaclxRRT76
qKy2dQreMjuRQwbQam9ldT1CWOc6S8Zj1Z3fUM790DivJaAH0wH0r2iDGaC5
zKUn8140M0f0AA0erAuUvP3sAgF4nKzH+si+ocaqJWxpry51V2AtGQTKDoSi
Foq4MvrSncTy88Hr8/cKiuiTXMEbddeJ2z0BBYZVdkR7QfeiKssrl5w/3Dha
TO27JS6QuH/JTw3lYMAoh1413gWkeKmrgzFa0rvUKsXw7k7Zw/fvspgwUkaA
9i7Rd7NHQsWjE3KHwDlfZLLcrfH69HxquLf93Nu8CFIPSCa16eVJs/0H/tAb
Z0rXlLMv2qMOWbtbRkf8W8UdB9QoShJTKtL9LnV1jeuBV8FWdkobFxJtEiBU
e8wGtBaIvMCf2q5RFtcxT+FeyKAvwP4gAVLrrVQTCRRKJDHNn9HVqrpvjOZl
iZXGEGiWYTVcvuBpLkbJ7YteUI2l5tmGsYCSi3NMaVKYbn+od9P1gK89b0ef
WN3mWhf7CYvz9+xtrAjtWcR63W/rcuYs4EebWBuAYVBtt5Asi8aWy6lGfh9A
6EoHThyvUhD0B8eL0DroBfABLW9MyrJkdO/koodotDTARIxbGA+uF7yQ7+ws
6g0ECt5gk5Zhz2FVGYi8dfgjIKrd0UOzPPyesRfOBb/7vGsSDVzbZtGzE1Ix
3C0jwELPL7KrisEmB2ZoIMch3nGS/Li1WOiqINhhBxhWx8740jQxdmvnJA5A
HaIGLH5jzCvywoNGtxn9LRX2rwwRI9VTeOAt79n2rq4rXV2XDDaTMZE2gNek
GzSeG1GiP/9Mt3jfo/0i21qzao7oo6bTnm4/q6ELWNqlFIt+fR5zJ+ABlpbA
Vf3CUk8q/KQF5weYEh5AbyR4HcNohmPS4ywhmqEdqBrhknctVdRFQ6qUDJo/
vEqs1umc6WvLoY4NR88wJylfsmF0OGQdgFrVDc+qDZf2jRaNpYo6Jud/hnvk
pSU8SG3fBp+nBSA1voT40dpCQ8n5sjtoc10i9OlxOyYKdA9UZ1gHiCVj/+l/
h37tgSbRYCUFnHTk0hWOUZFv3qU7h2HLRrkZPeAx3Lm65+idYr6XTZAQ5pF1
fOmPGGmzi2oxEiOwqfW+qBoNFpiW4jKVqDk7EFyJ1uKfPWzOIpJhdwIi+LZ7
Hi6uOZ8jJYt4Lobfk/yCQA7o1s75aSf79OHatZNAUrB6KVtNMJDQDUR58LHV
UJQkptmU0JP+Ul4qeFvoEg61ywx5FosqL2drXJC/+NUxyJCbDQnES3Cuz7D7
hYvsPVTvEHGgu0tZ3oRtONKxZosaqH65jFufJ7UNtvAFnIL/fmQKdafd69tk
EsXNe9RHy0Nng/GwHna8P8FXIP4QlEl8jLL8o74KCYAXU1qcCpb2do/KqvSK
GMVsqfBF1fXylhfJY6CSTTsk3+rJay+aD2bEASVag12KefBlxaxFVz8iHeSt
Jgz9K42UDh5YqknTeym0bmAnWLCv31Bc3142lpbDA9sVWVkZ2+0RRxt0alnl
Ly8X4/SEG8n7Q9rb2As9oLxMURtslT9Hofp/QWmijjNlYgN9E18f97AP+Nau
IAAV6XLXRGz5zxL6LsqwLvU+j4olxR6x/PXpPc7KGsDtSiAVgvRfA9XrnCRZ
0gUeCibAdaiSV6v3gAiarr1omhDzHxhwmwbvf8EetorzyCcdbbGkfd3Em9gN
h+IgD2HtPX7MCXUB3r6ANX+3/mVWpIOGWslBzMm5EsgS+cab6Xpa2GPG1bAc
uh+NNudvm8bZ9LNEMJREvfJdjKPo+83Rxui9jqJG6UO4dcDS+dCpe8ocIemK
r6oRIL6rKO8lvQgujTuCzBlD2o4CABePUxmsXxYTIgdUEH3rN8zGPInvg1MG
GoWQouiX5mqqOo5o9EqXO/6xb4yC6TVd2eFYG49uoFI6DjfWkMYRxVo3tXt/
JVpZiwYhakUkSDArWVN4WlQOPJAhhxpjGI5kA6YJ9lRuCB7DfTSdReqBBjOj
9QxnRIKUyeHeVioprzCWE8STbfDwqzZv5Jd9yfy5d2xFRkb2bGsR/q8wFyEn
+BU56pVHwm+GkmurePGx1HyVY2zeMlhC+OfU+iEb9BhNJ7NJc9Jjae3zZrF8
wC2NBCeyRCqSS3X4O7ymnBaJPHVNAUcAqxY3JuPcaZG6Ic+nSJ1yB8xLCn2D
EU5xAZw4DjajmLy5ISYxWa7kxZZoqbNj47nse4XfoHVI/5QdBvCPol73VRM5
N1PCVbB2Uur27DowOrrYkWrnUp27QZVcKQJjNIU8CzbcbX0kkTf2fJGe9EhB
VZw7CBGA+YELHnLjmQBUi4WGSFLqwUYwXezLsvgnli3/CsqX/4L1F7lwMDHc
f91oLiIHe0yRG1fTZyFYPLQye+wb3BiHgBys/0g51jy+3k0PSsH5PtxmvEFP
Tpi6umnyJ47ZJrTq+E3MwGM2LexPhSZbOWl6Y9k7874aJC4CQYYzhp5HEWmL
PYtKryVmNMUfw/V6E4xFDu9T+noA1szvhwodBvEtlKOvq7dtP2gmNnzGYERv
bcmKdcHHEFOHnjozxtKehoC5DXPBiSFXq56AHrJ+IqD7T9wXQHEtRfO9/Ubc
lArbgRZWtK3fmyWv91cRqj+IlS8oPyb6mUeOMiX5iTvoubOlVCtoJv2JKkbo
vgJv+Fj4DaLtzLYBCNB/chJM8ph0cvvG+jYDc54vc9jwSvBRgXEEj7RnAos6
P+HTBrcjIoJ9JcptBwwshbrpDe2wsNlyUROEZ7mboKoLZWKjSFqa5crTrJqz
5+7wklhPiqZ++PYyLFhd3qhOgpYFBizHwwscd9alVUelRti0mYA+mPItjD0u
EIqTJTXjDzHp33L8FizoNdYJ/cfOlQlGwlNbwRm6/afL6j7lCCYSUH0coeQk
hbcX91VO5h+HFpWMNe5hahmt9OvwvcQGj7ANrUDLHBnhGcr8cFd0nBrhTX97
9CCKQ/7EA2PTPVMieCCXEjszcriAQ/R/wmXXmUdSChZKo1PLG/h3TiahGQtF
qllAicx5m2HrP4tnM+O1T23uVX/VvMlj6dWLdQWW6ibQcCB39M/Mdbf6mzl7
S0IteoM+lfKNrXCQ+OBcgjlpluQdu0XnWtVsRxdfqiSSVIMadYE28Dsf+CLu
T2D8O9gpU8LjCuD3uyG6KMjZISoFRwCUjqGPmfm1kY0XRPAm8mUNRYsKngUa
UIFCZ+JsT6JFy3p/2QCKqfyNYtRFvBW/uzZZdeVaFr9sB79nFqMyLZskQgjJ
c9P31x4lzedxzNWZy1ca7CnBHJbsmvSiAcos87LMNmyFIWKpJ+XvJuMSFC1s
maHQd7ijL9J/+2YKShsFCkAIW3DOT/aAQGm9L5tkHNmuQ4Ukg0tRhp7gGaga
UdQaYlau/3ReARRVDWLOh98ajwN2X//OOY5A2c4NGeNk9qfqQov8BotAaXSF
U55s0C1ed5Sf+efRRwSgRVkk78W06t7I2FRIvzIZQxEIgK7yZTNsJJ8LprT4
/YpjxAVL+yyiy858gDqOD/S0xz1AAlxCDbPNe9SXS0aECVDzrAMv33pjxiAN
mFtOa636wSAlYL0O2hj2VZ/zS4zdzWEy4IiAtkz3W4S/MFde7TroT4ZRZSmM
hNW/+VDPaHVQoqkAaCYfMmqr6cLhi8YQu7qaaHqLjmHbJQnIJAOuBODvrjVB
MSLhRZpfkBXmzF3N2kiUwy+LpZk4ImfLGp3Y+W/Pz2ble7rJEYmBXOapTRHF
Ezx/TplLh0AXFTg1ojNn2kDTIBV0PStgqbnP/cn3u6GDqRt/xtHfvNEl5MvA
8yNFFblsvjAmX0ssO+t/4qNmzK2mKzNydrISJz2ZAPWFY2yEgaxk0J0WbIoh
rVmrmfc66kxZsypRn6qJNcAtV3mBvo1/8cjAkv30/agpY6eL9vxbmz3TtUpg
agfnkvVCXalIKKbj9WH4zctJwGz/r8TI2YkQLysWiCQJEfGgepczZEozrT8F
cJCtqdL4yUYQdp3oVT1cuClgN93Py6+qV550g7G9wpSYdwKOTF4PTeZnZo2s
xkwgNQH+awO3cviVJk/fGT7paCE7fkMrSDxEM9lx0Wv218x/Kw5R4GRdiAPm
52decxUxu9crlZ2BMWNUQ8I/CqsZw/nNX5CzvOmarm2Ms6o9wiX5LnHImTT5
0p9ZSuFMj2u4v94Yw/5em4Se6y+PnjnqTL0wp62v452//z3esHReN0B37rTy
DBtEX//SmJp/bAe8qF2pk7m/t6Mb5gYf4N7EB9akwL+ythdf2jaKa5j6hTeB
U9h1YaQ19hGtJlA9SxQBHm/EP4cEbgvx+DIn+LKf5rHhuUqbykdmLTgo2G51
LrkcQu7bg3lNM33f3wblYEdyw4p2ntYqiLx4+YrAiv4zXM+gIkyIBwpLVgjs
t6HYbHjZcmNMsjlzkGlBdPjbMQ6bzVvSUH+EVJQsjckfgsdXOUWkbRxMkjwu
FNBe2Rv01VMDwIK+APVqPJVSpJozbddWBrFouCNktDh0QisaqFnJl/iTLl8Q
rlK0Jk8sk7F5JCdjBmffdRFiKg6QuYb40TMbr4LnB4z71qdNfapzC/4tQYeD
9lAmMTKajCQKNsVcp7WgzLVGSUcLS7K/0uWg2AMl/BRzTV3msID++pP1GObn
q4kKbHQjTX4Se11PGLPqKw+z9njVAdo7aEpgTgbf9ek/v8HxggTIUP4dhLMO
ORbV4VJ7Tjy/fWf7z44unhRrOgYcfq4TcJ1tRAl3VlW/DSGWX8bgqnxcRWJy
Bg7HAYkHwl9kRaSB0MhbhgmK3HzXLiPCUMvoGFO8we3Fz5UooNFWzs2zMz85
W/0tVk4QLSYmy5Tz95p9fme6QkK3Pe+T4e6KgmstH6qrnWyZmDekuWuliT76
xDjuvPVVF2hmaCb2Rv6D3dtt3Ex2QnQ7Bm+YYJvDZ2RCuqZ4pLzXRmeCl5wW
Ja/cDg+bNK7SbRbYlr6zZHd2wHJWyxeVZcg3oEoxoCeQIs1fjwa2mfri/Ejl
ErTgkQORgCw2nTxH84kL4DLG6CX7D36oECoAeB60A2ntruuHi6lfhXaFSGkG
Gzl/EPNQrRlFmMJfbZve/ZYR0opse0dwv3Nw6dXdUq+70jK9fcwd1p9a3yiY
mBCm3eSpugpDD+OnuzwXL5p61PQ0hFp3Z6TGqhi0WEWcxhctyVxr9Gx0u75E
j4pDQ9ZvHMq52BmkOcPtYsX0PgT4f5xmEDIrloPWXEvB87nqaiPNs6vfsIpd
xZ4FEwegHdGTL+z0CRYWvcmUmXCUnFv7tIAuMrNdX4m/TDxDqcM67EU9dFPO
DHvhAY2X9Z87EUgNUQp5TEk+vrrv2+BAGJPKe40BO7O5U5hOyN1b1UsRtqpe
udyqablQ3fhxq4NTlz/LFXhEvhQJ8r7p5xYlMFcq/gHaKiT9UbrOcXL+mHzi
ZMusUCyMbwifoJEL0XVNj8S1flKo62e918RKlH77z72cqvNQNwmDVdkfIbBr
syg/+taQijuenENErE0adTv+dE9Uu0ZnSAQ3wxaGQe0/JNcYtEONJjgum//i
4NjRE5J0FFECRHkOkzFgrGS4DUIBqztRmMw/NJw9ini3+QLVEgLDKxcnmXX3
wWqhP1/bfyadhiWPbScRGjdt+DJVZ8nX2iZalV36BrKXei4UB4x8pM75ILUo
W5MpobKRzhFGfsSV0j4+8jxsengc+lb3XNaEPgrWZ4pE6ykZyiXxa9ZYaxWh
1n4dR997s8vqHqDH7VhL7VKDkGCLPiZ7Jh9OpFIKwb6oqWj1W4JdNwkp5dJw
pi8q5gL2wOY70nYZnirpT2Otw2/9EpB4xILlQufwmknamQIKalQtLt1G33JI
+epevlGc+xTP7YjlWyyfBdhkxTMzypnB+eAN9SA9iBuxU+pXK8AfTAk3ySAZ
vyulFQNXYjsygDWPoz8Ma01bQCAXa9NmLtHimB7Q+IunNvBn0kDgA2xR7h94
jQ+OhGiNzM/gzmZAsUz4rl7CzB1llvqvOJ8mP2bi8kECo+pwlQirZ0VYMkNO
u3uE6tirWfhq77xoYewcVTy1/wZxOJ52wT/CKFAsh8crPxRscWmc9rg+v7Lk
mqjs+a3rDos0nszFipc14tjRzMD0NeZrcV3zI92FoGBhI72YPY52BHsxaaWk
aIySzdG/c3CB9g4wJjYCgf55kOoPcfCBw+WG2jqhbkVnKdsCB4HAV9uBF0hn
TRzzPupYmzfPi1A2Mo+sS5F/uU25J/Ick9VoeIg+xBGq2DLEY+0MJOZNEQGi
/glPESIr5AMkDvwDCvGPqz4vWXYsPNeutJhhKY6jnpuFBl9v82H1GtHIih2T
vnYNbsEoStwVPu8ZepzSZ/y+KbSknR9s/8n2BvnV29++xaOsUKuFl54ai9rp
fpnkOxgHaRoJcZ9X6V7IqOTw/2Rkqe4kVyzPS48XkM9+CB4Pjnod5M8yq34b
xRAWTKF66R6QOysfzXUG1fsvJcjSTrlefUuqGRYvvtS2gV7LIWCAqIZ9xJu9
8DBhwHIdOJ1jdxOhkhYyK01/8BgNH0XqkbX/2Vbe4vuJ0kW+LfrkQ9k9UynD
CgxmKkKvuEQnxfVsZhaQ3bm/yRBCFDoE/EZTLEAcYPzZiiOoMr0YloPxFdQm
IXy5oB22Vby4Pybky4en5OzZ8KsB3A20TmSkOtBuMrt2qfGGU0oJNp3Q+o6z
In5vpj+/Kk7Hho21NRI7X1y+FGxIwB3HyDZALbD/WdW07APIrloazDK6gMyq
qpMcRUlQyqMlDgyNyZyqWqAs/7AmvzRjwQOLrSFtN2HnK1NLuToQ5lgrsr3D
lKAKOA0biwnp5E/Kw/4t+blT9iYlDZX317AMgFI77COtOiTP5H9qSFw/Okd4
Ff/BaI4AYtP1tTBlo09+U+c+VoLWet+0SFus1x2A6NbcLTiKsOXZOdDZRFvS
C0KPn9Eo2Bm/BDNO5a12YzWG+xNkDykGxM/zOysqDX26fEFWwnV6atvloOlK
6ISryUkdzj0lXnENN8VOtaG803DHVcz03J60G16jjpm2rbjB4NnajXo7/xt4
dkk/rfBpiB8SW+hOAKliCJ/9eHw2BeAOLRtwpTjga+FqAC+5x+mDGN5Mwu/0
7mJ9adylKmBp43sse8k912VmfZ3edR6DdSlfKbSGaGmmiWodMg2pkMYKQmlC
neVH/wqguA7en/2w8nsQbOusdOrkCv/MxTYy51jMTG4GwrzJoZqKGFWyMbXl
E7iYhIDE0aceKvGUzeLc3fw10TryVVfPwtS939Foj3UP0v1wnJfoDJ3sI8c5
/d7+AbTPTjhVW4wqjWOwKEtBIqP2WFuOlbDk3BHjfGzR89JwW2CmyzuA0Qgl
Ud8VMxDTj8G36PIPTbXqc3f9ljnJ3YlbUepSj74UB+Sn2xtGT54UDE2tLCV9
BUTgl8eWrZzs4kQ1kgzzVzsGNFWPpsWEmsc3gSVFxRkrFeYk/7ehBxuhWL+z
xtlobLjBPfN+oTlcOVbw1jg0C1YRM58jpLaf4bf2LrWxhphP2rYgjVbCnb5r
zPq+dhEpcl/fJcyJFqim1q8/rgakO5tNgcC5N49vA8kfrF3T1uEIA3QVfTf8
LZPxRxc+Z6HKIDyskUANAB0C9dCvyaun1BtHxZ2T2uxltkJFlqrREk6DAcdI
RoGkhI4gdVWrN3eyh4pOEy4srzwpAwNla8THNiZYpaBK3NQkmAPZa4MwqqXF
UWZIxJvkThq9dvCL+Yg5c1l/gxrOcqcQC8NzHRFRaa56XTXck+FrJzHRiQLQ
fKxzIJk68H03BiPdknrUpMnTffwUei7cUCd1+jjWNHFef9CqpLAtqulXduKw
SNU3cE3LBKXpa6NTROJ/fqoyejh/OdJVFt2glu5E6WTInt8zu25O/qYwAQKw
TTnJ6bdhyzthA28mAmCKD/RwzLr5badfLyCMWIVwtmr5OxvVqe0YS/qJzDaT
wHqaILJ88VKOvgJS3TewLVn+AapCpw7LPXW0vMDEIxtqifNcyaLiUuBcny0g
iA+09rkharxWvSb6wQXWolFQEBkyYYwBXfjr9b72QVilnuoGTHkpFFS9/e0A
XyRhDnCRB5ZAK/DoLo247uUn9jaFO9HAgDzQBLrLsIx011699WzvziaHKgTT
ihY4gPoQkQMgVj8cdJFKmpYGpSZhQMpiDKaz/lZdfETkvA4k28rmY8ztoJ2y
8zyWoL8fwdAIlap0OpYwLd2NCdZSVrcZe2VZ0DZ3GHf+8VyCmVdwvklz5oIy
2w5ugOn4B1AqGNaIS3tqFA3zaYFw3D4EeA6YEEDZgOyiXs/PA7ROyfdlUZEm
bAs7cNAWdMcXkGVaFIwQ83QgnYYhk0Ib+tRAcnXMXb+9Apq6i/mqEqJmRiPE
+BDa6W28QtXktifiuByPnNwWDvYfuXsVac9/fSjmO9RLwN7c+iXMiddxeV3e
xn3KMz9porNfcLFctxl7tiZJkF7UaQ7Q0z65TBDhkmW4+/uIhGBqEDIsGK31
MQki58zs80bZ2gXWrnYgmH9W9XCnkEfyHCDFbCyIEe9jZ+qj9LEY0l1dkvzM
O7OtkgjvDodZ3vmMpa5Sk1p5293gB1aKQIwfVmJEJv8cg9FkoFgA754uNot1
mToknq82HPdvpfdH0VLF+vVZn/arw+gHebXZWqgUL4PXHgMz5wephvBXFDzy
z9uMlcyVn5Gnw22Z/O5c9hLQiyT1hgJJIWW47hUpsW1kzm4U9QSZ/VXp2Hff
lXYLfjQ/eyYHpXCcQL/2NeQS01Y1xw39U45kr1Sw1T3mwIBA5XEx/tqmSB8l
DFSvwNzC9Ldkjm70sy2jfUK3HeCGJzwfYdVLkdodv8RLvSG6c9NnzUSsnruB
CTCBfZ8MnntEcmwhe9Cw+OxmoU/psHLQBLacecdLdrWAc7ueae9fymWoFk9O
i+GkuFCAfhbs4Mj4tCl0YYHo6ievU60kp3VvXBqPA/JqCk4auzI/4vyfsYlC
UhUrgTs2zggClMrq3GKMH9EizSIlo5Ryv088OQmrGjcJWRnATScuGovldrAx
QJ6wlxkY5JnzFS/lytIgftGY6ewyKUclVRipNX/5EqHtmzD5zLOC0+QsxjmW
txa9yj801Y4neV371YvyDM/PALnsHqhhXJPy6kMz0pYUI1i8wacvVKu7G9cE
/g==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfQrc4tgpUGx90IG0iFTlKG8JM+dMeKHD9QSxa+6FljhzMMJEoaZoW7PNYEY5ODn/l1GXNUNoymZO2uj2bsB3H6LtCYqRSz+nXuGEwVNXeJyaQDhiA0Q3mpRWRzvoN68+dq1ln0phIKJN+fMYOErirqONiN3GjL1hPe2YPTtmJNdXgfPTRajxNVpTkANXd+js+NWDWV6W1fpZd358f7pX2WC40+8FFCP/voNN7oS7tgp7poUE/IUbNPbMgLvjfFEbXxrgkl6C7Tt2Io7yqJX1u4HcKHg0LF+dy5uBs2MKKdnIOs9jDac5PDX0Sf3d/RORo+4AALB4R+cLVzG9ngO72+7xysuQqQ6iUneK1CV1pcRsmGb6nLlew2HrbZGJ7qFUUMVhCrAa5C0cJqvgsX1Q5Qyod7DcjgABsndAerrmVehcSuUS0E9YbSucuDZt226x/NoKh5nGJXjzkbn0n9hiUIeZIhD6yteQ5PLd77F77hTROBpAqHk49ZK5y8Mn+sYUo18dd3uNSz/KsH2nDmUezh32leeu6ocwZI4TTgkM2/P+uX3qwSoY3aMyJK4+2LY9S+y/wtZvasSJE7LFU/bV9p/hB3M433TqAnOITY6Q1hQ9YullcqtZtDxAUU875WFL8p7EptktLsk0ytNqUn4x+ovD4s4XE3Iv1CLPkp/EXrvAKCYCGVMFZG3St8sdliokMovYI5gf60tUQFS9LAuOyZxcCqSzRunSDDSbFVuBHvyNSA8Y7aLf3T8NT//5OuactO0vkibY/M+wXydq1WXRYNF"
`endif