//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
FyKyYwP2JdTtAcJXIXCIQop9neuMI8K3PuUOSf+aLduNIUgsTZUVb6W8i6od
YiWG+qA0LTZ8wnm75mYJ3GA2iu+ANPtB8H8g3cxKtMv6Zi9/yMkSB4RDrSQK
e0yyFURt5eF25u69KVNBw6sgDWXUbU8QJcdZN3WRo70SzJoectGhqOFrHwJx
gg8BXmSVr8+y1/YtSvnpMWHz3F1SOqEpKYMwCsjUmpFp8tOevD2hE258LO7F
he5plp06fMKBC/LVFCrMuHMiH0mpXHzqmiqCb9a69zqVUFtTExgTB70kT3R8
AYB7/rdWcg0SPiv1VzNP5PY9ocKSs3glJl/tNcKWiA==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
p1zuYIxrRj/Wfy37sOSK6jC7fv2FcNcLfEfYDUi3vtwoIDW0jULJN+WTeMKX
EBJOonTO7GlAHX8clCDWWtaolrpJYgFPgqPr5PH2aNdq1WBa7AFXbGx7nOBQ
2xVfnNqXEvMrg8WGFQ/9fT5IH6491dJAd7jXPrYzM10ia+CM8MBaB2k3uj77
/UMvaWMdclCzwlCpiTDuJl4q4YZ0NSwdKQU1yK2zaRTQ58245G3Osh/n2YQz
7O7MN0XjyRM6U+woLazDalFZYPtS6fxRfUiMyYFQ6IPI3qzel3gz1m+1iFZW
nM7pdMbviG5UzYe2Xnr++niCzgyOc2Vjsufr1SF0gw==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
hhKSfAdtKV2QudQ5m9S5eUgYoHiwwjSbRFfWluw9RM92WsUggY2lzuuQEebq
WwIaMV4kjGai3xoKyFRxt+Roj9OvZrg5Zp6EInDIRAz6ixPRGXBimPvsQ+N3
bkcVCFkJEWOhsuLhUaVmYjQH3Wq95HgvHZZ0fCyuGPGfg6D8TXufpnlAyPiq
7FDwTntameAa7gM7hezLuCJknKiD/jF63mWqc7FMm4HMV8PssnmzNlLMBSNS
vg/D8LQUvsos3Wy5ZXH9E9HrfkghtZOi6G/m5f/fKK1g4uC9vzVtNpPLu0IC
ixGcOqXkL+RZFcx0pBc/K1Vey2lb5M8dq1KkNqHDFA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
LUon98fuqHrwVhX3uIQKE1TYbCoyUCSG8Wa5KCYnWJdjFUQGibPcJgSqeCIK
h1We3KO8+MkmGGn8Ckt3v9ctfOxwgC0vxYFZSKOkHxp/Be4L5wGCEL4c+4hT
GH1iwMv0qB70ZKR512V90v+pCg0bkorZ0hGYusYG8fFWzQKIAwI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
AhLyqa/SzQ8rP8wQIYsFk6agSrBEyYNgfmNL0vGz2OyGRkEQQXghhkP8rs/X
C8e1kt3jvav+qP0Z647bbDiG2+A3iPahgzDeflPqqB3enuaOQ8z9BoypSBEy
P40mondM5HNbgjJkZzywNBcTBTANuozowWe35ciAUUI5P6OTSCnfW4e5xl4G
BsAIix/nqvvok/m6KZ0tgo0IsRpp0bEt2gWAMN5yYYtiK2tiPRZhBedepfPo
9OGyCnmi3OqaeegCU0uanJ6SzxTEs5afp+gS5llvauwStBBT0rLeDeBD7t4c
JGlPdOR+vPoDcG6JciNgn5D9YYUYm9j1UgVCS95YRU9GB9Ln8NushBGe7Ste
LrdGRWgGJRuGMjARDPJfZ6qXrBXXUQ2iEqyiFotFotb3/hwk6/UxIEXk+FV3
+Ze8vkmI84SMrFiPIybmxI/b5PJGtRy5OzGHCkhYcmQVVzS33jrMGE2ZwJN+
Jz9x9CbL4coQRutsx5sm17oFIlGLRPH9


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
CTBqFiRKwgPRQukfiFgvummS48zX/Fpe0S6fcMXhjaMiME6y1gcK4f5ZxCxb
w1tGem4JgMThw5bYK/85IfZg8iNKkITrAG8e9uAdCPluDyKADOS0hMNHwy76
1vs4EoGFFSKwkEsW3H0Av6z/YlpRjd8AiXFf4ZdW5zpgPPdV+9M=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
J/Bnu1Fhrj4aOAebwNGMTkjut30zZXEeeLVEnp6fOfKoRtrW4ZUuSUAm2juG
Dg2S5DsuVTpqiRXd9yVQ1J3mH43tJmqBE/PVDzqualZgviQqxmkmwDSLpaXT
/JYVxfUbfKWUh8ow0YWEXHL5U4Fz2Eksue82c3ZBEMaYPVMROls=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 95024)
`pragma protect data_block
gIfArOZtkDmnLhrSdb6y79wBPg/5dgXCjvYrUlMvnJ8bsVVtRJRlRdvbRS54
Lq5nO2xFscz5v6lWh2eHTb3Qx3wOVA/IQk74SXKFZ2KMDWpvlDc373/+c0yR
QwIQESkr2FXQT9QYFPwpR2MBQk4pMMOTy+gEFT+4DxZeD8DVICiEG0fPLIiI
X9B3rBYxB6zbXLz2lVzEkb14HlX8XpIzM5yDCSx1w04L7w7pr/nsx+G7K2uB
WZqbYTLCjpMTwVZmngG+vxFh7FvaEpBVDtkqeMgXT3BFxV8wRU2tmWvQYbTD
6+X8UyOLRlbeJ+gob3TRYeYdu+9giq/EncurEtAt/I7IsZs6T0V/4HbdpQPV
GI64H97q/NJoeWhhsTTlHlYBMAz8h5frmJsGC+kKZCuwQ4c9PWM1495Yizl4
YnoUtZdNhPPWJBOACynnPzWahjAPeF+lyhBVHnJwmJvoPXAbCpbZtvT2thd/
q3hP4CoaEI1Uq+QEJ+GX3JPdyRpj5ghg5o5rtqH2JRUD+NP1X6bFsbsWT65X
6Wr9yypPMYD+ZXina1decFYoQL4rQqIb6ILkz/cWpxWfVlofpEQZ1qy2oX2y
F/oVDRUw0EcDhWXqqIi/LrXf/21oJq2TgcaUfXQmlSw18iwhAadBRii08Uy6
FWY/nVWsrtmumfep2Vp0vRbwyz6leqw1nmulI/z9YdeZsjTGAhMp52N/hSKz
3TV3fG1JacV4RaoRJPpAnetp4hXXzbtfDpL2/j9jVrk4TC8ephXWfJtAFcfM
Cc8TMc2WSk0hpnK1oWTKf6emDgxZd2XJwHDSIC3aUHefroSh4n5piKsjkW79
EWQwnCUrHAABVxOV/RTnvhyFT8qYxzVnDho54T3BXAfsD12m4EKGWg/H1G/u
bdl7M+5RUCJ3yZR281DkhZVEuXZPtTEr9b/t500yTBqw28alm9ef4IVCRGpK
MrHlwWJSsHZeA1LIF6RgcvfrSXxVI0zIXkILgMjDG7w9lUmxpEtea7Ul0C5W
qyhjcDnvykxyM8KU72Fa0kDNvTlyvKnQt3JYTyBrkPSz7yHsjC51I+hv0mCB
9QBSV1lzNqmqFkmGcRWpqUEO/mgfPEtm3xwT7HW+yDSkkzR3+vNbXSiO37Ih
KeEvx7rzRPtkgLyukuWG8X/lxIRZAqRKQw/k7Xl3Iu+HC//J/u9N9m6fnA6W
KZdKPI2wvMCApoj/keOrJxNXW70iNO4wtz22ee1/Oe30Bb9COIWbf232LnKg
vNEUyJk+GnK4sKV+n31Ex5L8SQQDtchtyvLVaLN9wA77a4YiY27KLGkeKjbs
wmtwIqGFzVkZOj6PkdMFm23GUJ6oMsdaGKwym94ewwo87jo7ZKkX1wS0pIwK
mMSB8u+p66KCul5JjfwERA5HbTt3CXFDcRYBEZThEyA9ojkcyFE+7fS4HL3c
HAUT8i/8sGmo9lH4JaTEfhhWlqy2YCUfNDBxR9mhj3RBYQIIE94utgIcdLi5
RoQklnCw8NIBa+FQK3TNw1QEGjSwfDye/M+3chep0Wv7k/70iyye55kGXWg+
NDZP79XBDIS5Vmh8s4F6hbL2lW+rs85TjUnY+EWvPX1CeCdOF7d+gcbdbuMq
55r6CXLBxUk/hTkJa8qTIovTuSK3+VmHSBvIBQbJ5nxC3t3sd2G6cfnsH0A/
PcaBt9My/81spUNClGllcHh4HNrGcxOOf40F6GzIM8zEszoFj8Uc/vXkFlcV
cwPeooUf3WteJL0S1UdH2TvpKUEBFMkAMcMTDJ7VqY3I0KRvjhNBjDykHyOi
mSuyfr/7cIhZ/9JjxPee5Uy+zvD+m6ucRxOPQp9KflYRK7UOW2C555y8aCEJ
d9yBnCPuqNxqZ1xPStfSUbcd5g4Zp3dVUz61LIjL9NudSqGzGnQlK3k/9rvx
Vn97bAXvwLgAKV/dU2eK2VjdNPAtD+g6md0vj/+fBxwJu9hNIiiAqQQ3y+Hi
GhO/uo+TufL7B7FC6LxeqQWai1TfDQ08rs4TYUy3jjYP0RSDohLPzSmfG+oC
NSj4OSDZpoATVGkQ7FJWly5+EmzKqa4kEOwgG9kyfAbXxk5NgwjHFCXMKjOb
c7cP41/NfF7KoDF4Ff+3kctfuYVdV8I+d4V2Zd+OY8qn6PVDU3hlNygYahZO
K/TWaX0doR10Ofq7KeUXZrAGaj4Gc81JIePZih/HFyvJyJaAIFv5ZR5n+M1I
2YG0FM+WUQVzQCZ2mOc6qTpxAqrRbtsHI413FjJpDbh0SCEVjwnnaPOB0kJF
4/zrDfCBfVXTkeeeSWl8NmL/Xar/gPnYH5JcDC0+oba/IgNVcoxLx8+9Sn4G
kwPhN6GniGmgfe8/opj8640gPUoxpAcI8CEqvBRxHV45GSqG9T14ixYsO5eO
NuX0wamn4WRzYFGQPfAOCm9tAzrw0weM59+211WsvpW3sIY+zHUpvdUhyFWx
d5kMFCCsIMZywPRZrfvySXhpQ7T97MLY2EP4HtWxEkIprcTxgR3PgY5rR/DG
2bnoi55OHMdHf8enQS9vGLQsn47gKEw9r8SAz6L3RjMi9CEBHH6vWHmKR73e
3QJvyeeEKmijm+O5b308l/qT7GWCI8zqxrutQ1olYcFk6n2akxMAnAkpd62a
sIjgQsjUZ+kM7RfdRWqqrWtZORFLbfMG6SmHc5U8tAsNelJ9RF5PshgzjAaZ
TCu0Vk93HMjdvpGNm+zB6izywbS1n8n0N8dP3FhV8SqPspVHezh9XKpIgUbb
Yid9q1fpk/ySMswH22H/OuBJH3i7MMZ2X3QP5lB3fkBa+PPjmXRpS62iANwy
aII6xWzrAFN+7mJG9S4JFHMwbDgTiOc9pxAmiV9SAkpuxLPFADeaGuQJM+0D
CRz9yJ/Rxd8f4AgilO/n2TOkVq5stgjUaAwHkv3Ogf3fDBm8NoiYi8vTXYhE
oHMRoBeMUsZDWgiOGstdGaQy1gKYAzu/wabZvenywiuue9IfX5K9wszco5aK
8F/irAkhUskYkZ0LRT8zK8iHhABvAm7PpyWppZM22/GhzYrKatHgF5ZO1Bfr
k+uciLxEU2g/oWcAcX6Uq/iKL3QsPIAc9sdjpGwFCsqq0Ppull+doGkPxcyL
NImw7w2M83qxB8x0HlKEx3cVWDJ6/uL21AtMi6AEcrd1CRdxwsop3sV7eamY
v7TOuMdBNtOtMCUnyYnAe+k9rIig2+R6bkiThd4P293bGj6MTlq3edxd+tuc
HMOiYSEOon07RcSlZFbeusGGBEcccy8+N/nXwkZOOrWnokg7/WbYKJwFQrx/
6+jca60tbhDTBK1aPE5wu43SSqjKd93F4FdFODG+BI8irqDy3/QkobHjJbPn
CzFkwiPYHwFuKTkmVIxreRZ1tEqUh8/ikGEBDqYl5qSZs8LP0bBNrnjzSEIX
Gc7RTsX66b7sGwYakq1H6KpcXAjN0IRsrVOqW11k+3vPL1sa04RMrHXHG3DS
JSAUkZl8GZlf5GrL5D7VgD/5qzUQWuITT/hW/uvBVYtNIrNZoi+4FHIyVixK
luzggLOE4HdJMaInp3VnclriJ+tH/8vLve7jdCabRRXfJxjX37s7tMI6C50S
uR0WJtXR9FZzYryBlLBnzP7hVcUR1UHzh7IfI8Z4/nvHD1GoAZmG8rDm0r77
uzN7CtzwXtfagtLhIVTa9gLyiSyaQkesh1Nz51OwFoKrwSgTqy/M5KLr/1GE
dEvfSWho+MijgenWlCu1zLPiHEjMOXHresHNSrS+Fc7bbjEreFvZw5Z4pxE1
fEAXMfWTcc0WZ31nCfn7FpA4V8lQhsi2uXQvp3kKG8io5AQy6JdOnpDTXnb7
QNQdMPIw2Hyo41buU7BXPd2MUxORNyWYyw2dAXz+g5IjPvH8fFm4Dqr/JdEb
IirjpZq1QqWM1lOzmbnYGx/mlONhjzfoi4FqYf5PUfuSZQk1wm0zKlYrNiTK
5B53m2nv2YDFwpAG8XNFO/0lef2bHm69zppCQMSi8FvIsHvMSh0gfnIYAxB2
WjeIlWV3VzzOSPx/m8T9DwkrYa2iaAFec6w6V2ECQI+AnV1RQGLc2LkPAXvC
LG9dwSmYljEmcVXzdi10sUuMK2vLkzuCd6yDcyqj9XsErwM2iYaClt4c0Vxg
NwCJJMB6shVyrw9BE3SWz+M/fAaazJgqcMk4GNZnQ0n8psWZwAcHTCLByLY+
TaY7okjHS/oo3cH4TpeDF+ov3I922Y5Bfqi495Jkn3iMQ+hFHWl/7FC0CCYn
SIfdjyZf4Hi1tN5hOxXL1Quuhv2chrWg/sY6A4fcberKZkxxxa3QUEVMpfFT
jELfunsYuum1PCFu91IY9pcr49Z5SxZdQ7zDvztsNJkZmVIfFJ16EMdvZd0D
lPCHeBSXV9m5Sj6cz+RveFxFmBYj6YPGMrSkoUvSyCi2FLfk08f6zJwI2gtN
dWeJOziT3PEKmt07gOEPTTq68+zVDX/Eq+2cAfHU1Wd54LuoQbgbikRtFfZj
TPMd3OpCK95urcad8FlPDW3RTbtoSCOYU2wxGQ9WoyjCYpkzk75rX7fQ2lBn
lPXwG8ewmuy/5hcoTXemWvlyzq+BViPpcUC+BzEc+9i/25ua3feQTzPPDR8d
nFXc6RF/hLZOJErjJH5ZSksS1IHkoDVSKgtsfJG7eXNcdruLP0akjHAYDkh2
qOsRAF2kAx1ySSS5+CjZEPlD0KlNc4FECP8xUwCz5F20MCUv6WqivK4/jlew
QRheXZTLQJ5C9+pCYzNZH+lphB8Da8lp0LdA9ehQJuV8GlVoOIsRCFI9hLwJ
0i3mybYLh8HB/LuCuAcDGej4kLc5F3Dwa4uk/lqM6vliKRRvCFkalGvNKXQp
YsKmHOfQcoOgta5G6yuCaK/RZ0uAr94lFIbOaPpVV6FuoDNPwGFvYwWIMVxj
LRiUNGWa3rJaZ/zINN9+b7R7TEG4UPgR38tBS+r9qCX9keOXYjPuep9dvVJI
xBzHEp7etvMtEUEkvHDXZDYFAuPVb24J8s2FnO2OXGtgTKM+pg9QGxCQ+Gsb
2m0LfGR0PAmuzRYkZKSaJ4U95LjBI+9Q0Xt2id/N6J5VSrKSJdVsz8jyHOa1
zF4yo7FRPOJ6JQDXCIlCaoIjn/VFeuPih3kx19w/Va8I6yVNf1YFEHHuiqVe
lbcHHOp1hOd3Jwujd2vOEIWJxKDChc/csPbTIEe2/uqiM6M7v6kVw4SvP+cW
xvIWtafbBWr9xRM48nQcvEtQTV/tjA3cFf2P9/qVaR8GO3+34elBdKWcszwi
9qlPNPQOHNOugOU+vCFbRuw/1da2QeNAEuLjVIgPaBktJanOFUmqG4X92jcc
wXDVcZiJW9SrNtgZn66aa39jHEr7mqxCfE9aKG1uRirEVZ5U999P5Fs/qI/i
aw7NrqDXhRHQLymjsKrucuoUtbVgQSWfK9eCtHChN55PU4mFvuWYAhZXCENL
YcIIGdeTVv6v5HxBIEpQllGiHCWTkxwTio8Jd3s1OHGI0o/laVGkL5JU2Pz7
isi1XBMeZ/32iCwmoaE4RqvTlVvetUxISA88V0h9b/0YU4eILcHJqG3jV58x
0eoa/MEjBj7PDmDrbQtOozSEqViFCYqsdmQ2LWqUD5WgwlaFN5Asx8AQ6CHq
5EE4Wuw33gXbsRa8Hx5Cy1yPBUHHHcUPkd90QM6FXzld6YxKCNgX9y0OCnKG
wxKzhoHrTXmrg0v5D4ALkzTf3pE4kUasyf4uxRTc1rXB0jNfr7rXTg8sv8pc
xWtWtFM1AbuUnfc91gLPacGk65ayT2mMYSArcnxmiRY3bgzsmXPlAkxvzL3U
v/0cVVHzVQT/1qC8E/fu9SQ4lb4SooTg7DGczRU5dzpI0TItrxrZWhAMLAqS
I0/ajMoOPubIRqftN0O+UWDNF9xTQWOSLlDyGUJcZvzL5UfQcTE48fxd/sAM
JCFFn7LFil05AyrcGHlyOtANyITGFml6QcfjzRCHF7ziJ6O7blY7R/F6lljD
JMu+kZXYYkTUZfsYBmmxYY7FyyBqHES/iIAXBDYNc7fbOj9cMRqddW52p9mG
zrtqmhS3VY/xkIf6Mr4ycxzhT6G//Ug7RVedTEIUN9ZJZkHhJDUp0gYHbq9n
ontalkk09Lf6DuRXRPp95GAEBjzfvYFDFV/rOrIKGNIz/IDp4C7AeNYMN1nb
qSdWfpeV7h6/BcegsDNi7N9TZTQ2+OQp5QNURey295Um44uYtjk0RCfD2k6a
/CfiuMqn1r2lzZfYZE6H7D1GeppwCv1RC7EHMyHmHEVArbZc6Uq54pcfbqxa
POI9n6Vu193gXqd+O/Up77dYXhU26WCJ0s77HvaT4GbCNi25kYkTdb9ZVec0
e1s3ItUzGOlqAH1fmNjkQPeaKwa2MqJBVzMMGn2HEQeX+Top+lz2WgHu2I4l
gwB8JjBwW0Yj9pnHEMgk99FyNX1kcYIaAdrD+jMn21IPjOLIJ04fENEAHVgk
2G8ch92t/NIIQoAkiQe6j0BcedU3E8nczhN5uHh7BHXGHMogQ2KFa4oHw8Lo
ZLlJn8DZpphsUhbxx1QFjAsvUnY95nB7bGNwVD6BhyFd3yP/zXJbrMxAuJqM
hDFlocwTxaRy2bApBbP4Rv8mlfbHE7PfZ7xfu267Eot0sZ5dIOQ49i0z8y/l
hCF83FJ0eaZIIc0n+0imKnR8ETiB636UPjk3UpCa13RlcHN232J3N3y66Ig/
EqcW4X0OE/zWzFteI2WDuOHJj05XRwPgUx2T8Bocq8j8phEW4UjBWbvcLnmd
avLh0NRD2BvNKfnTwu6sINXrS6OZpBVps57458mfhsnBiRYBYTeYgfRkXtDv
zp+jMtmielBZ7U9CmVckhnpAtvTGHSQBDzcIjaIFJY7pitxG2BXsFLGeDZKi
ordHlNo0uSqUqtK8WnOUPRiRniZL7DydJ+XRBLN/xjHqsUc4Nxpa9DavgGcN
yY9Jl9SEtv8zElVareC7COycbasaEArYC+PmTsjxvZ3SJIv3wZnxAzfASCvA
r/wu269UecixVBEgEux6jgHjACxn4tzRB0Dzpx9PZz9iMPnIf1Vaz8QnaOgM
BV9P3f2H0rdj+P5bNQarG+74f4oIt6cfvmE93XbWthEKA1AfJavndD5GvRSV
/Rv1dk2lGy6BGKd58uzy4g5D8gVAAOGNIfAAJnQgPnbAvUBFDusXPjgz7LX5
GmAPxNfzXptXyAsj3X09/E9HIw7hjllSnPedsoeY7ki+qMV8UYXbGeRYu2rU
gJHCQu79pmk2VlvmCtRfK+pjAY2I0Vzny3PUiSwtVfYLmZE68V+YM+ubZ2p1
we1Y7lcZaIqk4fiJ5C++hKg42oakvE9qcOjcTktQt8KdFmZSKmynC8CmTIvK
4A05lGz+K3pdV2Atk3Tsu3ezmnkwlaWRqmG5e1ftrNN1KcSlh2dGC5KoneDw
55GTmcPDzjHYszCuvuritRDj9Zzrw9EpvoCFhfdMnqGcLPrTBfAfc2i8VWjb
Kh1hSYE4MBJOqAJKYKyGuhHyx6taAcisWsL1js5cG9V0mzK6aRcSimY1Kbyd
mw3MSz2JnLFN2EI4F71BO+HeJRnDg7KZD5o55rheKc2WIN4skbuTMIEUTYT/
KeHgqwFF+7fn8Ks+qAdOh3nHinwmbJ7TwcDIJ/6L72X+kw9Zc+ngIfAMGZiQ
KzJBneM4Xr+DHAMsPAwS9cjizWYLwqIamFvSDFF2HONodri0NdM+Yb5wkTdT
uGrv8IZVT0i7DJ1/iHu9qbqaAEkE5OyphSu8/OE/vXr/7pMmJLAd9AoCyl3b
/OfkOR05WrzOVmMn0wNTS/7UOyxprtY+1tolEyeD+fj+jIaUT9LWI4JwqqGq
tCfE/L2CgnF3PAsjBifR2QeznIqiEReFHlrKvr3WJ2Nik8H2OWIXeiW0yE+g
xUVNyLnK+ddT8icokmzEzqL8r9TkQ5YzcwmuCfIDCEsPvSucoIUogl/uWbkS
JrBcE0gMhKx4GSyzrJz8IcxVKW6JO0M0XApGmHrS6Zz6+AI+PP+5fKnHmHnW
yuudxPDD2/fKgSSHNqfvjvtI5wgwymkxz4htjmWGv/J0R6fEc6P4V+hNuI4h
1zGYU9ZTVaXQ8tKkQBfm4wG0eUtCF+BkM5D82z4vH5PP5K3h2tcJAiM0XwsR
YJCDKqXyVtQIKzBKY/bmUS+hWOB1k2YOTvmVXdIKsR9Db1qvOw5rGYJ8S22y
DRstKWZZ6A3NB8CQSbfjrfMj70/cnS5b6E1Pbov1+VSvrgBG/ya6ILGhTAZ7
HjXwdCv9pMFyBlACQ5LNbfiHYB4oes+OsuIgq0yac6w16DX3hPVu+NfbfWcs
UchECBaOiMLI3oX9jTN+LsLlD75Kc/j8g6JWxkSyigb8UIFJZQPb9Xr2kP7n
MVxrV2EbRJdT44JDX7n2wHHvuWV+ukY9YvMUTxUWwyjPEvSHQYdtUlR7pZao
lTj+IwYfSdBq6MbsU3aW0Y9SvLNy7zdq6Y32lHVmSqVssutG+qa857N0Rxd0
Hr6iddJrHH+D3dEqdDvKP2O5JLYbSvBSH8q+HOQvmt7txXbYZXqZ9A1JPG09
UlLCJ+WxYORtzDZS7u1XmJhbAECQ+r8FgSLnI4Q4cHkAOKvzKwspfFyx5cCU
mi+CWmCmCcNB7RDpnRCvNvVKxydgzgYWMf24Q7ZeP7K3zg43OwvCphQfeKD1
6OjZwPMyz6ZDkN4SFstLNikCeLUEXNwZp8d8ROYs9/z2LA4sfn6wrxB0gLRo
VMvrII9akuf+UhMve+RGj1TvOcqziEy3A9htIOg5UQqZ4vFyzvfZMk/5Q2Rb
oNmtOTNj6j5Dd5aTuo/AlgLZL0WtV3tfSLhD4U4pHxw0OEPKSDLYNNbHRl8d
BC6jcIjoHkNo1wrFWuG+q0XWe2xFOCfPUAktIHGu23dbS0foCeBjpPI5xECJ
/PVwJ6OU65EICen5LvjTJPQja3tiv5t2pw/zQzcYXQLfv1kh5ySQ4unkJZqK
OEBk6JZv+vL10nEqdRX+MD4fV6zku41cfVK5HlYcVyHKEJGKgh9p2xVyUA82
3XDw8TAUmJlhOPPfEy77+lTUu28ucSCBWz3ITUwx6NqLx/ayiD0ZkLq3MDvv
5Xl85BKOO6k72ARiDW4BeJo/eGrSVIcyS+RJqoJbhdYgHIok7p1yNWA2spaO
OH9hHnGK5nMYCtO2fmFhPhLqerElfStcyuuYiABB4gcC12OkmI5QsJKbSr1e
nU+O0nslNSv7q/r5nvQhrk33h7rQR7lLx/H5gvYrFoWIxfBdaXYI+QKzhx7g
dNVOBTTAxvJOjVrNuNIYspwqLo36mn2bY9B/fx/BWnFj8GE7r7BkTE4qsoy9
xzXjZu6IRbqJ+HuKprL2Fv410IPpUShvL4/XBaLd22NABxF/C0/SzIWmWmYf
p9N+0Vpt8hSj7EKC2d6+7sSIPAcnB2NnZzk9I/COu2UtOb3RvbB9kTnJYtdA
648HpVvkACnAgLCwB37Z+dzeo/8X8zMEYK7meJh4+SiR90z/F2K/EiMbqQp9
gI6+GuIvzPBENgBCEgNr/NUH4uVRKB8go+zOPFvlr5FbsWJE3SYpYrNlioiY
gC2FjlCfHwclyWXwexORsK9MHKlJjLA0HU4JN6dymVrEbNysnNFUHsR+/hb+
H3+Hy2CcADkrTdT11RcioQ2cqAw/OYEplmcgf+Kq8SoNQaYpRwRMnDAcl3Xk
duqwrMPN0ZlOMBIfD1kxR/r3M/W1UoK+8YRW7tPP9fUHk4SZ/PrDxbaTG8AV
uZrsPEIFqkp9MM6Ae2FDuttnaYl7BZl8NTRw5dMbpy3S7J9TTMmw23ZbNkpT
lxskPkZBMlXovwjhVDa3bIluBFYmbM/n9Kv91hFY4bufAdK1KQcRwZT5SLfs
e7myrgZl8uL3NWsUEwN0CAvjIWSHUi+Nvs74DWcDiWaxvM5U/5BvZz8Zj9S/
ZrJ1fBNk5B7lmXPNj+3aNz9g9EoR77ZbO2LJsQG5F8eDUQqKvGsx+1cYs2Ol
9bIN0frVHSzq/kAqljSShCoSZjsxOr3kE9mPzbdwJC5y98Ej+xFs9C9rMx7p
QH7Ng826TxvUTUByxtZfwa6zZS62Bcj2SunZ6uW1u3Dn8fmx3KSz8qSkqDLe
JapAgpnKhM/D+GViWBX2hGlxOmHl+RAad9JSCc1HUqvubf7RKWmdGR7MhkQ3
J/uJxhtAIZa+cRXOcya/z73DrgqvRAo+/xIMLwZZq1ZYg9bv3UPca3jwcIeg
/9hgS7e01CNhU1Zd/cuoBsd9WalYoqAJJhLiEe+SFD/Mgfu4T4az6rftEmsE
Gi3iZ3OQIHy5EOaMBYvqMvMG+GVKuK7FrL/9MtRx29iRvg4q3myq/rBgNOAz
926UC8lIKxRnit7lVKhBgAer4ZhwwmtrZ2r/WBbcwb+GtqZydMcYku/Xkz9c
97cw231iuK30b/ozf1ufEnfZZEiNofQ/o4FEStfyOP+SW3N9P3C3dvwPd891
LsWgRLtIcvbN7pG2xm1fJZztI1VQPo70VyU/X+k/lWFiTIA993dj/QZxNyMY
Cm50pxuxncsCblPUjPajrH9NZ6TgSnvdW9q9e2eSbpWsX8xq3kQJvu1BZVW9
sHAUN3OGqtBeKDWr56F9W/lOigGU8SDgA7JyQiiGrGKlMyxsFOxJr/x61LZB
VlVaz6U9GVU3fYuDYW1qMksp0DAoi3c1zKhNk0EDyEEnHh2TpqhZrqbd4ddx
EQN8KPp5x3y29fMkwfwE6c2APoqc0tqccEOcYi5USZ7YQvdhv/yptr7f9g/s
Xgk01jWU/rnDPhNVBZUYrLtVvcQkXS2/Rc4okGhClbK1TrFEirRRGZTUw4Ml
LJa6SCFiw4WXapDxNauEhQtQVV2oIIfm/DbCRSSwTUvYfHea/mv/5AOmqZru
2nnPGYpdTuOudTOMeo/UqExLJ/tAG6B62hiPzGI08SyJn6FDemFB19hki4x3
u4pWIkeMC7mT1059W3iJqfyE4k+WeNM40Qyd8HV41/uWOzjYUoJRd9VNLM3n
ah7+GDb7t0BZN23EFzSQubRMG1MhpF/zG/RyJ0D8GEOhTr+noTbvfJqzv5ou
//Dm2L+hnYNt2mv/thf8OcmwRDTr6JkvLrLP3vDsT9hfoI+UtVU77x46qVJg
K0Fq/sG/U9tz2UsvemsGc6EQJwR4M7z0goC4PQFhBP5BELhqGxWeVMjmQe2L
N75iSHZ1KtYD67dLBKG8nfjBxk1OHduPzmTatyoDngZlHYyPL5IxScZJ+6L2
mkePZxnYmHrqzndKFsKu027XYSAKk0uHg1Jb0Qpjtm8CQLmRdX6KNC7q/TWi
LIxr58qZMxLnMcQ6ILbDux9RcXK5SXli/iQK5xpYyvaFIAMtLUAJoetl+/AG
l7/NQ9mGcylGVQVvZCN/jJgBb7dkXBZZSyFrUjiim298VJBN7kVGDmbRsNCf
3bMzVE2KAKWkk2Xln+ggTgIEe6estBWzk2cXKs/VL7jNcSrB7IE9XQQxX7Rs
qRZh4Ilm0w5kjb6SkDH8ISenmt0HVEAODp2wtjVHQirJ+b5l73qiJ/34bOEc
83Uk9CL3rZ1mdEbZVv+VwdFph8w4HvMDGEfEMV50E32PtdWX0v7fOqpkAwK9
UJJwnGA7eTjW9WeAHn0Gv6q1CF/b6aS/HJjJy89+ZJ/Dk9iYGUwTf93xVq0f
RpZBdYJRsYPsokdKdktZUMWGT5mZ8iIQ3JrU04Ejf66IKwnjHoeNtB4452Le
PLa0AX8CEPuGiFmYE8ky9mF6cdQhf8j64otEGY+5hIIt0AHYnQXyu7rjN7d5
ux7L/LHmHIDyWoB4+NPPKIrROYyayAEd+xccgJ97vR9bcKtbsQxQ0BzAE8OL
+E9Q1SUMobo1HqzCVFBlMGO+lYJTYrhaSM+1z4tq8iOiEgbh72ipsQkV7gTM
66SMuXG3BegWFnSNcoDGGXMKa8up4IEKjN3dMQJ8GjTlyRt8j4i0e5Rcb9MZ
ROWTBBoy3RCzRKF5pFW1ltJgh0B0wfYC2GwAalKWzQrY/jcy5tb+3RY5Lqr5
fg5YtL2UcQkttMlKvZ5W7D5t0cBFDMg/OI/IsGirdbU3JBFMweyN0/XCyFcr
GL7HZ4oPd1DLvZpvz+xYCupHzFCOMnb2YRQNWSyteOIv7JzeEP517Q3+jmqJ
P6b6gLHnAUAneewQUGJi8XA+20Xv71/nrjnIT1ARjp+HvOknkzrJlm7avgU5
7Fq1UhKSsMzq18rEdCy/WlC8n+5L36nJhJjx8FbsqmLzh8clpqqmF050CL1T
5+fFCPLUr4UEP/g1NKNpogzuhaun9xnrwi8qrgIZ8EyfGjk5+0oL8n/mQy5l
MZVnBm+282zvyJZ+8ztE8qX9BxQNGeQeExU+yc5JT71RAqyWglejymZyYZcX
B8ZzdLZfZLLd4osQb3z3WZrrt9KtH6u9TTzbRzDJvz+DGlzk+FEG0Hzx8Y2K
aaFoL9NQHER1h2BnYMjzyfLZD0hW1WPZ9eQfZDEj/zdhgxdLAXh9lZDRWjnV
NNiVP9hdfGyG2mS+G1/NCGcEFiQu4xt6pPPQX7PJuYVPvRbJJ/JgTUYPlnJr
XFHk3rIdbSt4ffOgoryCATfhWbuBmiO07KG96Qtjw5xOfz1UR+T/ooQGm1/f
3Sngl77j273QSvduXa9GksYAcgmeT0vFAcmKJyF2vKYGryKr3s5ENRWL7RSu
0fpXBNslb3GOUPmS1TH1Jhrscj8kxV8zWtkIExF5wp2OULqmEB8IKzhvpyBz
Pu+EGFrtG94cBh1NfJAu4Djb0XOyfPKnU2zk0zXPmF2Kj5q1NfQ4e0Yfv9o+
EgibQeGV19wmfVWxQBspHWNvJTvEkxI5npD4DN0vNN6CncXnAjK3Ike9y/Ii
pTi/CcBIQd1hCFOaagNK9ogRuH6jJ0WRUlc+h3CwOTtG5MINFG0tk59AY1J9
JZAVkRQuusc+KWkU9itygipeupY583elAjBE/SA1rfRuNrGZdUM7s9Iwwm2Y
HvlTalC6aHnrdf3r9JdLkdcNl13sN66rwo66FmDGVtNm5QSObxY0F0XtqXmt
/pKn8PNOxc1dkVl1CIOhelYSHHoHRs366zmfPutACex187uUQToAOUVwwSDN
PR3ojJuIMISyHMTYZfF0AqDS15gWrFBAP87+mp7tC2sX3PtZ99L+Z+oXgU+1
/DncxPlecDBKwCv6NRljm76D+gxy+pcqRUe6fRLMIKfhAbw47X3rmR0t69dA
3wgRr7Xxv3tO2btnL0ZIsRiEr93QIYOLKgku6g4A+cHZRc8jqIUdAYk82Ax0
eBm2J9YsvqBfQBUmkoic9CmWzSeCZ6UA/P7JtO5Eyle/L8EVlEzd97TPcG2W
973w5kbAe8g1KaD9zUz0PvM4EzfQV3J7z7l7g9MI6/4NazrlYKpRXiEq5cm2
3EnCIfZSStSLUs8UP3TYQWJ1RCuJwtkzOk3zGP49gyjhW5RT3nGJauhlDXAC
ApFElwygxwIlW4NGZX7jRwmuyJPyDK40eNHZtX5R/2B3t9sOhdC2EDyPJ7vQ
IKZ156bZiDZmpJ+kNH6kniPSu++cp0Rc5V2TYwAYnxd5fpL78nVYJBiO+zhm
w8p0pHE6HW6UWbRgMA/7nekjvGWUA1K5C8RyZCDYfev5e2uW0z294v8kdUIQ
h/k7q2cbv7MIEmwfsrZiM5cMOIXDLJbc0FtLYgPb6Xyi/uM299ZKdtKMXGyJ
GFZaLZ58Xt3UHwy0ZWPjS7DgvmAUFx8pNFDpie/DURefH0WXnMYPUd0wnVgO
5nAFPz9VG5BCWhcd8j7pUOC3wVqmw1uNNmqFbTJehmELJurcTZ+U8vBOAhZe
EGfrR8wPdyPa3My7Nzvj+xMVZzS+xliIpVI72nfOivOd1w26fKwIU6yhToFy
iOJM00VhPUYj2tEJkL7cFjzl92oNgo7BpGcL0KvnUDDKtDs0JPwY2l5XXldc
FkAPnj3b2qZzLJJuq5nDchBc7vOuxwqGDDbDBHC8oelltANAz8WmfQz1CD1v
42j2wrHj5AANyWZ8qvagUdNZcbHLuivnTTzYgH/PSOXGxxmjl5QwEeoaC+2D
cWEp4Axx6e0xlcP65h9a9NgMZgLQth/tAyUsrRi/9MW8M2qOn6UCijiTD+sU
4qqdOZnuXUfALSQXicUIGXLIGDn9qHoCMaxpWgw9TBih7smmw8V7MMYzay/N
Ziy6ohwpTFzSVDsWnVZa2MqNxEJk/uuoFkWeNdlzUZomMmx6HiCqLgnDUyhM
Tc3BhrIC/foVCe/xXKM51bTMy6U+Hrqk/vDUz2ES/blytCSxlv+NIQK3m6gW
VzEs3isby2HmPqw1xtdEd1/4oSKoqVYisvLOzvG6Y+uVVXfhDGt75JT1uKcx
9q8U2qS3OFqQ2hFqWygkASZWEd0eT6xjrJYxCsc+BOV3ZxKEGtLm14BbBmO+
OtQ4SxgqnwPIl/SmH00ypY9jVYowV7OyS+LmwastFDvPhhJQ2jiZ0Nm/vtkg
qeJNu+TBQxEQXh5bxei75DW+/c1LJximmq0omr1YmScSn3vKk2rV82L1lW0M
FtlNIw7i7TqrkFKAM1LNORriB5s5ZX2ubsQjNlsJf3pqwwAtq6qxr/dmS7xM
EZU+X4wDQdFcZnhdZaRi9NTzlXisIH4viZDxstz5bmTgLT3L9ijv93WSTmFY
qn2gYwtp2xJ/76FmJPLSZLmZpY56L4cgJfX0n08cggK1q/sQHnIWo3j1pbDV
WEJ1ULUKs75shoaBu/AfXoPsr6E8YofCS5lNME3LshUy44X+w/h/2M0uIs2M
HE5Y1OCMyOeV220U5KaK7i5ZKj6RYH6M0WOfiQvsJrlCwy5mSLUG+KDzPCJO
ubh64hvghODxJWxWfvvTnLjZhajFnTqUJn+5MtyTOZy9IeFTYBKp7duRZWLM
4uM6lj4PNSMzwZ5OucLKIfvkk2sr3OoBkwvSlQj7X0py9kcQXY7Z3BMR19Vb
ZLk6EZ9yr4mFq8MNkvcZLFHFA1mCzNgxPPZmaaFJ90sAC1jrgEHrd49hN6Yb
1A/aLEsJr4vpw2YGd50T7O3YDRpxiV2aBMxO171T47Uq6j1Ln4bEzwg4Lbe2
N+MoNjxqP72ySuDmMwpL7xI95LtSQJJa/z25xJ09fCibT+mLlTzPFVr3Zncx
VSfWd7WuGXtpEgriLzaLQi4QMvRQ6OZ5xD47wLOSqLDRfJrocMP9lEPLlDlT
zBX+OQt02ho+IUJxLmGR6625amc+RyKv5SP3M3vR1y+26YRIC3Bt2FLV8rJJ
fXhKIVuJ330x/pjmMNvnRn94o+gWpry9Zsq5lCxjEiw7L3QWLHtMa8s4duYG
5VoZ7Fq49bXssRlIqR081tHpcA4/Ew9v+mVrKECGQ1WhEf1X3rCk6/j5IOG7
RSFbvOu+6Fes2cwzofBCAABYG39U+vJtrTeQJq/5of3XUmg2v89ux4aNRxZW
pqsEEPF4SPl8FbraZN0KM4u/3uZvGd5Z1vDe3LED2RIHMP7eQu4ez0VXXwGe
lhxChtnd+tjknU4THppvEAOWOgtbNFRzUYxuE+/cWlSYON79y5AJp63L0r7m
Of8wcRFt3sMSDSRkfRTiSSoC08Fm6gGDabzYv0kCkS0h89N/GwwerkYQChgu
hzkZiGyXQe6ljDoC7yfhPtzIR61n+3mxfrlr+21ENNfvDfjpQijsLphYv+OA
1I/4fR6LSF9+DWIuu2krMNutPFL152xexUiFwsw9xIxU7WKAerwO4UUclxfi
FE9FOwme++/BQI8CVrXCD8mbVW9Fy209Gb8vpXfCcDj5rboIG4DX7gL9aJ3V
izqu9ceOZ3/bbHkoX7dil188m50ZhkcrVOOn3xu0cSiXjN7fzkxcQgp1BrMB
MArayPFUK0NdwnL1aSpdqc6BJpqqihiNqUIJQqZBmbLTAhSWwfvvuRpzSKMn
kuMNlXJIhU5L4FoNLPc2eWNdufpy5Vi6rp5iBXoT5qmPfWo0Yzy/MVv7wt+C
ZiKUlzXsumk3u8+i6/LtMjzOm3fPnly6+5rKIl5TzNFL5XzbGvkS113sRf80
6+ea86thqGRPfKM89KjJYNJvG2LIdmOfT05UEEvsz6JSvnPFfRbvqusOyR7c
knis28pnwu0aDdHdI5Hey2A+cvXTuthYsrGOJh0KWJ4PSDF2zduPXk6Zor7C
9JE9GKNAzEL0FkzaFa0XQ9vrhtHB5rJZSCN+sEcp2RpRr5KW4cNJIrx92QB8
JOUY84T0aF9S0NCeNOFHjQ9BxITP7Zpa9bsKByiFCGvZH0t1tImlNYUiGSVO
gS1dOD+fXeXcGw1aJURAOZf7Ops1nwwVC9r7tIaJjAFLk5FexzOdMwSv4vFE
R70pEUjz9GdgaTkZJ1kAIXLLyASH7ibm9qKeKpIvYbRrDHE2uOgqyBfB2+hF
yHdOo7SeCcTz7RLayHDUizIqA5abxCZdIXDq20qKO4tg20/gr15gu7JBQSjt
0xCPwWAPElxVDfMwAFbpgXnKhbnfoOPXZh4TdA1jGavdGhDar/oB4wu32jP0
GiHTgkVgOxTrY6ijzvJ9V8ujgiyHarahgDIcu2dvgNSAlsbhQ99qI9kKlXxG
45ip9e6F9zmz+hlsNATCVEjtw7z+wn2BTU1mJiHCfG2hUzadjoH4wxYNmB/u
keX80+9eDnH49v0x6juGdvU+8pc7QnpTym1l1ZfDt/N5PKUfq897bb6Gx0+b
yusdKXk5IgF6Khnt3u9+NFMjLI2k284qD6BnPekOrDAE+o6RnuxeyjHa+OL3
r3jI/DI00vZ9v6VWUmDrBmNVJyAVQp0T29GxH6XP3xEQLux+8gwTD52ysMfS
cLEyR4dYReUKMNU3+AKgp0sXWfduXPgymHn/CmzgJSvSnaf65jtAyt2uaerg
vzFbqeRWfd3wPYBbF30QQfGucJ9naQLf9U9QghxaeDji6U9RkMfNc9gorKkK
8AL1akxSCUkgGHUPAe02xjcEfuPlgymgo/Z+qBe75R8SJNZ/l9s6URceEVPc
weTPo11KjT63Y46nA+iqwOiGOfbijvvGWIvGAycW9mAaPNHI3/2KrhAVJRZ8
jMlF2JhpOyEoBzFubaGDWEiweMS6FINS/mpi2D3sPHPKhPaFl19xxfH4PHxW
KW0mid74xT73H9TatCnPunBk+vMXb8xVYK9nXJDEhxMiXn8EQ+dj47Q4lI+k
0/mOg2zrB7TKMMAb+4887Lj97o13CRvqkN/QCV4sxcu9Y+1Rhy01LA0sq7Po
JVHd4ZQBcQdzPjst4TqdkDIR7kTVJiEpqkjsCCg3dJkNs6yRfdKJ4dwNQkaC
UUOWwv19y0geP/M5eo3DeWJCRZpo+85+MsAn0S1CUy3ZBd2FzAzo61bVB0wx
JejifcXi4mTxn2s+Z8F1A4UeHrCt1h1WLE125kd4gWdQ3Ck8xqvnYECRfOwf
YCFfL0v6U6jMH3OdO9uhh3c0HF26QWK+pc4wzZF63TPVS1vvfmO5BliwioFJ
0d5hA59oZ5XIoGo0c8bj4a7IQDinnDcIPM+Ba4nbJoHxx5ZsdsyIn4Gk9kxf
tALb/PjHdkGgN+O8bNSsew0Dwijq2bH0PytnTdam+fdxkXsoLbX0I3usELTa
fef0Vib61t2lfS1yIQlPRguOhNsiir7YHrZ0quA5fQpsJww6iU65RUiOB9Xi
ARnMAuAI77Tkf5Ndpb34VdryfG15D7snrCUILCdx0oScpgZbm3O902LV6jMn
maHZoruu1+em40zbF2V3spQ8Iwg74uViZSiyO0xotGHxHOHONGsIo3lzwvLB
uIe5NR0Lj0jSQ3A3SygBFWsf1g3iYy1d+5hfw6DjN7cgrk3zYK+tFYAU4I3g
7sm1SnKc+wcpLNfuQFhCyft79Ejky18kaAnmF7M6tVC4KTl8SZt2vlfzkEFm
/6y1Ha+SeMM1tNIKrtfLodz9f+vUMC5dGSgk2BkIFQM+qPhTUUqUur0n1F93
2FDItqprcspN9cCtHxebpkTuWU9qFL6WdIOTa+/+RqJvs6z2+nnVzKAVquLf
demNzSFqUFaO6KFfW2Z4wPyomxb+2YvOZr7fp65wkPNydkI7I/3jG80v4R7v
VpjdgVcweuekn3wPP1GCqCyW5fboogitkcK4NqJ/Kdf5AkRDXWvBq42nlmhj
XyPIwa57RajgUex0bDAC94rdrAYHjd5jLpf/7frp0W85G+cOp5tYIiXWRgxm
Bv1al0jh09FyBJ+KIB7Jwsn6RKYHxheA+GyUSNnQeHFAWQ0wPudAqDgL4+9w
fhG1hpk8i+Lvsr2zP+19EuHmXjZ9XGthMuyzpgynsDf9b8m3XgUpWemezufC
qTkb+aAN8xFVPe8UkIut0v2ttJJOHit9yW9nfIy3WeEu5k8P8mlRRtSGdgS/
Wl/Tf7WNVh1QqWF5Ql4GFml3l/Pcit/2hfwOZ3CZIS802AZtxfFXswXaCTjf
9pPzG0MuUFjGjf7ErxYZXETC5HmMeOBBHTwEIN/iWduJewR3p9/fSTePXU+S
3ECFDsON3pzQdbgSGCMpuSC242/ISfn5UQ95uEBDr4eabECzbdBk/x8M7sSS
faroLd/6kRhHEuBVM01AxEDV/wwWD7TV+GXYU7BX0M9VYlXYq62XUQA7vKRj
wskD1EX+umUervuDaPD9hFx/frd/uZwFuOkR0T3IQv57jF2vYVFNlEIZ188F
t52mnZUz8HGCKi8GhJIRkxcbeQnrzyILaplU5MlJtWg9SShs6gD7r/AWXQyc
49h1t4IKXvfa5sRybj1S37UtUMCri+GwJf9E9p1+KnOeJwc2Kiv1amCXdV/d
vMX4w8YNM/MrDEI8Ni0Dt54ufp/sU2U81eQyy5/xgl5XIEuNXB2FTrFjt235
W9hRPjj8LltFZo9i+vo8AgEPch7RdRf0IIlibOJZRdOnlnNbIvR/Gjs7oCLm
1hczfrdwF8avR5WIUSktUq66BX1atuX5bFo37sNxGiW5OUyukCnWidRQsmOp
PHUTbrP7gKDdwYPeklCO0MDeWM1wxRmT9NZg8F837oddqD2aKF23FdHIaLLw
eeWl+lcxVEqyVCRECWZrzq54hXFSBoQfyQ0427NogNSkunw9e6cWgVXsJOZQ
+mU6ZqT5WeAx5QF06TcE684Jbp4Y42PIvGnCQN3PpAsUsHwCwKSFzggCCbFg
wGTmuwYnQ6g/WPCCkmd+2NXRIyPGp6KOtd2XYJRuxqcksV2TH/5GhvScMFzr
wotOsrf70a3zSDB/OD2BLVgHoO5yp0BAJrKD376df7YtOMpDFQEwgKLR4fqE
dJCDWoLbH+ORjC+laq9oJMLlE7TFuIzoGup5zohDXdYv+4ldoVDqZo3u923T
KgnLcolVhmSf6VWHkJpU/UPELEQ03cH72O8z7meAnuq3IW6OyRBh+gviivyv
tTUoAnraMoJReLbFdJLTtmNAcJGdJmjitiO80YCBfn3aanwVAEveSYXjypSS
UNlWTdJ9n1ooDNEes4ZlTRROYN/gWq4HZz1x0jqXvGum0+k4UF+iEOWMLFtz
mrDS7Hnbj4bFsO4MawcrCeRj4CLw7vbb2/MKLFATfGZ2JZqZmhdLa5ytLoyQ
SrSM7t27MvJXj1cu20jqUPqDaZL+O1NPH/l9TeNyrZq34mjFE38JoGoayXp7
RSYMhTh1jUWTNxL9SEgZgrI2H3cm++/ftt/HZe8t7xUmLh9Ekpf64WMB9sVg
dDFwlPnIY0sbGbU4SD85jFZbLmtx5eB3VmEOyBQKouKQQMu/OxT6DHBAqmXb
RMYIjvI2TaVjVERiL0Mxiuwq/bMqyJDyHS+8rjotCIeT30bUBAAkRerilSp/
xdEB9DYCo8qJGeuCetD16ADSgKMb2HDU1CR/BwilsseO7Ci3qNz7L+DiZHjs
JHvu0fWxW+bd9TAjldHhhb1kbVVUxCEFUlXX94EDq01PzLeCCgSsBEEtNN1D
dbvsDFXZofo3qSbcX6kS3yrBzju/Tdg6N9+VgM6ZMwZmf0hT6/K7hjdnyRQL
cUpgch3JwRQi1cxyDd2GC/NDxY+Pr4tgK4JZ6ZvX9KUItdXHFXB7lQ3+vZfR
h1FwwlDjAM+p5L2u92oNyvzPnqDeI7SKoUclnq2iiay+l7xgoACVRIk2qU8U
xUeQo+iXOEqiE/rf0xX4WucvI5O7yoxDC1MNz4iMvKm4HhCPnNPUzCkyn5Ae
UlqA+/zHy2MxvJ8Ozul47WuDwAyd09Wa+pWOMuxU9L6elS1ayAXjVyzQ/fxh
TOEjwuD9bzzkGQHgfjR8BXQvmMva2DktVra17WOdpF18wMZccYs6ANhZP0yC
nQ0+cp5pF+4wZSov0PKo9ZcC+25BrXhNJSHn6PmMO+pPo80snLqiIm94vHon
jQYVslcp/J5uY9FPwCEO85iY55pH1M/A/59RLgrlnuM93KjPwaRYUBxCLR4+
6Xdo+YX6AolJVIQHOjFmAfrCXVdo7FbUzEgNdkwfvKX086OqbBnbK4Cfw6+o
yoeaVc8QzMWp567Oz20Mpk6GLfB96jJCv5FND3CwFzvfovVcGasHWWB3SOQP
FkPAkf71EzO5L/DvjpiGXFVdZGvzKOz2HRYPMsO5p0G0RS13hYiaTQ9AY91x
5xORVMe7MvP1IIrB6VjVyEdnLg8OXLR6moXQ9jHEu8zZQWuYJJviwZAedYBd
h2VFlTYIm1lOchAE5HyVKPvDKocpJu4cKX3p2zQFWYVgCLEKACUGBxl4u2pd
t0Nei+mWgKqvSZrq1U5yrsTjmGzYMp71WU893662ooM9OEGjz/D8Niaa/M4k
QDvxirWP5Ffd9I6RNxDlDRWzm0oShkXYqXnN69RZl4svY6QTm0hiVNlZPYke
TjMIqS2BSDVP/l/oMbPaibXHJizIfg9UbYOvybW4CtGcNnQoQU7qqYIVqvjY
c0OZkpm+9mpVk92KmrTQxjfnzVmLIzQUWkOV+A1dBx2N2DrZGPcZj9Z+1eAl
wvXN6ZhrACZrqdJ1VztarPLKZdJIdhOHvFYIPUCQgBgpxhzpLYE11TpQMin1
IIv+y38uRUy4wg3CGa8epLlgupzQphfddZqpQAZ++EPhOdsZ1Cupe5KZq2BE
VDxK6ZB2aLVHY+nG355sytSTgEThhVo+yCBCfHG8qBSQUhlEcs7zmCcqfv3d
5gj32CH682FS8tYuG78teBCe38m15II/plfT9LmcTMkM8TIicYpkhSNUc6aS
xGeGHZuYqB84Hpdwsg5E1hbzvzSi4QJxXdsE5CQ6VFqGZ19ohMB/ytfJ9fxG
qf3G4+Tyuvn+t3lyGYMYODOCnP5z3qqAUlj4LqHlbqhzVuDVt9L/j7gxDIpo
fUGDqHrhRROQAZa664TWy5lsECDIoqClmBIHlLcoY8iPPbXotoU7ggJuUs39
uDkrVYAf2FW/1NTDUOuIwkMfbZ1otBqw2EU12waHp72UoQa67gK1WAPxF+Lp
wv114DIpjkrm2E/vz1VrK/tWdapdM7Kipe2tNL/Izh9S/d5hP0Se+MExSKo/
N73DVQSfqFwe/mYXB2fp64Bcy6nddRLWSIqtZZcQylPntOsJFwQiQcTFeWNy
OvV0GJIY6U5uELyaUcWLbilNW6/DMg62kZJJijOc154VpPL/ufoc0Tcw+a1f
vx9HZpGL5VwOVsilpaz1aOv0pDkbhi04/p1HD+oS6TuA4HmADtkJf64NZg5W
arKvrdHVACF0XmULtqdir/WwrLQrGN5x0c5anxn3WInJWQURBGVwIwAQzRj5
io/RqdVpNlkyCWEm5R10LkJAlTAFFB8uAyoJvm52xzfrzNyGB0XCJYkMqKfO
hN93LVedn+o9Z91Zq2Lo/Gnrf02B2ZMXQ9UNMa2X70TZFRg1g4pnaJbKBC0s
1FJcizV8LhvAW8/xQplXF2+zxnmu/q4C/A7sqkvZBvXQpX3YnhJgliG9UQL0
zDrzJJu+C9wqq9xNw+xfGFo23e1TsNYEPgmge3X8jVxp6ymDDP/Hm4kaJYoA
2438bQ9KiXHqjEexX1B9gDragQlNXEk2hBZeXZ44at4/l0cw/9/no+0kesNn
fAcNK5TacsaOWJjPia6m4FOt7AdgP4BhHN/t5JTs14KK9CyrSyG6h2x0GJN4
th+myovsYAihvOY+QGdPO7RmIVcOwVevCacSsNqiwL9rEtP447EObCP5HUwq
7vyufw0MYmIIUXjfCvgAEN3NICaunL3RM12ik+lC8BNqj63p6TQo0mlYDfD2
+dcnh/X6IuDnbjQymrAiQ4yuygaCRfodq8eTd+KZ96wn9yD5iTi0OaUekru9
te9jfnI+8nCmGdiW93hlndvogqsox4XsUriKsX3T6AL9oV5KpRIhCZVRmr/t
DniKw3LWfPq1sAi5x+FvgSlhUdZOvwJP+PcFc6AnI/9LoIgf9ac29bwPBqWG
dy5JqrZ8MzptjUvwmfyvH808h6TUJMI3MNipfXG50lfY4N8VWTUKVXDlrKhH
lwjeeGECY/okxUANYFcN7yzbpyfkK4LJUmgSWNDObeUCvyuKH9gqjD7hjWFW
RL0+CxH0zIKYjqf6XW6gAfyYau2KRDFMum8pKxgmhJo5w2uUYR/JdY2wkb29
k0RynWw90DzKsLwbcaZdL4tY66V43TJlD2uk6Bwyq7QM0k4NFLJGQpCa9+/2
vz824R7wHio+XPBJaRgr20yFyxqurqCiW+lZ+kIs3vTfUSHaEJ6VPrewp6nK
vsGIMyO5dScyLYUTzZiVCWhtB48QQhwdZow/Z+s45Ns2Jzhw/M8GHVMTj5P2
yrnoJngWHUVtx1nyEGL83OcGKZ0qVhn7tj6I9eEKioTnpLSeYo7lNoRHTa/r
q1Rc3fam3mcFNIYGg6pmWhY7RF/WPz5STX7NEcaF7WHU0p3vcfGK3t+Q79TT
sUTz8jRDCcogsSk1uMuvCbbFrZB55h1T29sFLB2/NGrgOwJSMWelZXHljT8L
cbL+2vOI3NBabELwjiJ01gjkgZeQvoZtsQI3in4rmsDrjiWKGZdARKpIZzYd
EaPfPy2uJnSnjnXbTjivgWbQYTJSf8Fglg/4DtX/E57z09LMQOgW7JJ7QN5P
3LaCo4so8lgnBuj9jyBXEzwf9oVY28C7Etk4lkQNOzTCpc7s7jfMQzZOARKd
6SrQ2ozWL8daI4kKKEff280MsaDPd/nAFdgZfxE+mksBAspelwslUOSCUwqE
1pB0nkBLdWk/tutKoRWMSJ18P9ldQwBeScwq9cW3HZlo2Nd72HAQVr0TsC/L
iFbMXpseASeF1x4HMA14tocGIsJnFg9c9PlqNXWVqg5GjsuA8A9VTzAeCKk7
FIJu/kPsKjZaMNXGTb2mjkwKiNZ+u+ZnQUJsWge0OhDIhlp42Ior8Rz5Qhvd
y+X3rsjfCgkgi1OWS+yJ9fmwLS4l2V0Q+F1oEmEMtBPe5/yNRln+JN7pogZO
Kdjvo7933b7Wb4Y25LamwdgQ5SydvHYQPOdW71fXq80FEcTuvq7iqcIuYHTj
tkvvcQlczfN6sYeHG8kgPoc76vWwrt/14kILXNPxGAA9ao0lioUT0Nz0pQ1W
VioekV2q6WSkvGFBG97UXseKQcJyaLd/SkIKo/kPGzfeg22c3dQfZyE0U+hJ
Z6Ic9gfxy8BsZQlEdNc0fFa6CdXvsXxIgLkTPLFwEXpMbwgL6v50HulJXIyp
CJSaq6CCmqqbDpVA76KAY4z5Ugg+9OK72RtjhtpCeJKPL+N3upasC0i6M7vq
XFTa9UHiDQqyRsHxkoS5bzY6j0lmVHyQmNEM610586i4qjTnKOJVaY+HztpR
ct2Yz593hutQtFDvjMqHRtOtUwpr+2dM7xwla3PJPQDPOvPUKwsNJVzXuEn6
ulqi0XRI1i3+DytB4pkiRMaqkH/51fqXorrQ6f6zEkRsslKscFt5ELV84hOp
2ssNhLwZpDrkEjYkCt9s3DsR5G5MN5dBqzJNfQKzvcvJWpEOSYUunOBZGqRZ
WrwSdFpBPq+lmJnWV6kPxlhoT5SgRi5VrDE+lEG4vy2sjp8qqHcCo+jL2Lbo
gqNmpcP6BVaBgK/cw8a+pjX0cbftaYHu9qXZsszbD5Kaljrk+yA8Dvrp5/gh
cS85BiwguJI8FEc0gGwRlreVXhvUt6zhm2qfDmYPiq+vQQQ094oSLipyGn7S
iqRM4t4SCgg/WLlUJI/JWiOmnK5By7HcqrapnMaMeibnK8k5yb1Ii/QXEEmD
O9P75jnBn3Pa6H7U+vGy7mnMEF5TihuKGvTVyqAhHLGl4K6RATt0AlEWbOPc
lhOMtf0lDvDIvV4FxhZGpVM0nS2xkE/3bJM5rYnPzR2JsGjyGEcDWGnZ4R2D
stFpmjFYPinACBpiE5bzX6+9bSeRh/dtl6W9slkBzHkHJK1U5dNn7dxeW6qX
S/YskTKBqStasfIQN/Y/krTkrdq73Nbe1sSeumREsYSUM9Ap16wWEbCrSHP3
l/f6SXAzzsD0e/EK+I9bMuNx2sAW7muuMHa7ISgm6eN+dhca9gd4q8qu/FSo
P908znAbKk5a+/W+W/LshMUVGO9AoroCRc6eQlnfGWMsrM4lPZ1ZfV1lIkFZ
3GFpcpU37tO6U2WrHFvXCYtdGwpMLNUelmRCDBG+HPXEb6JClw8XRA6tsNlV
biZ0une30N7dZugE482njR/TNSoffya6ShWSBniiDwjKUpzG96NLJmOCHQPP
nCXctr6ZJ8agSP+TxvJfacW3ANkt+zW+JN47Q5nC0bh+G8o2LCIugb8SA5jH
CgpJkGmRMFHCDTeR5knFUy0adqsiSfSnJ8aSdHS76tzTLAyh27giqtCiYl+z
QoHZOPO0vizFkqj60vIClHAEmEUmenbAbgJu3+j+67w/DNkLslZG7pMtVmFZ
JvdaNAPDgouv+Q/cfGYq2dJjYayQvaNjRbiI+B5lhF58mXEt3oqwWi8pQEua
2KR2K7/6TQpCaUcwzVLbR8YJ/XR+b9p8r5i6x3c+ZIPd554FYe8FF6zAh3sB
xsMIrsGeHCMonxDh+VLIvT9pcoDFmoD6DT5NzoynKUUS9/DkiTlfA362FUvt
vVzMGvlhZ7cfpSX6R04NPRKw19krVJr4vaukUzw7FVxysEZyi9bGSpGS/RjY
NQ0JWq1FfDdKKHoDKpM0i0y+eevpltAu6ws7UvxPxBq1l7ciHa/oxkg0IiJ/
Xls4IqXUUieIJTin/88h/aAH7Qvf8s+83uwiA6L1CX4X3wh4QyHteRrtQ1MY
2dlaLR3ZjjED7z0t1ipUGrkTIg43v1wQS5Jv+tqiz5RoXKC6XCEsE52+IAFc
iDD6AVJEHmeurLYS1brCXShoFYAEyBwmRwdDtBsbVwpOZG12kXImRD/0GDwu
rhH1aBxlIg8eOpSgbPAcPQtX7de7fX+H+ReJy0UteddzLEK0a0tGhAL2B0ul
9EUY7tfGfWa4EfjK3aaW8OTkngoY+24SdofbY+snJUKYkDBcjcyVSSiyZSeo
GeUD/SiJgLZsHnvKjGRP8cSySR5BtBkr+DpL3n1Dgdz+Ge0bhH/drO4i1JNz
uQBOwA6uG07VJMY+JGH/4zKawSgXk8sVpkJBE+qfKfnYcjnZCmdue2jhjIek
xxGcUdkEyuC4Uu3U83kapNXthVSTnr6PbDXo6E467ohukuRVRFMsaOL19mS8
i9hjvS/bKrjrdIWSaMFZtqQJ3HpBpd81eGg3zjXCJW9DQRjAivrAmWHsuaG1
nVxy7qg4vGQa2oHRMf8yB46Q7x0yohHuJUtFXApguEhI6cCVWlrJydkZhG7e
6g0I25PI/NJ0S2h4uPNaIDd6I4DrHcwllmThX56bX+jpZuE6YdKvmWMSw1aY
FZZwR0LrKXZ8wvssglWHpc49BTQxaXrCz/lruZAF+vzcJ2uyAw5an/s91V3q
Y25eujwYg6NHKocVCRanXYlMwnjQ4CfPCe71AzmjWGiuRVzBkrCuZhfTw7eC
3LfLu6ywxBP8pxQulDBHArdc1i+xb3x47WvHGDL8GTrtjIGgQSyA/3bf5Kke
xgiUUWcQwvRjSkt85kLwDU3nsxFvCYbGtEeupIEy5t6y10c7CS3euRKhpWwI
2f8ZDPgGWVBMYQKP0xYsbd6e89j3uhhhjaqja67ykiiFzxNKu43lI3Xm1/E8
s+FnassxPg+u8n/9+HUQfCMvWK35pEBaBEWZEK/w3EasfwE2xaOhFveR9PIH
LmkFQuCsLdq/l4IfsXy7Y68SpyLx0Rvj4FpkLJ8HU8WMbWgsvRfUHK6esbX0
YjzQZsj1xhcYZzqb3mh2czILiZZHF7WONoopCjnMDD/oHV+QmTxgxxdO0Jg3
9XyysqyCvk9LJ/FhSR9HLeoWwwLyvfVAXrb2Y2HFnlAdYHCzk2ylUwGTfpT6
LAVzlsarU05G6yqEoKHwwd4lRK4ztD2nwaB13fo71/cm6RFsHvRDqtQbJmNs
u3UDhjRwdikahBANCXsGECcNNVcMUINswpRLiCFfn2kW3XWcPKQgin/AEKAY
nlAjCj58qD7XBx06SFTAbd8G2HzRDCcCbo7f6OSNqy672XbQP7d5ASPWIFCX
cBeqhy6O4Q9JIetGZguBRiqrgHiWETZuI6t0VJJFqbAnoEwM1Qd0nBPWGi2B
f0TYHZUcBEkWFLawOjNoFJMUAMVAoR+1igv71a91oYas0Ackg918J6Sao8zR
llahUwXu/8a2R+ACF5XQeO6bjUX0fhnlbgXK07MFJcsmCRm+cOXAYJHELE+w
pSCx0BCXefi8uPwFan9spTnrG8AMncM+JFWRp4DOaP4ZK+7CeW5SGXV0VtFv
i4yUWseqnKAkGeZZVmFv5MohAwBvbfoini143FMcdXN+h4WVh2btxDn25NzF
w9zLKJmh5bYNFlgzuAqualUXe84DTDuAah/Pbv4askwaBx24QHFR58FX2aCW
1Z/gp3m97c9DJxnYSBEG2j+HT0xOSqZIu6pGpNgML9KkLxAX7KKD9p6I9fDA
bp4laQOH+BeP+QPJHNxO5DH1N7Jv7mxoM9hKykOqrMlYrEI7yrBVuNOL20kx
xHOucwhMDJP00tHV5zpTYNUkZVZpywE6epoElqmDiq9klK5R04PITuElF8pn
Gtd9vNNGJlnW0DBHg4msEaS5+JYSN8F2rftHD+AeSmDt9vg+0fU/nCrz6EGQ
kIqd9uqZrQuNTGesJ38aXrvzSZPE0kjyqlz/w0cgkxE3G4AVf0C+TKUKF3cB
Qioa38a+/2sMsorBIMrBujzs4gMy904OVcLmOOsXzsFOjPZvVLzBaK0A1Gab
uH5WTfjsB0naFJSXN7Zq1wJUi8dPZcUW+DiKcT1k2wqMDpc6lZRfdpeZruUf
si/ayshhOE1MzTaJFBzyNsocaL6LPXje1j6Aj7RI1iwa+1KFAPTwXozYxViC
Fndmg8TysxGrjy/Rr73GvFwx6WWxACA3mqKlFrCWLFtModTHaSHObREGewWU
6yTpk/VMj/a8vsiAYHKIR0lKLG5k27/JjrtUN8WRme0QiHqJcFOn3YCtAIeB
FiLj8lup82e9EFDRVq8Q1oghB481ygCuWPGjL3b/VjqiHENT0TH73NgMlVDW
8p3mDsl294OM0s/xOQy5pN3lUK9lBeEAx1+nlZz5dvLh7GISXp6js783MsT7
e0/0s6XMCccPsE3g3LcOO3gmelBZqlfW3l2Wio1DweZ2ikjeiVOoJr2ksot3
fJCYm8xYlMLVLlKO+8xLd7QmQuDHMm6bWf5zOHByMXeylV+pGcoOyyxC19BQ
zXm1Lyb+s/CCfTICG36C1B4D1XvDEqbXtSP+ThVWFM96zPC3plwU/OThFBC4
/vo8pc8UG3RDToqN3B2sN5emb7oTz2S6sxy2JCgYMyhDCo5FixcmTMLr1zq2
J/oye3yJrjNurBHGd6ZLb2n7JnIj27J0Q1tf/RTpIzppMlEJo2S4tqFDTXEP
cDo+oFBgnI47Gr2fDGY7l7D6FMYbD8SA0q6I0T4c7xO3csAt7KEcLEHDMGUt
NtV67zZ/KKhQ8PvVREZpg974t/zMwAK3eg31j/zGuxN8lIsuGLsr8etflh78
Qb9xuTLTSmPv98u8H232oYUAugNZLkQ84jKxEjElVequ61QaO9I/CLU3pFwe
KYua1FQ2wigq+lCFJzZ0zOz6+cziX9AH+jq7h0a5ypkgXzADfq3SzO3ATRoB
cdsbmprUCgwLM4hSe59nlUd2hn2GPjcmNy6kxR6zjoAUUwmVp0o+QCuZabdF
ntHINzjGw0ua2ClfLQsR1PULC7qKIJLlukrgFSxy44NaDDCCxiFiPrruHNUk
246k4POZ4QnQGUrW1tuDvEzuijnz0b2TakjqR3hNDgR2T4FbQT95LmSwoBIa
yaSBU4aDMhMsLqJ8HQFPTtozzOCS81bLnjP6oiRJah1g9Q3xHVB9OuFYezoQ
YkocZFxhCqDqayFKl16oGn0aui3qjMYzZC16eFZjxu17fsfPODJocNczRenE
vOLfHEWflU/GMXQDpWGpE8JfLourU07E1XMY3Iqr5AEOdAOeqPvlJQvAIaoZ
VBYUrmF+MvBJAEZZ5KCyjPalRIUjfPGj14Tv/60Nd9WAFDC+m2J+UgCdoTUx
eigyJbz0vDd62r0LVOqn7EIL3FRBTMZZrot9tFysOfr0t/vbJXEM30ZXCuui
9u/q04SOF9xnVJal/fpuPs8IwP1foOAQN+ZswA6MvKls9d+5CbXK9e5JCXIy
N+om54UAholj9QIHxNRpATBjkq1twwJ2LbCnEhm/B2hzk67zzrDN+4rT8iYw
AmED6cDgZKlpBVmJaQYkscRwpiBh5868m19favlmUx7rYnSAP3zuBbde7W94
1IXT75dzh8yw+a2r4u6GUmuymO5J7hiW7sdT8x1TdVrxwYP7wNviJenjUe8D
grCJ7Res1P1kq2MmMwPKW/yBWQZTAPT1F66eWJW8+gL+UyTzVK2Rl4IQhQba
OLCpAvRmrPn1GHpi3a3dX7/Bp6h5PpviB6BqsSZYqf8YPZ63nVEw8S9pHVJv
bprp4C4IYtX9AeMGezYovS8c5Za59i/JiNendpim8iptNy7YWJKVOxtyrJkj
bgm9bc3el9m/OOCw798zWPgYLkR12KvFSNQnXld1kXZCZY1Wb2KyfcMVmg/T
deVKgNhGv+zGeCj/CiZRZEjt8aK7Gs44lhEmvfbPq3c2w1gZP6XJd1bq4/fR
GHrhF2NNcnaWMyDvVDm9BoEH/bQDSIlFJxfdPBIpdWOPPNrTprDAdyMzNeP4
kHUO2AniyE295mcRMe/MhjhYaiFAX8x1kQiDd+gmULeXf7UfhVluMG5HFmEG
vnXoLrUFGa9JHqxxtY2+k58VMCpGgbSRDGVk+gwf+gtzR1eSqStVk1VMjwKA
8lx4H5t5QKXRF2GIKEqWqHNr6W7or+cAB0ENsYs+3A2TUzJVra1rTLy31PvK
0yKo8LSnAgMZcYx1gJ10p/LW8ICmviz0lH4IIoMjUqrfHl1du/hAdF6g2fcZ
fY5LZNN/OO2hqewmBa7uRxvjlxAbNkj2dKUeVlVXErasABkdQ7lcmTLcIEz0
VXmQpwaaHBxKCeEFA3+h9g62tpoZ/b0QqdD51arrktaIh+WmGWTcGhJx+VtZ
uPHPSP1hWnq00DRGenYQJw1RJv8ewFvxzMO4H2nb2nzdGDnL9xvk031nMTri
1e80L4kEg79iBEY0aw8Zy4PXWrL0w2hywZU4VdnSWTlHu5mBB6/2XDF0OPYq
cP1clDaithns+DkhZon74T2gsfdM3H3YopYESotq43ZVt/xH1zoNRGMdkRgs
j7RUZRHmkxobwJDUQkuAsKBpfOuuB73otVuWgalBcpbNoX6MZsL3v15qncYF
qS060RzYDK6J9s55fm5+Xo3XPBigcnJVANlhm8mfr9nUDKrWI8yac9krofBv
/qhiFtXwPDXHe3+ZWLUsCnqTw/VpONhTRjV66MkGNauSdogKlpgO5taKNJ/i
GpINHBW6uuNVoLtaWXsiMcJCoP4hrcOcZ7f37EkJbFVYF6w+xzUzdm+LZU9s
VT0AMNHe9ZLR/AhqNHTKXDOBfDl+Aij425lV6TJKwrHAJbS4/C3U34HpoljT
ZYcCpWL7Xo3nkaFuGwyIRn1mypT0KiJKzWLGfkZMCEILrXliINooXHO2W4hY
IezXcqBq6FOfHkxrA0vblBhPjy2AZW5AgPU+JbE56fSZmbdo4/v/YiBwM4zU
yfQtXfEfJvR8CGarw6m0V/iAfDIRw+9xKYK56xhBaGjh+Cgo4NKaBob57lvr
3JqRm2Sus88mJY9+2Go1lmIu6Q8MnI1auoimhOQPBjKT67ozB4oGS0AYz9qS
VKwJvx7upSA/PiTfBx1Z8rvlDd3kbVRy23pH3XWIbZqElNafUFQl5HxAJgxn
JNhnUV07D13mLaNp2Y4h9/yrwbLxKkSsTa4+gw1pITrqrIHtbeth+4f5SyW5
4+LyrQAIF7yGARQAh63+PRxHg4EljSFU/Eh9YmVYBjtgYDvk5s0NsQXFIJyQ
jKjXerT44ydfQDeFgh2hCb4Dtn/YTaWbvRakfTQSHe7zKcTboibABBtSKZL+
dWgQJjkRQJd+bSKofzvMHkMD4XPDwBerIPIiwUa0ay3DAOgFmWOMdg5P5det
L2ycZ/ByMN1dSDp7E45pee+f1+vMyU6AyIG+T/MAZixCNShzRrz4ZkR23yO1
OHxzRjT9Zl5yTIqnGn53IemUylw+9pZbOhl+y32YiYwOPr0+kfRjEeXAgRwx
FuL32jvLweecEBL7GhcXm8c0jeYxQQvwfpSbDbk7Iinz0jx+uhg5Otsn+sEU
UvjedZTsRNjakT1XMQSMBB7Wob7Vrg2E2cKKOKqGG3tPvFUd8O+h5tGtnpdD
JTXt7I71lvu5YhL3MQgaxCoElCUZpkoIcA165nKXRLpIfVvEDCrPR5ZMLw1J
K0I2lw74C4VSLYd3ZBMqIBM2hml2ZZ2FBgaqaBWSIHU0OPrG7NFCKaOkZfq3
CLOgVL2d5uvmbfmiR9CfY+/jIhqrFp1F0Te/t0JXEjF9Y9s+bYlC7npk8R+0
gld9m49oY23KBaCpJCvXGxIOB3roxpQ254B1w8lpyiW1THLVPZHBrWutApk1
V+T/IYjRZdg9duOcRjbgJYqLn0Xz30Bf9YJpC8OijbDBfRQkzjF+Qdl94QD4
NEO7Fc05b7Qqy3f4A1Gzrww40JzlL6xBQt8hr/dWJ/GsgeX9GoHWPNMBvxfC
XBkD3boImHZHogMGdoZswNiTsEVOo09ye+iwPzCfdG4M3hWL/3EPXslSR0x2
vpxeEayLm5w5otjSU9Zxw/66xlqhiJcigB9tjlsriAK4+tMFB4cwGHeh9qpy
rmw5BMqoIX5/oyNQCcmbSFt9p3G69hQeDxpjDKj1imAu3uAvyfE79UEM8Qqk
Q7DTza8Dm8g6eWgr3V9C5yuG44xMLHA71L00Y0m6kwsp2mL+ik9KJNdp/OiG
WgypD0gdcr9/E+mkoI2d12Ychq6mWSRbjQwSWxpvH7YqWBqkWZ1WTgZY3iAr
0d81Sn7Z2BH0/mOlibw7M+68C904IT308PkhUCbhoCD22fP+BXgD3y46rAq4
DoCcs7JpyaP3JkypFzSDuyGU3DVzyYmSsbvBIIuGB+711QBvsJwB9nHp4s23
8IEQi5GNdL74WFLkpNuSi0StVt6TBmsX9/LuMMgDwCnkwebZM+uzOpPTHfs6
NPfc3tx3vKJ2bT3NZ03qJVYwn0b6RqN1hG1wHSgRglaXhYpG1gXcxtn/VoOT
6yqhT2YWLRuWRfqHKyF0ZnhDOxkHIsX9DPs7W/cuVxwEl1FkPo7O/TTWw5lU
Fm181MyE93hWWV5iYG+/x1iThigpY0AvSyhldNCwTgecYIW18p53c5u/lM02
YkGRuNlLuSDjdVRWzsCdj2iEmaEcg0xaWwcdnoM+N17ih5kLr9w2jiNh4gUH
OMiByZ0WThLCV5eTYjbxMlq6MkPVWwbRumBbp/S/PGP9zHXbJ8Vvh39n3hzS
lHYn4Bpv/ypLhvG7qA3j74ZqHIxXYkfQwTKp8juPkZJZpR1jDpEMPPn+b2N7
IuQE72hKrFLcLwoquL/yGUNQt1oh3v254nRCqZjWcYHAUiy49hwp200VGEZN
QTP4QbbJ2VHGjnwixf10qh6hkiBXZNTltyA2r6r9RLq5l3Y+2/+n9DfK4t42
cBvKBF0tdgecrm7yM9QVJcN66BT/6fqrQN4zcbG52E+CMM9zaG7SS3F5fuBf
/NQNVNSiJ4XwdW6So+CbF92xo8WV2LYc3iIomYLUd3Wyc3Ibceu1/+NXwbFY
f9vqV7Gp9qoAQAjb2vpcujbHZsq9iZMRAQ0lQVta9ILwmzkmkMvu0+1BVFDy
7HyEGrGpoed5dqjbuEmS3VSxNUi/YizLs1Ymny8yvelxlaYxrhdZb/If2EY8
oC8JcPlOtjZcF5UUZq30iX2npdozUx2Ue76VHIoLODNGtuSdB2nusVlTFAhK
+dlecA9vvVQ4hiAnE86mIHy8bv2fcfIqFVCBRolNFkIqx0aNkrmGV4RTx85r
4wcBx5DqyndWfhLWrL07jv0lf3hZkGOcaHPBgQghMr7dDyS4HSUsrvD93MJf
KE4J4GNeh8MVsxnBH+m7tMtEr6qpDKnxjQ3nW3O54qAFjl6/e2epPIs5ClzN
BUBPNiouUOO6mWYKEUMqREju2+ruEk45HBHO2Sjqlh50LGyAVHa5yYfmyw6E
dCiYrD5619w1A5yi0h+6g0EThOG/ysQJG2LQ/gGh5/+RX/r1laI0R4kYjEUL
jfMW9mPAaI7en0cgf3NqUduqjWPQQaCVJRBMOBWeRhliro0BbjagCIQfV6IW
C8A/297EpxA7CC9uUq3HTm4EKs/2gmBC2R4KVPWY1zDRN6a2a/N6aBLBLXa+
U7vMQ6lLBFbpaPK/R7owO2xfutSPaDwyM0fmLqaPS6qpc3S8gMTzaUUlhCci
pwo71od7ttwoWTK/hAn+CFazyhZFv68VPGssIWry0Vxx9gSn65cNkjHQ74UJ
Y/5ryRS90zI7pQjCJhiOpN5L7gde0s0bLbacTu1G6vvqoMUz/04dl6yH2ezA
IW9IiXrjgCMkBgrfpCHtnI2wW5mdFL5A0otnEOI3fEZKNqcUOmHkuDxC10eB
NpL1DefdbPCJozsWdyKNelq26iQTm30svP1290d34YEvwNA4oqRAkpd86p4n
zbL7oaisWAKwy32VhlELTNRvqNvCIGiKlXjlvpA3eM32o8dLYlDSOcQe4+ew
z9aahPO4lsWUla2OzFcG0yx3s5BiygartoQ6znwBiGeOKHutkQhJg2yxFpLs
Nat/zZFMRD8Z0ohCpQY8dOSUTaUDQguiHWjQAxl0N93r1zcw+l+P//P4LZbW
GL7PNXc54BVGkPmEXPo5WaeNExeBG5+Q6gnu+TmR8KJkNeERebr30Z6yuHuX
BlsOGpi/CPIZu4VwgAJ4jJqHo5zJRJzzLiFrabIevDtTrcHxbCxNt7CgLL9q
foZ4yHk+sBXlu7yukTHbml0xZba3NPh4zFHq6ZMkQooRh/kRImIcjrEAqSJv
nEOpXqCCkbM+xt3jjIPhJmFRlY4V6eSMEO2G3psbDye9mWbkfbYfwn03/0Xg
5ACfB4x+k9LLUC5uVp9ToPzD2nbYpGtPVpvzef557+/6ftyiofLdY6Xu20nZ
QjsQggxyzWZlsPF5ZGUGVVEzw05mQRG+kRHgoMRYa5pVpk7/s6a6BYOeeZpS
4xi5Wa0WNYXHpBEaEQ23+TV97r6ylGSuWhGIgSocfLg6nIOGk4xk2TM4W5wE
+fueVGJ0n928dM9uXxcuyg+AtcR79wZ1kwVEWDYPkKV6snd1iWA/fptSkb3L
gb0ZGynEREUW3LFb1mU51R7XmsJLNhXrX3rsr3n/geaaOBzPPPMm83XFIOP+
/kxWeixeEX6VWKSD9bcc5x5ABqpxAg0pc1JKChV2hY0aWS3MLcPwthRxXb3O
7VazWwQZFv1I/I7+/ZrN9WRBQ/Nl85Lfl2wZ7oUHtqjnK2H0Pw1yQCpJ4867
6v6IpbDaRGIRDjz83IrQilYC7vYcOi6ckPXDNytm2ye3u2zMN9ynQ4QQiWIU
FB1fCvlS+EWmkvp9+wPzxIML2d8D8dGdQBujFA86YEgUCTpwBdBD/hFclgnd
THgWlJwWcFXsLbqL8PNEsI1ZryDHZKzuvoXD0Ei4/zmPoLYQ7V5GHBK+771r
5G5PvE6bTNR2mJbxpdhqnqYMcZsqkC8SZ1Sq4V1OulSqdcCHhXL69R0gR1ml
8KlwQ48pQuh+HdpvvFd8zudLs4iXSKPfZ3Q8jg0CbyjomrB3NS0fu9+G2CxP
zAQ3Op4P4+B/UuVcb0t3jFl/iQ+Fn8T6lqeIImY7oeC+OuRIIt79gNdXmGIx
vo5XE/0k+/dtgQHlLKlkgTLljwvKZzpHepne8fBbui6vBIHVAXIG1FNOgZ1W
hhj/zKSs5pdZTER1PHJgL5w7s4IeYXK7piUYVfHhcAy4/C9H5jhE/54ScqaG
lxOhdMckJSvdbOLKZCdUvKrbAPHVzPEVn19MH/z3L5dFX2VQ6QCUKPZsKxQf
94fzv1h8Vz9sMUw7kPs3efgmCkxC6fAFmnCF9Q6M1CW4Ouj3Ptq5U36yOBD+
qEBPSoZesy5wyewKp38OtQtqsjTKgoUghIa4ZByjykfx8rrmZ/4jgWFlQ+FL
+RYd0s+lBqdpKrbMnG5o8VIqT+3Os8odX5F/EO7OftXvMh/Jz2+6cGDlVHOu
YMH9OSHOAu5iWencmb5UlY3FkAO7g4cbx+dT8S8XlT7nREw/icWJ60qkKX5+
+2GIVWBAsdWLHzDoHfw2Z5fGKXriDc9XcnCo8rKx69iGQlRAfXi3TQpgQSit
WSB1bLvmIKyKdKREr8lt6I09tTgPf8davXaNxPRwpq8ZZqK/idRk/1xhuJGk
gI1uLzk+0CpLbE5C5ASsfDk1+Q89FKO2btQOyc6fQ9ougboKxLav+ObPalPK
vO5uPfpOTmbKiWPke7kjzbyoW+vbJc7BLTqy9fUjoNdcp4DLqeAU3FuISxkv
Y5tYhkq0en+mauPYR1auonVbJSPe7CuZQlcSqPce/d+w6cnkshEDEC6lMois
0tkSwp4mQosU7rsfOryx/e/vY2SPWLFhP0SOfOtB924BzK7eb6AKaFPGPbgt
MWSNe+l8KVJj+e31PiMcROQCZfZy9x8Ak3nGDQQPYf/8h1W/Q9kCHVIhR9PL
pM7rDp9iyP7C7SMYv4wtsF9Cejvv3CYkhE3Ggt/SdWeWQaaAF9vmzDNMbk9+
qHRBsOu1aMFUQswWg5jton3O+1gr+455L3lKEKS/qidOgmX5B6vX+qW2Xy7s
xg+mzj5irMLYkOu1OtfRoMt/1zRbNlbrvCV+1NkVsqJkGqhw/KNNqtflbVl9
/OlhPH5DC57YppwBIZ2ahtRIFbMpY3/0IAd8UxyYO4qiq1wYaHzi5qxEPOZe
F3IUmozFs7OR9RfSmCN6JcThz4EAZTjl51Ae56X8zmS7rjrYcdDPqfh29w1a
+0/LhBT+Bg4h83fA8PzaaTjmSF9ptI4xkiwC1G0pSoOMJOTQtOEn+nuCiIvD
P+r7AUWnfRRjsuDLyKNKuAWqWsBG5y5DiS/JEujN24l4LJhtc2d4ohVp/CGC
vMPmdHGEYtWttw3KXWUBjGzu9TY3W/en7N/U5NMApTeW8v+YzAR20r+ljaRf
2QsFvcz43PcWNfcCZdUWV/ZUcgx0VyKhQIBzFHfRjfkx2FGjP6dM9Qll5BzE
yCTXfwknnN48PJn66RfEHus+zfkCFdKnrykkwX9Sd6EcUI/Kly082TLtKmYl
WtRj2QTL9N41fTZCfXoOOexATMhLgYDa9ALQPBeCuAC601LyrWVgXxAj5+5v
sMY31CbtrrXpp+0Ls6rvSJTDYEjOI8cmGMV+jbW7qf0l3VErYmnyB6w6pY/o
OpAVIsjkcuDbhA/3iopxBzpTmQ48qVw7WoZ2XVS8RB416vCQNG/nQ4kSAcuM
TL4v5WzbVYU1+atjICIWJwNQtH+F0RFWuWeYmN9JGZE01JxVx2BG+mpDn8bv
jJCicTxsqBzMNk6ojgPmZqSeiEEtiZGeW+frGkl/vguDUatjf0kZ1B8mZq3q
G9FNMu787yDnVaQhLFb0Tdj/d9XUZ4ogPRSa5XOUKHlwGX3HHO3fUn1w3mOG
XM1zqPC9h5m2jYtfTkPYLAwfenDpltgBHrS/eSkjHZdaJv7YK302bymjbl8g
18gCJFdKnOrMqH26677VsXEtwUmJGuqA2DKacKlkyj8M4/pp49LrS96CS9pi
cZg/M4SVOEETnkpHnBCpOzeIofPIfvVQvPPaI4Cy+Po/1tC6hy6ZHPKoqChy
AgcV7Z79d1hAwfLUr5T98Kl17XloN+PzqPaMLNM9/tDGBSTdKRYuD/srBTRw
B8PB3osFSFi9+m01zsI56mQAFSIObXcF5tHjCv3G/85zRbVz0etKyWnufGcw
EBLFMm+bmRgyZiX4NXnpVp1b2p0ssMRAuRwquhZQ3v9Lm86QTFyFATJFOjY/
vrqywZ0RnjAUE5qyVCCUg/L+djf7ekSfFjLrFEjA+yNs0+LjXl5AXpE87vgD
vrsXb3lBSd2xzZFIFofsXMDFOqyW2fOCnuEQRTFj2KOkKbzAwEiA2CiAWxBB
QTOHR8ej9HKk2rqoHrtsIqKND9RJPB9mYGK9wEOd6dB1u0mV09rBIJ2Z9890
bPjdTzf//4K4rJxvXfCJHhLQYpma68KNJWEJ/GACDmBEHPSjGSg1mA7HVwBu
psVG+9f8o9xQqKkR49OZXdI6+XxqX2/eTkyoOdZX7ZdfrnAfnj9Yt3CJg/Y1
a+fjWmJoQZz7yo0m3Ke70mx2j6naB7bm7TMU71uct/Rb5u8b4U/2SuHa+Q2H
+o5wjGaXUgqsheyRDmfs3o3ZDYF4bHIxm1LZ2ELIgPUCgBQkzJ2ZU9gNXjCX
LhwUEAohrRlAAxPQmZhWcxdGzc3E+XrKZ7DaHVVa0Dr+uGAVq1BkHuYQTcnC
X8cuavsoIiO1qCgh0CYDGFi8wBQimkJ7MbjNplfDih8rkaras8BaWuE9lUXJ
Ppowv2ihPmj6mwy+lXsdV8E/kr5gY6gGF+EwZAq8urNKFC1O8ix4HI2ufU4G
hltvnl5gczeO9qQl5zEXUA+cKaHGYGxsYj2UI4hzKIeFgz2x1ktpQNc+QsLe
xrOmAJnrm1nIK76iVn5fl1jFwdVdU7Fev4zPkM12F4VenAPTGGMx23HKdAPX
fqf3YMsN6gRrfueJHEfu0PeIk+k2Rsx6UNqW3GAUNbDmH4+bUbaSU6dVMjM8
FqqaMyV4PHVI4v7afYk/TWPtdIuIYPKHtfTg5mkfYavk/bLCpvotxjUUdaoG
1ET3UfqUXjPsdJogj8o3wLa/F3CUTkPwdF/UXAij/da6RDSmmdtbBfnOwnNl
BLhfrPvjMTIa4tLcdW1lAPCscENBKvPPfQKxdeuQUMGtIBF5Cz7eRrhCaSiH
q0snGpOznL5r7714jWQD3Mm2Ig3YYOfSMbgtBE+k2koQftH4NTPrEwa0Ch0P
UTP7/HshZz/rVqA9leqY8iNIFimOkxiBn+GjUksZyusBvutclsj3k9GZdCNG
fQwAJkFeTLCns0vf+3PqLvs0p3G9pIo5FOSGprVjpzdzd2Hi5M4VMENbM64/
ONBs/u8SiLXE36cc5kFddTZMsriCHl282nxVYGNAFetL7JHTAxrkQK80+lHY
qhxT5A2ehyLidWB43i1Q0GBx7nyUwrlRbVrf6HQrH2zTU2YPA2fREYOleuwA
ioarJRdHtK6ujxndex9rOQg1wq9HzwVeafT6ktMFLMgEjUhKXZSFAqa/xrmF
CC9Zs1zPm7/VgTLmdIKWLMYKvgNMMTr4+Fi1riLQJvxoz7uWmbqP9sijlM77
w1TEd4aZ1uyg56gker0F5LRpC9IC4ohenlVXv2FwK5yTHZgbsIOi4GDnNOiJ
S3zlkN5+7Vu4nOl1f6xd/5Uu4nVapo2RwWI3bni3CDjGdg5qjFayp7wGZfr3
vNOwfw78VDqxHRT6YzQnFjz9xZP6wv9jR8cf6S0cv7LKvroURNjgdU/lvqEv
bR7Q9tT5w459DLFxZLyfIlHgzUirEk53hYtIx65rBlfpfMYQUmxnRDwtlHP2
xu/d7+Dkm4ZY2WAEofxZaVmzGRQetUO8Vkcifnc5YyYoj9Qy9Pt6xix8WY8C
9+QYemC2hqO6dR+1FGZT0LjCNIz74nwhRj0FHWN4Dg2cZrbnVaRH9LtqsOtI
i+SHeuJvZfqkNf/mWMOq3UA0qPfpSNIRZeN6h3lqs7fLnm7cTqt3WRyDy2t6
QiHuBKsake1pyNnYbwZzssvhlzJF3NMbnaUJ6d10yS92B64Lex9EMuv33Bnq
/zb2v5zAV11/9bRFBSntcrv65vpzYDlpqZ/C9OCE9qk1gDDIc/iB1QrRM8CN
3o2ieIxxXD7oh18OKX9WdpsXDBRWRLwyBvcCwxYUnAc0y8KAYMvjAOzWpmS7
Vl3NwkOWiCiykp83B+JwsHmhxXeaQj41T1FeJeC//SfMIhgk2FLWU3YhZDur
2Th/hHOnu7+u17rmUU3QX43c7BHveMKXo5CXihJ3H/N7V7u/d6KcQfxJ7lsk
gC1j72AquV/VJ+QW+QkqGSnh4bmk9wvI1YyNTJzRlQuUbIONLf36riQ2eEFl
5zn4+8jQt9NYEaaZQmG8LzkAr3wap4iqPlRW+EuSYfgVjxWx8UHGcxC84Z+O
+LFtVXGL1kCzDCvdfjUsXb9kH6M7PQqIws5xsyyMQikRMkudyqA9ESAUUv0V
hCtZivpFEt0inLNHhiwM6l180+uRFHwN7exAFiS2g3iFSIXgRlp/s6ZXX0b8
dDsT1BfeQ74MnPpLV6eZHX5GvpOhVp1tgSr83usmod5b4N8vJaWrMMs9Ue8+
ztZnT57mL+GJkhsoC2Cup7n2/Pgj8PPeKJSH/L1LFmy8lRHB2YP4tw3FWcB7
Swzn2xYx5YvesK/h3Rc6KVtiumMwJhf4toVCz/qpBzvMVozwn/QMdfB7HnMa
FTMP0kjzN0SkX9AYUPtf2Y/4rooNAUK5ccBBDXWssqXl/dcTKUeQb3sKjpt6
xblaKrI0dkuss0rzBRRGqyNVu7X+hhJPhQpH+spbaNZiYx4NF2l66bUuP2ZM
WiYbFrFL1JEtkryAN3o8Vjc8RxZdPX4HifOZvCRgg331kn24ldJZ1KwFk9uH
eotJQVEG9qET9B8NPkKBf14KaQRMCoUs7vToYwZ5Qg82pRByaQzZqMG8wHs2
EjhF82lp3/3gF3zBkX8ICzBYzAltQhasEHgmsZc5oxN2GcslUFd0qDb2STZE
7OxehtJXqP50JUYTakFy/fWteHTwX47mcqxHQGTd4Q7YoNGDJHFwFY6rN9+o
FtVqfNjDLX4D7YdggkDhqeCfQj8Qo+o5rNjPWH4WFZVTQimDmpX9zFUeaVHS
EDdSbU+fuHCvQA8ksUGUEDOiPF+jVGTnej4DtRrHtpg0/PnSzRe+QzOj46RZ
jnk/4X/Dm81tBHJcYse9XSyh4T9MAg07KWVc1SELkbndRUm3oE2qTtqbSPxD
dsFALs+/XgB6SoTnYx99zmiKpdz52Hb3oixLNwiNFNGxSeJdYFAXdqU63Yoe
KZQ5p2IBJoqJa2ulbMaFqNb2L8zLM/rb9jh6XdrK5HUZmrjOzCNuaQdqQF1a
C7IcpVMnz9tiG5dquxen8lmnZQg0S1KBKyTSIKDGSHmgHbLp/IULCFTbVk6s
LcZfnWHwymrw2YtucMGe1QCFVK6Uu51XCMTbwL+H2eQQGVTfcdhWzdX686ta
Fx9IhaCILtWghKPt13A0Xkmu8cXnZOjxAaJaDclbUhQqIKq5iUD6Ptfwq9E8
OS5xjNAFLAyehq8dZ9JEs4X9WVCz+WeWz2TUgZ8Tcq+UAnFU4qHEq0ETeURU
rIJX6ULqWtpEc6PMUVko0zg9FMLW7Q/u4nqcW/lUSdhZ9hoMFngfXv3Ewtxf
GAq2DcRreRBS4DnwHgcT5TF/LkPuEyF6BRzS5zUhPkIhsUnSSCVaedyo9DuK
3ApxKOCjhXsU8ZTuixtt9q1trssAa/fJzUpcFJuF4OL0UfmIOuBby55zRaVm
bcCWMMB9u/5c0w/Pvxj1znGAmL4loJ/ekf26jGu8VR8jK43XrojoHPqZYr/1
lmzfSOkFDgeak7tbExK5dS+IeT8Fou69IWGiwO3r86RK/vjGMiI5cZUZkAUh
b13cb2OODHS5Q4gL1nav15cF3pU9gjok3fSo5UK9JTupl+o0qsBfiolZDiMf
4XSFxvVkZtFZq2Jlzm3qNDdb9Dz3p6SwSUj2QRm03flygqerFMzP6ulA9Ys5
19xvl26Ecp0+SsXgp68LO4+gXNangAPg73encexaPrwjlsdkWFbFYW490dIl
/cr3KDE70bRD4r2oJjoZEVRIAwvai/3dMAtB9SiU9XrRSIGtsfePXf7F0+MM
e5lX5Wx8lG2kTe3YNV/XFYqSH6PlAh0w4PSwHPc8Tcumlohedc+FWVzaGR1z
JCpHbsCqt5oLIsYfwej0Q6STFiL3RwNrHmAVFBi/N33JXD1sBb2tcttstcQf
zbplSF2GVCEPixrYtm4D0qdPl0R0KQgnU1nzu7TptllveiFTk9jDDhqvKtKP
C7iJVAS/wHvq1oG8PgChwXCs+A2woeWH3z+sG8fck69vEsLllP6L0tf68b2X
0//3dEQqzgUzCA3Y0PzK5rQPyekJf98y5vxLD0RidzXrQpU65jsO7ovMSZ9t
zi6BG3fkaeI24yRXgwPfqjKXuK/QzbJ76Y2s3o9sZtL6bZsWGKrl9dLLUKfk
uSp0CEyioxxaGuNFQooEN4WOCoNbAanzm1s/Tt8j3qXnM2j43HlxlK0RYO47
USeSVLWK5vgS50U2zWkpA6xSK52+PmfgN5Dci8t3J54xYxNCm5Fv5Vi4+rKM
iHSREBRSHip9Tpf8CmEZDOg5wzyd4qW7WlSctdv8qFPtgWKSPbU1Bea0mbG6
XMfu4bmLACYlBGWwK3fgxBufU31gyDW25ihHab1vS1COT5DMPfROx7dCSv+6
IMAaorv2pCrmv7g+Ua9EAs9svUYha56Ztf3RWIpcAaXoz4brsJtWDM5sBUCz
95+VHqDsH4UM3Six3qEZvJAELrHRYX3Gjzzo9tERMIIbFso6wcta9NFkn9B8
RPExWNVh/DioTYiQx7HvSEkjy6WHfP2k2llP2fen2rVRapIyen4phJlx+Cym
qKhRv5zgUAzigLGKHMPMqJFqjRVBycKVyPCHTAxn4zm0MeTy1us0s6MhVAWh
HMIxiPQzwmp1Cc2Vim1i5nFpqFRNJ/Jvdf6STR6UYWCZ3zWbYHayTgyN8a+G
9lgOeNz8IEuPH0b/2zIEP7vJXyRTFJz4tauiXkMlLKP+tI+Bqxz9wl3gcnuk
773Kz75U2upX7OGYuWN4Ma5rvwcQ2aPGi7c4RNVaywlW8z75vxcHTs79mpvL
m72Vjp9ZDl/yHYAz652gxoQQomBT9PiGjPaAFern3MFCv6uKu2s1KRIWtyye
R0AiZl90MPqSB+aAueu4VNTOdI5qKXKagHQUty7ED19uXh2/2OELrg1uQNeb
p1pwB9GzPsM7y3x8k9Tjk4OY2oNPWjUBmYwFrzwcH4d9mtT/7/ZNwYyejwe6
0hkpTDlBOjjmQeynX6+VQwPmP5uOuTyiNavjntKbOVPBeZ2ZyDrObUAu4TX6
IMwBxOfYAjObfSIZBbiGoOud8/UkuUNHb4aTWl9r8j2AIHx72k/xkuc2MWjz
Sk8A3ICOvwhXu7nwPgX6cosyHC14WE3q5vM6WvXRPj6Hvzo8uuP8mMePTDje
YXefcaJGISRSn5rPGyVVsJ5AuPHb47NA0qDy+c846/r/Kt+3Lt/rPUxM1kyt
rmYBhCwou2NCAaZzo9rgHo9Cy1mpRSTOAGq8+CKNaEjBmNguoGEoGYbtmx4j
6LSZyjJNyrLzpEGqXxzB9ZRSmUf7CqkSb6Rx3zat20foKbkAZwt0PNVotr8c
2icTL3ttId2L6yS7vRfaFYoSypkdvt00qS60eGMbVxsrHGtNwo653y4seYXs
txa9i12IL+oIRWM/aWS7in+vrCZQK00pU78W9iZ3K20WRBE4in5huQ3PQRHo
Cik8QwIEjGHeVnwgIWtFVUiZWJcHZ2hJIKkdzHRpCeaeJLxhXYNTPx7uO4ua
J+v9ScKSNGy/IpU95iDX7Onii90kpj6yBj+DTMPzu57SQ8xErOLe8OFDvZhz
4ULDly7w6tsvdOo+HLTH+Gn+dMdvykFF75hWP5r+HnnOlbO3oo7eroilqPSR
M5Kc2R1BRlqr4OlifFBkTmLdKnJpg+GEBMz4Kc//ZtfLMAhWEghFDyCmtNho
hnjfipuddc3gYZvW9193kKYeev9VBOK0A6m05RX7v7qJfkmklBNCzuChnlUM
9Teck+euncUtmupepy6/DfXP533DLSMwPKaESsCpGFObE6vIevks/kDz4Llq
f1ZE9oYjyhQ2TvJ2ZIMKxc66Qoh91o2etYYfhM2vAkVJzljC5jNBSPstDU9J
ADHyl9f6Y2h6Ydpc2GSCBdEnqj0MDscmE0SyZ/d0gewYlWgppEFQzzd//jaE
Ifvr00VmD9rTOB2kx3fNokClrPjMHRtH3//SlKBrg5gBseksOXFzGliLJl5I
TjLHwAuKUjIo4lUFF2wj1Vf7TyNDoZdb9Pyxe37UDGJguC2Tkf0vhqLx2Nz4
l0ZSHRToKxkgoyi3Gji+jqQVifpY35wflLsmKIzKN5M/ENi9MN1JJ8dz7H6M
XUohZ/pyEZiOkLjqcCDxY47J9O7GkK4efieOeN2MpITYZCQHkJxVzrRAhhqD
OpmsnjLtQTjCWLQG+Ir7FjDhuf6KiX3bgynv0vzWwXlQoAeT83us6QvA9ZqN
9TnL5aAogKXTzs1bmQUU0rsHFTgHpTZm+5CB/WFbVm+iM2ADA0iKR+UMNDar
lZ+j1ytnLh7CvFrF6hzkLDn+wi7up3U0KyGui1GFM5zDTOJ1VFBrvykmBFS2
dGV1X0YLPKRmcUhswQmbZoZln8HvRoywj4GIW6BIBn7soBPNgyXPszG2Agi7
5L/zu2lnkYe+WmY3Ge5Hx4803o0Jii3YUrBnO4se/5iSXyGQqxekoXlD+K7/
keEhaQXyMOcwl2kRJM3Ts2kffmnCyA8xC08xX0Aqnnjg25FfE7k4iIo85thk
gzln1HzjoTfGh5n+TW7o0UDVLcZ9WKQsl7z6vBoI31EvikoQtKGbXVwQlLOe
LwaurEtnXvyFLlvLf193aCEFIg7rSAkg5ZiikCbOM7ZALnSNH5OCcLsgnA1b
PrR8nPI0Y4CtC5LrAXbzfYXk20YN8Kgw0Ep/udl1WTzQ1b6vRnegBfot0CU/
Lmk6lR1fS2ZUq/LK4yJQEWEUUDGFPZCcGnLlzBrFMc3YsFxFHQHHeQN2Skp4
cEMuTUDAQg0q1lV7gRHMhtgzNDRVukokkDA+MhDY/qxEx+RSeZjLNzAPVtcl
NBws7pmaRRPKEJtvT1eYGo7HdAKvtUpDsONnxIKsNdkXV9m046GtWo5wbHIM
YrGzjSgMyoOvRh3OetafTnY8h1ehp2VBzUmDm568EyfoVz/4GNvoO7rDiotp
01yhCxSBNQYIYeDMFu/8bg+ucNNlWG9LE2XXqTPvYAeZ5nRxYSLcXRNu+lBk
YYRu2c57V2DuAS+8hOeRcXD+Z/THkyFMl9lERBMxGxt1ke7PdiCu3+77ewIx
PumAhXgwjY5lkc4UJHZFsfUbJz/m2NTRxHf0Vp/9u9QwTuZTPEW/i188/pt3
dPgTAznO+pNa1hL6fjmDTrZGBptUFmcomrwrK372UxIU7AVoHLMiF+erPTT2
qB47/WtH9UdThgkN0ZX21EUtx23YWA69hav0hrjanxvtwzwiLMeQl5wFUrKv
GmlkJOWbP5PVBh9OSNTPT/auTrkUqNet0B2x82FlEfA+htOiAfeztc51FcN1
IMIPWvFjL/4ysDRZ+nCvilB4uhpm6gLvawBUZky9UIxK+HHvpCffOD0d55VV
Xehg4G7ZBHirnobn2HARqdOObCSBw/OJw1a1LOr1ba9kVujXvF0+Bh+KLyhu
ri92u3DXyh+JjVdKM15vCAMJwohED54/rOmcMV86p9wNzWLmieJc0+jdBaFm
vJBdPE83fc7wOsQa0eW0aJRPTximbQEcjb1f0iXfrDUA9QVUi2QGeYUynoLA
b1F3FEUtL3yLAsYucwlgqWLMZJXjQbIVTXwylH5KDvMeVGH1vCBUxXhZiwHA
mQV4L7d3sKBPJLQ6RUMBgiLZKfeYM2KnaVWhI0Q3IZRtZvesg0qTF1IJ/L2N
+hU7TReUO03h9EsJOXpnqbdgmZhpPuPYDE8j95CwIMK5w4qIgARJWCSlJ1Cf
ZvwaOWiF1hz3MegbvZ4dGTJo15QAQgDFZO1xz8/v4puxYC+nFJoHRuAGpznv
ifidGC00skF3/fmUNkkztH236wUvntyEzfpPul2pfOL1DyGI8SOEDUSDl6Mb
3LZ/l/JY9mzhv4J7kRm5mRp6JrmUKkbXZ6RweagN4iD75t6/yOOOmeh5BaUX
OviGlJcHRDK8S6WTMX3VJxdw5mB8w0EpjQNgpLWiSEMfplE9r7lV/ulIVZLh
TyiX1HxdpEqG/HaSbadnncr1oAf/kaznGKM+4Cwz2GHaHmFO397M0DVUmd/0
NdPRxQv+CM8+wPrmQo1vlyC0/GzRxNVbaRV4LWvYmP9Pk1JdpD+hx8aF58jA
QQP2+3NR/W5qEcO97UssD74cR6OA4T6tTKYPebIZr1+Dsq2uxINeo3FV9CJD
S2I5NiLfa1Ub0IKcRTzNiNDgzZzApW8GMn7hRQb3h0ku2w8+Fr5osZbS3pUI
O0kPSOoxgToW+j4YndPFwBCQgHqx6OFxnvL5SkJUKQHs+ejGVETWvQV0nH/y
EgZU9jvY065FuIbofqK023I0MCdEO0v1lu0oj/YtzZ3eRG35gBSB6QrqLRVX
qTQgtZModgBIZ5B2K3V3C4AyVR76CK8qHvAjyD1V5l0DDv5dhP8C04F4MITw
k8KQQu/QTC/Ew52LwjiKEELpiksL46NWf51Ed0mm0Xh2j/FhvHMMOjHsjGfb
+K16VEHDaBVITFYDizxa7Ga4kaZcuZDIhJ4G9gDpweieRmNFmEKiO6EMGQSY
yfH6SLnaHS7g1kz+p/6m4pkvBSDavQc4iPyoRVRVKD40V+vnl7V9eX2b4gWa
Kn+Z6LmJ3ITClHRo79S4ZA3Pawzo1VN+0o0UBiahU09iSInfdwVG0FgbUBhz
Xn/GosaQxf+4IfCtRYlpAF4Xug7uC/qt8UjnMtpp1SbvhxGLIDDDUEDp9zCn
AUG2fwWexABx2LfPOkyvCs31S19Q4km1dxtP+/oaDxm4lY23ogIbQL3VlVH1
kv/naIR1CyWPeYVIudPzUZbu+0WfPmYNQGL7bK4Ob003gn4Ohregc3TzaFhQ
dU+Nayj6n1H6CenEWx+1CfONBVaeTsk2/6XbAvun5bmzevgQPx1FY197TrzW
/4W5BQF+aOXN35/MlrRrdsizBAHfZnVPTtl9je+YDnxTJYuP7GSwaNCOTUuu
WwgGWIUgV7Eo+F8arem42NnHBkNgzVaFS0blF6/gcO08/IC3ocbRh5ghdkW+
F6sErHGNtN2+5WOINY/vEcvtcaQ1Ktdcy01+vPijQHespXadNQvuZwhRZ7x7
BR6ZUqCUzARhu4IKHmQxWisShwHQckeQjQMtCjMHvhn2aGdaCaz3Vrw1Z/n3
Gv2XvmsqlBm8jo80CNhyisRJghFSWodl5iUoyaKIYN3dOQnJqmaT4RbzozzN
aZIU8SWJ4i8fQfyGt2Wslwwvp5m54e5+bSr0k31NVQvdgfDw1/+vcjwHw6ux
0lniEF7DhQMZAbls8IBu5aDjZHkEoD/Mv4+Ny4K+eVt/EzyWG35l2cVJ89Rf
MI1d0jTuP1a+0TQ16klPGqSRBS5om4wS3JcvibjksNxJl4H439EhO+DR9BJJ
MCnA+toDjt1oIkJCRZSeXKCRwwt+pFqshfitiDWqWDy3xiRa75jlDwPeQFaB
ZrweqA+Opn3nJIJEhgy15yfMHyOfW/nCJwCyqSOsz55+ZhmWICUAO0YsnLaZ
PrzbWmPr2V0DSoMwchiKwDGI7JE9nSFxOlZXk4QIFnbRZ62gxJv+Xbv6nQh4
eqD14nnGAgctJcwjmQxzQeAyGjnoxsALeuSXcD78mcsfRBRPOntrWMCDYZ2g
lhLgi24Nrz4XVzjjn8t7YbQwHAuRbkceWARGKZMAdMa/kN8scFy2CG/kRrEz
h7AYuKk79zh09cnyrGfsKExPStW4fFfYXue93bM0ujqhofzgtt53Z3fmOCH3
821tYU6myoW6kHj60CUJ8cQHjyxOM5Mpo8vQcRAQ7AmC+oMo6khcvunZkp96
X+qQ2vMSh7P8wAMDg0FosicPrSoyW+qjoAS3f83+Efp9HbaxBBA9E4UG1oMZ
l9/jatzEpp/d5k/axACReyMIKtI8BJqtGRXb2jG2KB+EtoBMxv2i7BMQ08sm
36wATS48/uzRopb0WFboZ/zyEdT4Y7cMVaFJuH5UWDd4YysC36gIBjV4Dlfp
HtoaJssdGegv/Cuo5GG1cJYXwNjeFulA4U2un1Dz8kGk/Qv39a95wkP6uBZW
GBHumYBFep/9mbUe8D+VfbqD1Hr02yMAmfzTdhXgeJqRNPqetk+S5U17XexD
4/0mf4EAup/it9L4na8oyA60HnEoIjD+ORa5y3J0OAop4DkH63MiXtArBPsQ
UvgZL9O224176h6rCuMRRlwT/KuBS79gEx/tdDRvC7WugyCoiQb0Ogtyi4Yv
V04EhvR3XKqI1Nkp6SVG2/LcMmXobczQ6yiZM2iEypR+TQ11yUf+DKBynzCN
aL1+hrQFLuwMhwGgKnd0o34b8EgXTCRGhnUejipWzu21wMkUrdbHFZs+9CfA
nZzLrlUDRYBCXxSC9MQKx5xEUv3rG6iSS+KNl81W03VvM1xlab0iyfreaHyJ
/TkEot92xwBlVqNAvbEs5oApWn/AbWEBT9ROLYorQN6/BUSHDISQJGKa/xCP
UVJ8FWRYWx5F02eCec6qWfiqk+CAXxO9mJgRVlKMR6zSD8sPwYTV1l/ksOP+
l/54CIqDizAWjU2roZYAY6lbqoikQyxGOlbmJCAmKXiV1zgygG6YZB92wd23
droKPNcJA2dXwlo3ofdWjQ+V6XcbXuoAg1O4/4+MFt+yYFqERY3YalTo+Tmn
R5Qlqnhu15L8Id12YfOkPIT7f2XeaB4RxSN+aLL86IRbaepm/zI/D/2tNEfi
SJQ9K0rYdxdfsSJovwbcULyP+6cqcu8N5OrprR45ZjKu/4GhNAYwqLhBK1Un
geYLIE0h+vuvM2Aaw9eIrt8Znmo7KWA3Pr8YNAYcoDNFhYbhfMb10AxMTncK
ECB3AxXKTydo5br9AAoWRn1shPYW8YhnwXI5edO5ZdgUQDBGDRKdEQ4ooHva
XTp7ymUgxbN4LEQlWSq7xuVf2sHV1juWoOUp4fbq0mSzU4ARodJtXQ+EB9S6
hKC9fGmCMmKFS9Ri65cKR3PN1pjys2zkhB518qc2HWbTH6aYI4oZsrT+w9uz
s0Mhk0wmULx5MqS0LgRiqLCvDanfLPKqwvH2J4rls4x8Gn7F86cotoXNdS3L
48rOH+av0vblwJU9q8WKxTFbYLSETv/XbdfCm9ZjJcKu/BsqYO791tHJE/di
Exff5XPT5zoI4+9J5C5qwLE2ELzmRZ99P9kbFieOiBO2xex9lcSut8wjOb6E
wiKuV43pdQfZ8kgIujKOfuQQ+RhRksvs89WgUrCKoIzy5mHWvq+A95SpO0YQ
0v+y9bkspvxTFK+bSWvutGhRhOobkY2QJLlNglJ3y9vpvOakdaKRLIgxAdJG
k3wO2iUJtTSZnpNJRXnPdo7JwO9ujIdrT2RfMRmctj5dtwgF5et0LpVgt1EQ
TJEesMeet4xMlihwmY8SLQCQp6KhIHNOSUzmDUzuZM8fQ8urmhctH1tVAkyZ
yKvlq0JBKXEwTbbZOFAs7x8DjRaV8uxZYjYhx3p2BgkeYBA4LRQcbja0k3TK
fn4HFmZGH1H9Yhh3Zuf7S9/ttqdwoovjvDpAQgLlwBx2f3g2fxOQl/nA7w3n
dMSZz/NiMPaMt2KLHGxzHToYaNlPqn3nYvKXmaEgKJBG3gmmtjNsixJr1Llg
NwXyuiULU9oltwwoL3jKUBptsO/DTV45eZhfHymQEO4Ts/Mg/UI+G9G1rx+M
vlwe22K8hIyrLaB3wZL+yKQKN/ZhuMVvWswz7uda+rcdj8n/upFO8Kkyt5jB
nTCevTyEvGaWw5WXxOiG6HS5SMI6RlrlXGLf1qxav5RIOvgRQNWyQwqoHyiU
uhapsmvm5RBIewZPjHDdILVMh90iGB1iZQ2qWPT6Yc4Jovhq4o+Mv6K3ka1M
uMCFm6IzlsrEi/g6J0WhB3zQxo/ZyY5WEyLFURwbVORbs5kd9nb7oFo5fV7r
ONwztqxr53mikDgF8oaXMeQIn2FU95Y3rgGkuEIw+Dn7745+u2ezsRn/3yPe
aRWLdzLBg4Ae665es4zJtih8QfhNlX0hI10lONiGMB9PycYwykZ+ad8EPA7k
qMzGXrg/7CLs1VU0p9rqeq/0K15kAo9SnY/7n7nde1qWU+fM2PpiTd56Ap6O
/yfk657NzQ0UCZUPdd9ox/CNw4RaDf4cSEtLijn/wMFeGqCTrQOFCp2tfmTq
q+whHoNyFsFu8ScujCN2juKbkXHwVqlY0jDmddpxJEIDdw6S6v+fhaS5Tp79
32rg9x4V+UzD7dOL33SAb4wvUtT0E/gWW8tRbKbdgvnJUI9//tIqtIK1leeR
GK85TQkuMNJvgyoeOxt9WRPxAoqBhGvg2fKmKbL93AAHQs+xdqhNRgBjesG6
zVAJrgLz2GWKYU6eBI9jr5s3NROD1XvBTsj7h45ehjyGIGM1MHzDPRjdfQQO
OQP61bNoplUyhN0oDYZCbjORhoC9yv2IxNK7yxD/z1wM6ehmMcPEaSDdma6w
7AeWvQaT40ptZ066+X1hRxfLi+T+MV92s+ieh4Ku7C7sqFXJb9T09vEgwtUM
YN5BehMlT0DC/6CPieYK/u19+fYSiQW7VPY0o/ZrWELSA+Cnok7ahT97rpNW
cIdD3jVq7z51+CRGC0s81i58LZu2ud6hZOUs5qPuWLprKv1Ahf3Q3wtiTc0Z
4km2o8v0QnE1yPTbisRTIQhh0yk4YGisVahu/vshkVMj0zCAk87JZ8e4j9IM
cP6OHl/ODbVK5fwKDYDgnK0TGHI/EKDr3TQ9vWWMa2oWYCodVlU0x6VIHKPs
Ha4wzai4tMic65BcD6rGcXSBoGaGTt7UDEzs4IxevZGtn08Q1QnNaZjEw2/d
e4aIc3BUrxH1+xk/SUZDzkBb377/CV5yk1xCpV570NbScOSZBCrn2olQ/FQm
xPmJE3ma7WCD/OVSzmjxDBgfboZQL06pciBEwYFPWWADxjyCPXZMFHSqNvaN
KxKdcInOAJYa4WpIfBuBN6VNsj2rDrfjkOxJX8CaB0rYfwk5WA81EgCwCqwW
NhR7LCwGcLwBDMGtbWzzH4qSsda2YyAUcIeqhEpFuGPwcTwklCHgL3gAvWqO
jFmFAGjItZwDblvWW1KQ2sBnaU98+siuYQmQQpCeCRq7vhLu2ET4NCQUVEuj
OKJ6eY3Vs9OlQh2iHcevJuxTgGMhkyUa+zGY6IMTX2geYsSpu0bBSu4owRBl
zSTpOgr2h5lJb2/OOtJQ1wkBo3Jt41eB5GFyFFhRWP2XD873X+N/B/6q3E8l
/YyvcB4w1oRumBgSsj/KahyugDfRKv05SrZk8Q/bu1n9g/at67ml4zxDH7sf
d90ybAp+wrfserWq+eObHTyJo/O6LhcePMzLJbGvThO1jk7q1rHaR2IyKFON
tAM2MIBZv8a5acX8TT174Dxfph76tEgqY1uXbUUkh/Pj5y5mkTjAM4lqCAtf
yLh0TnEjf0bK4sqnNXI7P1C7Na5U6n2ifus6UHFAUabb3ugFETGg9cdbXdBY
+M1mLiYRxG4zbw1b3CTy90YV5XdoyIjEquuUmTySuWWCHJbdzGlgBLzndM+7
g1DnN6SzTpYcZZniJ+GNlJhOnkfdWICgnHdIOFwmoVHvengR6ZX7bL0z/jec
w6N+t8b3SjFh5woOYLLFLbgj78ZfZKR582DbdUL4VY3Tjy9kbsyZxw9dBKxI
L51TbrAPJZSmoXTf8zmNNf8JLqfk5+XYjlQprM2AdZxBkS6nhuIyS9O4UgKY
zI4XhyW9vmuu1xBnx/L0pT1BTwjMnqyY4QpvHrTzML0DZgif3x51FTwkGhBg
J/Y2QOpBOkeApbVruqpmMXzqzsiqKcGHysGL8f8coDExoBfv3TEjTWKdPcpI
+6xHl8nlEOBZuz7CvkV0Jg8EMzsV6sRvkP+YTk9Ef3kRXPZIjCs7rp8gxV5L
j9gRyBUJ1OSJcW0ACL9lmPIEXFWOuTCvuoiWEvdqfdasevs5X+XtREbKyTld
5TBaQYGycQPep46pVrMen3xPQ1GO/Ea1gWrI09gFE7NBNavcjS1555MfA4a+
9DZS+WInJhD/nHDDFcR1L5BEgruhalziVJOQf4+/0/5KOUYxIlm0//GJpDWO
LbNrg85m8aWShOClihpMfsU7VOvR6mGJ7K3tE6Oj+RW1O/TYwAMicO2lJu0w
Fup3vsDAGABNspJ6SHAlIKhi4QCsEtvjLkEU0zv14UYrTusHC+zJ4oXI8RaN
GOjHO/HOMPApnDGJBg84BHfO3G7034JujaM3KBVtTTXgXIhbHmmJKlFpwKc6
c9i4S3qZjKL3cgOSOtJNrcNkBllleDQ3aJksIKL+o6fHtmNTrOrF3fKNnIRf
870MSWeaxEg0svn8jYZ+QQdO6QnVNmonIa2M1dKroKTtbYErLxlHywvDz879
zyES3Jjeud4+ZPoThSb4AeB5+R7BTgL6jQwZZ1ghTjkzpsgRpqV0Czy9UBVt
8XePdECQxgw0Uqtx5cPerYeW3M94sCoAyv7pvNJxuavQeLAS+ND2R3G6vJql
HnTKnx0lNeR3MR1Pb+6UKtPOkgIJq8TXcX8EcZUI9JqT9wqBf0btpt6V/HBE
lv1eSNB5L79jYUH/F999WDLVVRzSbb5wC6LBntBQPKgQGq5hxQr8Wmu6/n8H
zZkTz51McHPScC7BQNk77Qcr6VfJKzm8NDA9qUHRv7y3WuNMDvtikbBs68ZV
y/qM+x4soHNiHhP6WbdZS5ZKNAQ5v/mSluD6NlUBA7yBAhjcHz4TBYJZkrbv
i/MULw72bc0CThjUwpjLJECGsbCvuRTEw1DsRRpE/Fo1jOPm2sUph8dbRdd3
G+nQTDK8qqk5VE+F3sPtH4MS6t8YlISbRWzquQUD1cxZA7L8kRhYYiAl6Ovu
hbjH4hwjREYElbsMom9HTtxxpg9dK8qAcrAKzDILGs6GlPLXbRD2IiwdtsRE
QSG0nCMLfx7WtwtPu2iKwTcLL/AHNlF74eeGoSl3OBgVaEBspEsinVFu8ec4
HfjJpL3cbfgwQ6Hn/MJi00ab0CUIjU54GWqr9cBTOfDX+3n+Kpz5lAH4LHZB
FkhBAImwSYpFjlhovCK7VirA6A0lQfku5itExfEQiXGWmPpoFlmkgdyYYSQg
m0OHR+7sNN8ZLStv0qUNYsLvnWq8JGM5oONl6UmQDkgH5NyKr3hRniSOXLbf
ne1KhjG8lYek+90VbT4Wvak686DL79puyItOiUz1jpEi3qJQWUcombbge4jB
xoMfOxlXd8jOnAb7YYLdf8YuQk8t3RjMJFgADtEqk5X8+AwvDMh5VmsEF0wm
TRNo5nChFj/STj+X4YCDFagj/HZiWiKw0t0t2TghfVqdJk+GyQCMQiKii13W
IP2u0mY3BOJV30sVkBEEsgxBq80E6JmyfqhvrPnaFXjjh5w+W8i+17cnoAxH
daCRfl2WjMXkdNuTiZeXMqCzlS7tkiKwaViq9uBqoJLVYpeu5xJ4tHmFFErb
qf+WK4ll38hzjMGgV0UcAIB5cDsovSP75902T9Tm0ZOH2HrdtvzONnIP5MKu
U/10YMjPcn08RHd0J7/3eJqByfj+dbQ7KJ14WWRL+naupvpMxvfEglqhGHgP
kmIYbNtpzdHE7RCEfqNWMaw/soioEH6uxP3uyyS3FrkA/N39jMem03QN8pgm
FQoOA2N6j4jT82w3SyY/7ERW93xj+cr9WLpWm72L/RrDA8YY8R5nOvqgT0Yh
cT55R58WAtuNjHe3AOksCnyt9Gnf+MangM2NK/w+cHGKNPImloMMQNA6zjvi
tskAScyCZYKXHQCcbqawLX0m8CsSqH8Z7dnmA3L0vmaS6M36oCQP/yN4g/O8
YYnjbtlgljZag9JcMSMMSyvPsShGvd1gwMftlp+xfB9sChh/AEMvAIyutdSw
kJT7amBCXLYiAhi//Tvad2kNmB22A1RTBopBk/qTiiwk80Sx6BBQOZruAnVW
hEMMz5zXE01ziJcImrgcCjOC9BwzdJThSjj3kSkmNICRbD8TofGbAx9298JH
OXaSlZKax3Oefydvtr/b1/a/DlGfYhqV3V37UbItGWJppzIxjz8uDkKBpHT3
Xp1ZVG5j6EqSV8Dj4ZtXDSvYyfeVzPuOUwZ4b+K06ty+mMXWVFabp61jDyXi
R/LLGYNgxo+5Tt3kk6pfxDndOOa61ImnUjxnzkHCPQlAx56Cr6GfppoEbN1Q
RcCRU4R28xzhfLc20k5svuysVIz4l9rsTYTyEy5OU6YXR2IsOzYziStEBYCz
UoSRHc1Vtnju+ihOEf7czFDTQAoVOwcBstzLqh3PWt4vVQtLu9S/Eyk9DuTQ
r6nsnwq99eGbZRBDWvbMBGizoZVpmR6PGr50QNqqTXrGwnRIugX7V4+JkB2O
p2ARYOPeJnmXmyWApiQPLgC7O6Nc3wNQMTzDH4b+rYVm/Q3bfu2MYAShwWSH
JZq9vA2pSD7EkNb6Md76dABSIrk1S8f3ai/UwPV08o4pYXdTcl5rwGTU7C/y
aS1sZJZRsEoUjw31IIzeTGbj9CfbMxoWS6DkghHpXdX+lTXZigc84RTbq9tS
NdSN3rfJM4NBIEa9zsyhcjXe573ddIY/BPy9O9uCbF005V4x8G2BkL2+f0GY
mCmo3756Rz+rOXqKExZPGz4EKkXxTqnjRR/zWXCl8N1zNimaw6F0gJmTQCAg
5BHxx/OFKTbXqFGiHJLfbX4IeLdDpvnx4Qv53eATnwpEAUsFWkIrRAawN25i
AU8ib9PHYUC+8kQXbBxxthLFkACz+xGsvxUhOeUSkkFa/laLmFqmxXCf9W+P
vQoCE/c8iUVU1a3j/ZxFcQtaZOForb4cpcr//2EaOdH4v7DerP+MFAMPm1IZ
Qyz+0kntFmdpJ3ds02gMeUHSILkaqCu22ZXgSrQRxh7+NdCv7JlFXU/2HtBe
WJmDHrplR9nU8cTUMyHBtu8ecTRnNs3aDGMF3tprG1in819mDLyFUsijapI1
mjxQMM+UcHX8kiShtyKi1+yrmeampT0votzQA42lZCdK9xHlC0eurgSlnQc6
eRlVdFaiqVUDwpffHvUllZCW/meTAG/oahqOPdWWHp/ItgTJjFGmltzWxk4H
A0b0aBeWxsl3f+PCkEsEALC2oD0vD3DvS2Xvc7YZzbtWO6Gkjn3sABul82rJ
92NpduwO1ZZ2stJcEc9mZOaavbyA6ioWcpui7Hj3wouSQyH4whUG/MEH6dNt
AyYqRH8Ga05jw4oOvHd8qHaOKBY4fAv2XoPpvIb+Kd8aN5y0vgfjyJknxkgg
ETrq52fHrWIcbn/X6pATk+Et6nTkn6nwfT1Lm2cpbF0kppGNYvXIGBGmZAPg
o1ro8RJuT0jnhKCr2Fj1kj7ns7IILW8GQlrfn+vuScRotwJiiqLfflClvjb2
TyU74eKtcmhzu63Hu+o9dzWlS//s9yV2Qq26PfwUiJazsM0CPdLREXnu4nAF
lxJMOaIoY4dkOcDXYGJr4s7vrPxOwp/ZMofdyWRAEnSXm682PRrZtEHaVn+k
grrHtc9N04sW6TKhi77BltmcL5+WYCc+QfhxUvTjuae6mvRpA+9uMhzYrVW8
Gy+fGueM6byrhqncep+DWnWMK61NQPKZvQKiFVHUwwb1MU2Ab2jxCXXE8b/R
fh12TJ0+DMrMm7ZFSg/bO95i/u0PR0MLKsfBN49gBputRV82Ryz1OS21fjv8
RcfwoILwJU66rk0l1K3oHqHbVwss/b57J0yJ7lMi6RaOOJqxL3cpMQJbXRY3
b8s7kVMrsBG5IKhwXLXp5jNqwMsLqZK7xOWmj2q7wUcvXG9cTOl9Cww8j1qx
HBy1WS+xnpFxN1xXfsMoOHZVZhmQ67QQcb36Jg3pGXkxjWTZbKefY7hAOD0+
wTHeAyXIasA6MqtgWQ6Mjv6wyH4O+xz3HwUQQfeXBcax0LfjDZFrgtElma4y
gcLZzVPqGK7PEhcGmTI2Q3IbFBQ2PijMN4ik8xkIshmjo9yn8/PPtEYiZRkd
os4xANK/2NWQIma7TOmRncsw5dxBtEjVofevI9HvWf8vfrBhRoR095Tw6O7Y
ygQgYcO6DrudmJdCKo8PdTIGRS2h2XgmnvEdAzls7ZweALpm++wPhNjImB+y
506E1y8ch8FarCNDQtNjmLzAl+UKopgVbt2SaxT1INHFI1zjuZKxa07ozO58
dlCN8tcjGQKQecqmX+xWg5R0tYUPnlgHbn+7S7WrodzrbEFU8s76xVLHWGPd
1WeZd/M9neuXOgH7ichxTf7X9E4HqZV9CMumP8PffGspsbqRpM6xljvW8ZN+
e+8qDVBolhrxMxCrCE60zvYsgVkv4WDATUsKKGkpfUWT61bHV7GxJZl4VW9I
abEnZOpmiZyXw3qdO9YiEnBO8Am8Y6rBa7rEPVx+CPStg1Ce9n5sYfWXjzA3
+V367uwpLbolYOlACf4yAjEJ9Ewm0/JXDgoBS4N+soSrROr/tvkNdd/ohlME
BPGi7ILpHxalwbzSeEn5xZeL2sFBdjw3ObLpuLVWmG0NcslZxbjsAGXHFYmV
mQJQqJfldi2wNP64B4iDE668JTYI6gVWJdHPbAb0DvSYK2wSyRNM7WmHv69h
r/BErbZGzosZM5Hn9Pu3PNwCYpgbXnD+6Uhz4uwwd/tHPCoxiw0XU66J4Eo7
Q4R8NwpEAKt3uHyJOoqvbY4v1aeSPuCvQ9KwXdaxyZTpKwVSCgtbQ5trQ1k7
2nx6KvNDTjKkT1MNniWb4Ww+yk2/7n8iXv6OldQ85/DSLmDY40fRuDbSY9xV
4LiA81AWlCeN7KqGhn1oElAS852FaW0pa6FbuENkEO9UQiCbjfip+YOodrm5
D0VSbmIyFLIcHNlig7MZsY5cKjY7OtHLCNP6/ZxvmhP2QyqCIMJhpYZuJI6q
HrcgTpmWXTlC7xnlXpq2TYUvU6Wg5umdBizfUtmFknCIgxzFjtQ04uMiIdsW
HM5tx8wpfUtWcFJRn6vFxPOvPn6or8mpvKL/IESZvvZZXXH/wVv8doyg4bPw
w9yPvVTA9T6V9U2/176SK0CEaZuWERhU7b9nkmvcEUF3BKTONRdPQ1tC18xX
4GtX/fDTxRmx0V0j2t77lqk9Az3iK3hpDiVOt9LS/VMEpJzEDnJ9731PilH9
QVjpsb/wBmjRvizgzrSiVZbhAPUeQCnPZ15vnL/gn2wmE5Z7g9AX3n4OWA1r
1zahA2ZaIG+XvMJH6IjA/KDTYfYHYo7UY857tiZwmnT9zsGm/P5dkbcX3klg
yKCMN5Gtx0IgftdOd6uie1ybf4XAhVb/nanhj1KHHWK7ZDLvssTD8dJ36oNr
kyUmyq2Y2F9f94t57UH1EkkROj21xxiAPe0it54H/N3jnHZyC//jHp6pV17w
jp07AT8cjmsyOfDRkqS99yZF1Yzy4ebQANEHP0XHyf9wkMPjGl0R/KWQsAmA
udV0VsWQnHcdjmgoNiIiipu4V2Ru/OrfSFw5USaam8WPnooY3HT7yrCTVxm8
athlN8J717k7NOoTnAdowJfbq9usx38fzEHPnrb4+Wv0PpuE1n5XitRRHnl/
8+ji5avyaSp3LAmzNYANURqov9J8tpfWtIMrEOhWLI41Trs5Lnm8jbaXiamC
U+Jw3wza+1lKQ/G65rECZEufR3t04Y5vlJgrHiwkG6GdPLGLm+tJs1mh8UA7
cB5U7ZPkcCjXYr5Ak1YkFzl80U6vYWa+BqFsd+0eE+jAQLcqee2fq3hw+fUF
6R06CKJm4NVUJwtnObfKOVQ+aMp5q/TeObmPQHmowx7NrCGTiNfeOT6y74OQ
qwbZW/ezsOCpyIGAaw3JRN2vjBvl5H3sbRyI8W0f1zqj4Sao72uOYCG7+U7i
yHpoIg4tzq3SB0SNt4Gpfkibv6RG1vyHM1LuHHhXDuOR9v6koQ9igsXRnU96
E63y4/4CasmLCuAE9o0UsawgLXd2bOE23VC0MfdXHQ4cQiTFlYC5XA3cu1MV
TfKgUIMx1Eg5jx1QTcEoHOwPa1mM14mQkUmSvWFTfuXWbX+iXAqGXw+DcXgK
lAmg/bJWuN6LuAFXYg4wLJCZK0T+kyDhYe8qBy9E+b1kmO3FJyMwNcPsoQnT
rhXvUtDusTWiCmbN8O8KUJFmeCLtJaQRTVlF7AY0+kVs0BABzqJmHqmbGDk0
5cJat6OeHI7R4/3zaUBPCmqZ4EjD+Ji8h8GS6PqW8cyk5jFuQbGPHOA8zKEQ
UPE7RPQXPEB8etFMDOpwZieniaRKfGF7V6ieWErOw+XLliOtuVLGejso0b/U
fibCgMZo3yGTklvt4rcvQdL16KoY76t+kb8Oz8nTz+vJHIGH7oBeJ2XBLKRl
GGyz/XYuQ9I01GUpxBAP0x0ahCtNaNdHvbF7whIfq7WVQfXb2bUbhGMIYlu0
YTBWkfh04sQnk9dkwvSj+QqF8K6RRQendSrjLs3P4U7qzZwDwtZtgYIE39pO
FjS4E7za4mb42ozhUA4Qgcc2KxLzdc2ucd/L1YxiUSw8vi2iih+TQMZr5ueE
ey1F6ahz5RE5H0nabkhMyrM7Vgp7oaj77UNpuMh8tcu5YipIe3etjXv5FfZV
xtv1LZpcSyWlYsuM5n9deHbDHaV6hhDXKnviL92jo7Bq3QSLlrIBgo5q8lAP
VVzAvkNUhAk9Jqleneh32U6vnwhBFs5GEvxU2UoNzsTtqI9ckLa10nrGFsnv
Tl0cFQpsPDV1vGCG1AFp8hmE8pzf+Ra3wwoeqSd695GdZ26M7da/NEO1cN0h
rXmAppTrSIbPQOEMupvNLBYuOz5y0MumM3FTwvKAf8tGp3hFpRzNJrEslhKh
AOJixnaQ6E7RyQVwfTPbdEfjIhWpG0XIJmkZvFoCM1mdvJgQpKrMiIAVbRPV
/vxqpiq9hiJpFW50FZLmj1MGtsHMxMmFM/Swl05O2Kvaq8o8v1n0tTnGYxlU
H5qr0XNRiEs40QnRx1n6hh0PBUee+S0cSB7V37TyoskfBF05ECo31IXKh1kn
ydPpiwsa1UsEYC1lhUysEueVjbRzk2ka4/S4C4ZLq0B357amchgqRupcP7FC
T2egYIPdXR5zYrQCUoRJyfQFKvMdw/OHHW+7k+jfh68yc64AFkVGXlYJD1h2
ZkGHAkOibZXmIhxX7xYdiS0ppoMogMqaCIaMxMfEjKitaGsQtySRUmGrgzDv
8o53vOjB6roW9B48USCZqqGNJ44musqaLnV+9EQVOze7uUOuG46cVyQr9b1+
qk4+EiqSynioZiqmX+way1TtxMjVGsTbpgMFsH/AzqNmfrVXFCi3nayze5tx
xs/QBpKhSp4rbLBxXbYBo469AOBK2RvK2Avckrkf8L3QpAn6SYGnbIEkUcI5
bAmnDKLoSmqlSpGAoCy/AT/vLlgKzMzHoEIsFT375X+wgHyTnxgK5ho7SW/i
V6ePn5QgWXVvckKUYGNHL0HFxz2LhQGNndZ+ixjrLLPtO47EtsjShwAS41x0
L6jcG5IyklzRVoRz2l33HgyuOHPZpoSv7g4fOUJ7mK2ljumALyY3Pr4ggrvY
913P+Dyho/uiS5BX8h435lWB6T1y1mY7zV2CZvlsFDdCkpNcwA8j2mBdipKs
FLmjVYk+3LOXrr4tVS+wIZZPhuNKooAa32v7udV5VG/ur05KYbPfnnvrIXpu
LnBB876vY4jdUBwXIjQLxIgR8RvkHoZhdBp3w2g09g2uOU081SdeDnR+jTrS
WD+51amT75A+aUA1vm2QCaRoRdSbzSXHAc2oR0SNawyLNhid8SsijhT64HRu
RU465CECCht2qFsOdPuJDSd5Am9Z3LT699xIu00toPsho1xY0fsfHbOFqZHi
q6F2i+Bb5DJa0gkLBfySxTtDzs9AlX5/ViHmzqtCHjvlbEZEdqd09CziCKY1
lGcpOHkvMHVIzVrEsoOMl0rCrPUKoK7lZ2zquwz2hzwsUMaCS+YIQ41Bz1jv
HZQwdNy+Owf6Li3O3mhtE5dV2/2oj4s8PkUPqbwiaewAyJGUQYvUUw2/grEl
bpHGOu/wXSWYkyl8uf5O8R3l3egV7jEkA1VejI2jZ6FNLDBXs8NSc7wMtcV8
jXBRgYfsBFRRUP/Avb/bm0AGC8DvwVJyElhV1hENmaBzSg3o57GLVXdzeN9n
1C8em6xjDLt9v3CzKc0fAZMv2/CtgD7panfRcG1WjjOVF2iJ6Nicfmplu3Rx
9A3vKLWxspccGQm3s1jP7qRbuxCdgTtguwPOsJP+MQ/fV9bWGrrweL52eLDx
67ktEP+/Ss1+h3XclWBgu2T07Bq+bn+WmzlWaSAB/t6aFJ/+lIvl8eudV/Dq
fA45JFTGypDaxz7O0nLXVFBqYTD/gkAPRYTgccykBo0ojaonPVWbdwmLGBCH
0kckfgtso3Gg4j5AxdxnN4N4NC67NXdwfyumxAdqVWJqscuIEvLOVietXnY4
Nfht6vqoqrOw2EbozT94zGj13Rl8wROVpJx2eegbfnbx3apLGn+jf/GnLAt9
iGE0ZFzYM4ydtzGN3FDWciQc1nuVnB5NsD6D0lc5Zul2YHt12LmlR2aR6M80
EJ32fQV8o/WtqBpbZT6i1rEItPAv/aW9xC/bMBurecMVraANI5YRM6i6tCO6
NJiROj7h0Sr5JWlLnejVl4RfJ8WpfeleVZIh9YxIYvOdW7uGEdToujqp7PI4
ApL5ABQhpH80cQ6fRX03hYuJvKJDiFUFBUp6ZKLIO5qW4XTfPLSHQeABNGqs
/PCCnbOKHvjm31QubZ60/CCXWyhgk3x4LoE6Trmy/55X/6hYS4A487VejEme
rI0U3b2oj/ciJOmYH4i2D8vsbRnab6GQjqQXTPabtYKmdCKpHZtpfBo2bCDH
n4ddRktutDSqTdyJ1obGErvDDwYnS3OdeZ9NAwNr2j0xgakBp7RpM4io+VEO
RdK5ITnB2taKPqDx7+SUQFSNdgDgG6ZBchQCMsBe34udbG3pR+GA0FKumYiK
iILCd3033LZmSfGfbq63siv1SxjYZGU1vbJV9mhVEuCq7PB/1PXPcON8btTg
rtITzqmWUY4eM9xkSji3LxiNP4MJ7y07NiZN6tNTPczSNn8Hl9xWHvjV1rV7
z9v+dqQNvJ2sWNpuXgMAvk9iHTzxuoMzawXexvGI6cia43YZ9/QKXTXrJ/KX
64pakzHenLNnV8CtX5l2IYHOI9wyj+/g1uAR0aRpqdsavJYEc8QOAVtRQKTU
beATh+SVg64rB888C9ZXUEGjohiSDqyXT/Fc3GlDOg8VWokpLOLwNLLr6qTP
VKx3Se/P9gp/4Yj3lUIu3tv+xMqhHurmtYRJLlZQFS+txjPNuYoHgyAeBDuE
A+/IUq+2PCbjdBXCnDtwtPwNck7PM2zDo1GHD7uH2/9ibt2Nj7KYuUb/Ogfr
+Max9xdJ1LjvKlCbJrlK7RiCfSJPygEdvEj+hV10xxF5xefoNX/qO7ES5/9v
p/BrpTjzP/0o6L4F835kRk3ZprkqDwlm2h+SobFVYk4SuNdUSUkZACGcg+Pr
P3TdtEVVf5xreE/YcNfXq1P/QgYsMpS1rq3r0kgGneAkXYIR4eBeciGBBBtH
HRBV2BhjPxF4JIDi4qgt6oIqwgLbzCX6wFCJWRRcDdCiBVX/EInVzVMTgRbi
wE4/99qOpvK8FIrdBEE8eqds4M6VJuvp+QbcglL+LnHf4radsVNHdyVyd9o7
8DRODeHkhDcMob/jWnwn5rao6FFmGwOKwu5AQEhl7gWcYIR85ZQu2f3YUql7
Y0fJYBWsHANSwez245mA2UU019evG5PCI3WFS607wMzw26GaDvA1sGUy+Fr/
zsLaVmano8YV3DC4rdEobuyUsp3NG/79ZLJHTuWAVhLyZ5DVrTogipVtm2Vc
wOa54auhmcD3Yv9xseovUqhbm68yYUxSZehn02Nzu8cL0QMOjHrD49LNaSZw
1u2h/vxQhwJbbv7l/rQXNoXqTyf6TwL1lSr2Bd7NiGXzmi3qvTCMZ7KqYMf0
gOU7NR+8K55xs5oY3Hi5UY3r/jLkxnOKUDcCtoCV33TzsHFqp09Xru4EeJLG
U6h9Wi+FweffyNn7RkyCbqDkKDvMFFqnR+4nli0hmCKrlI9moe3Br3p0cQuW
VJ43nOmQcNiQnJItDLYhwoZ6omX9gNDfzofjSK9RyrE4SBzb6UFvLQxSZAWI
oRTEVeVcv0HwGoL7VmNkOYaojtRt4exKUWUcXHY9gnik3/38sSAHy5aUTnST
l5C+uKm76Ah/EL4ObqoIn1Y8btfAOIFFWkRwtayLKjrxnhosoI2328OeYXgu
3MhAtPtASSdHTbZZbniyI61rmtZp1z5iVp8whnaIlF35AtlnLxZHC4gThT9t
zgxkF8j6q3h5TrYjMaKgi+GPlbUeqbWRkjjQpIXGXQTXJ/PZsys0bqvPz1hY
E04mOyx48DQXL5GuWpIA81Ae4r17sCJFSHwxAa8FCbse+8naDm63zrwufoSF
QZpn23WmIQ6E+PARoi6iM+KLwlZsjOexRhovx4F4RNrXiuyEUaaFy/HOxJ/i
iFsq78b/kiSKh8srgkqrLchu+uvVjRezh09xclNIqY9w0C70bAR7OLmXYp1r
65b+TKfVaiI3r8DH+tvd302ZlLvhe+hqyzsZ70JIEBpEWx5G5qmJGhT190xS
NyT5BqV+VRR6sYzBn8bIImEwJsNmJy9EnPENhhMNUrEVe3qClwYv0Q0PzA82
HbblPksV++7tCGFgbCx4aPUu8wxxkneDJ69p61CJsTKYcEvsEbkAzwVTWdTz
rnrO0I0mH0VsGUfIMT/GkAXBoeMsmWMrY1H891MQgfGvUnt1gE5AKGOMG6Qf
tlF/WpwnQ7s6xEnGtzUpvZ6VmpsTOQYI5KVNxKb0YFCt25zaZDy8J29VZ7QU
zl7cHVl7t90Q2C+41I1J/QlFC/m5h8LWwfM8jAFMExRs8uat3uCXdk5Zken7
RzZ2cO0krckssRAlP4OSd0lrRiyI09be5xHTuk83GgihaTkB2puFgVUWIZ5N
3hVhNHDyoimCURUGVDz6xV2eYDNDp5LXXZ0mKeNipgBprZQ2HGMUzEfCDY2p
Coe17Lw3IKyleYhHtzJ1ojvCwbbAJt556awRyK2bMpZXdVN5h7kd7GX+v2gO
4ua/7mvb9YmFz9rpNWAJbNRjgUqeB4Y02toJ5EaFfh/pH8yyAGMngKJnqI7o
GGKZV9rbqTGPoay7uHxU30nrBYyCtsdBq1KM4Jja5g8PzqB2N2AWmod4Jl1l
xuRls6iCF9/U5HRPWqSDNBEb+nZZbU8UExoV3npJ1qvzb876woyOCqS+GTar
FPPSpm7nX2lWTqenOKFE1VLbIxngXXDyciXIDxZdc2WXwgVMJAghbhQLG0N1
qx6B1A7DVt7T+wBOZ5TfMfoaqTJlw80zPW1Uuw4j30gXQAA6n5EFmhYDYi7i
RvwmLyuIWLSYSGZBnyAL2d2H/uXM+7vAa84yYqbIDhowERE+fkAM4B9b5FOl
YeDQidWhipaEqf2nv7zheevS8JArxXVA14UDY6z61I7AElZgBhTu7jNPQc6g
KnYNJEGD3P4WIkGT4hgzUmst+5hUWVOdqnNONMKKK2RbDt6qKSxk0oVexaTQ
eDFOOkoerCDtTJuDsk8wgYafWbYi1hMN9pQM65W/8bxs6Kju8K9weJRPcgev
TGOWpRKjpuroikND5sZRInibXZ3A+juzafL+q2DWll9Uyg/iZ5caImjXpdpj
Y7uxPFMF4Iigj6AQp5lgKXM+6vAWeskTKsbs8dE71jp76bd0Z69fxSO+MPdC
ttXs87poY3oI0e5FGrOw84buj8qzJcu3sJNyREtE8j9XLyTN92gCKwi3EpAg
rzFtol3z39AL3xIgs1PIvlUUG5vrsEN4VUifAJ/WBqC5ll6cWrfF0N5OUrlw
GwAtxmLBUQcGOsRgCEXrRnqdIPAVbkjE2+/aVjNSxP2KjL+wDTo1VWp86Yv+
BWFZtuHT04wRNGWxnInH9neTGeJSmEh839yxxGqBYr+wfYTEq2rYn5QuWrNd
O4iNUovL65T6EAejlxlK6Q+1DKU7r/kv/IeL0xJsuGTPZZCmn4k17NiNSWZv
/aOZSrqmobiXn8Vev3PolxC1KP70h66In9Tj7AHG/9clgdDe6XZGocpU2H3S
u89wNwaOwD6p5Nr8sp5tq2GMKze8gQf2ZuKt4giMJPLoTTHjpw5y+tFZRQlh
jLVaKGboiZqAsf6T+Atmnda/TJjqpauIFrjkWO9Y8WH7OgMNRKktuvQ7MjkK
buXBN6MFE6ZDzj3NYw19ZkycfNNaUYihK0ALpY4PqXOmiQfTCT54Ugwv56Xq
OY7mWc6jUYTItee1u7AuIG5TwkrFRibYWsSUM24b467Aghk2ElOek98EFk6m
NuTf+CQKnK7eMfR5Cxi5Rmc+7RvQltl/Nb8BgVAq+OIWGmeOWutG//R5iNft
bNkCmiDNr5RFHeQmaHanYIVmAhBC/P7Im1UK08HLLb27nBF0RLV8NdwyYenw
nUVGXHNHnUifg1dRTpjqZooniRkiQRSO4rnZDilOCW7bU13A9aFu6qeZRVts
U5vCsHeES1Zy0E+SDi0CzTmwPiYeC0WONAc+jafqtUNrMmxmOtr483NrFnaB
wM4NHxSVhTAQ5MEJFCCg4BkVew+xisfavAo4TWouAThvvfZkWoklfOFvdoCa
C8/si1UotQaBZ1XOFXmi4ZH+WiNtodM6dp6uYGtVVxbDVJFJNBTALFdLkzDl
b2H34I4nzDdRPcuH2gmAlThxbNSqQU7N7NtqBFQproplJMfnQ/jmtSCqT4U+
VrsTdS/4ElJg84KInP2cpvQS2N2RgudoYiKQMhUWDcnyODb/Ii6IXOkwGzdm
L9i8hahq2OYEaTZACEnJCj2nObw6j69b+A5z1p3FBNSIua1o2TT4e/8i2QPw
2f/GAdBVStpjAalc5Fq6/D9/3h8bdH/csyfPDX7mYtKyU4XWKk4RMyPWs7gR
3fzzRqLSrcI2nmY1z8gDpOolsCh54ZLRa2tgCTQz61GWhw8PtSX+acIATALn
vaHKV/BSk18f4GK30K+0VvUtqEjSm1FF5QEf9HsXS8V7X8rOkn70VKjkmC6o
+JVcchOvI9dyO9tqZe2yxEyVI/rZcwKj2tMGQp5nvIpAIaZIM/JXYTGW9xL1
5Ocyxp6TBJ2R3XkxevQDpYcdj21bSe1wEPwEDvN6GlG24okp82JG4fMFzEfS
PLGIrPw7Z28tF86AsCJcwQT7bCAQaghqdLGSYu8d8VXvxApJrN+1lK3kHtYo
8lUp6tHRMzvGo+0kg0REQ64hX8Ov/XWDr8cICfjBS8qUxXPK9i0PfvYFk7Oz
OTSVaR5uoBp64c2MMvqGtI5T74TAwiio25+u8byHFHR7mr2Zgnpive6xIVmb
Y4ThJt0ysu457m8TVgRVkuewvoT6znpJ19jokVT/QDBzLbWD+pwTdSupSDhk
oXGJVRXo6SBwWurGtf5CvyqYjX/N1NjA565i6NN+JnAg3jT/b55qpqwhmOHz
4w4t3gnCyzS5Jc87zgnO+3qW049cAlVrSHz8+hM/4Vbe4gyD6M15u3I7iheq
tFudCHVk75lqbxkXuxx+O4+gT3FHXXQ5OXddSh66+XdH/0om3lHCgYZSWS6P
nF+iithYIBIOMPC/s9TukvlTBSnZrcJ81Mx/mYZEovVPlraiyG7D7Ut7RuLI
VuJjMk1+EsqmQ+dbdEdNL2zL9O2PAWenKgRF5LFqYPnhfL3V5KGBPCfmE2bJ
uoNTE2F0XRTL63bjzoFQS0urwP54xaN0q2JyZHPBG/Z32OFNvGyYDgctI06/
o0LeIdjqtxNlqhREA5jvSNMhul03jZJYM1ko8Fj4++LYCEdkFEpO82eoSsZ8
qIRPNOA3jYeHqAsFAnsAP4r57BjtylD5wr3Q4k4/VlEdsJ69Xz0oknxhE0se
wrFdFFV1iiNjJXQRL2DF8Rl1qLxdqai2QklHtS3F9GbcEmBNoywtz9pG8e1f
ppOom5UpepZBXcwjgqdifLVArWPD0KS4s/Tf20OENcWF+SdUFBa5p5ijZNRk
+P+WRE1a02EGHbhqbKgqTuE1qpiC+ApHArXOb88RlTReNxqVGINSK2wPgzXc
CaJFE7c6B3UhffnDM0PorOweuG2bx7jMAgy9QPNW448d4bWExrIJfTp5ZFFi
6Z+rCNH7qyv+aPGXYJFvoaNc0bVoezrj6ynBzIpEEXLChM4GSuc9lQrQkAaA
5pHSekmsUIRqLS8xMHIxPLEKF+scOElYLP+QZ4NcOTKDAsP65l7lgT4seprB
NTEFnws3UlKm9yiMtzbtmEkMnKjnJRjBCOePsjYhl4RK4bB3KsvIO5OwUdM0
UAu1RtkXpEogNhmzMU53yWZ3aNXqVDy2teYA7L9puZGe09j5aSHOLTKuL0qs
pOkk+a6XbqKa0sw9m/lIDUHduKmXAlq1WWNmlLvFGIFS64g1QUbx8vir43eY
1JSETmsv30GNWCQ9MwTGvh6aMudE/dVURU3AKSSoRLVtEgwlvQnUqA//fk4k
AvqMxHIV8hdyu/tOtC7rUgBEVfN14xfGOBPFTPLKLutw+5qDLe6xXro86LDE
aB4EQgtbEs4SKGi8ZT0Eoy0Bww09GWdhHxVjE8rlfwTxfQ4XUNmHRlSWrd11
1OW4nkP0JjULpDTryzYzo4+QIRIFtjTUIem3uTI5InV+vTVo1E/C5Am7dDQf
/483D85GVif5UAQDIVJXhNVQGkdDBmyEzhHDoWUmEZ5FgD7qghBdkx/eCA+2
j2lgNXaXmsPUxkzozwwjciszanW+R7VTKsBGKbIAAKv6jF21iXC6oe1b/y6V
eZrh+VrE6gP0M0C+stYIkuqAY2X7M1MsU2NvUUBa0uorTvFUcmbke+wqbwf5
7Pe7nQ9qaGfmMLStatgGDe6cbFMdo4L+gV3uv53AHQX9jRYH93tOM9gh6V78
otDqWWEDnMPt+MYZb2W1zEt30ZODVyFzMStnaAVH/QPj6dFlRiOP2XfqUw9X
k0gWsBp4K+UcW6vqyd1BDitOXhWbNULhJ4EzasI5dlP4G68i3hMw+49prDrU
fFnmTpsnHXlCRlOf+Qr4XEFPIdoX6HluxiiQVCTgmTcpOr17o7uLRRpkX7uQ
Z6yY3Rx1A079BgWvUVZKi9VSx2pXMMR9CJgaAEMzMTUhjmfWxeyxy5yQ0U5e
n+MAQYordK84SKceyMAGzKZdmSlT/JpnSWy30MivVWn4E3GsmSCl+FKqV7ep
tVuDwj59YiWvTJDg88j+hTho7lmXRTmlBllZgAa6D/d3RSXVohfae3YSGdh9
nb73ciucqqR+eit3flWLWBEpDuEaV76JlnVC0KfsDUGX7XubJewKBch5wQCk
SRb93vGcL8LS/cjz2ALM+JfFwQTRNKInRoPsMX6maAKKUTzF1CMP3PUKM3AA
Pti5vf3wuhIx7pXhmRC7fvYILPTzFFjFc1ynCZlr/hWwCVhrcM8pDNcisXPI
Q3Ix2HuMY7d7B9Uy9GCXLIqvAAwBkI4XWwcrkz2BzaUO2z1BaDjY0TdoR4e3
5VsS2rmYnb8WsB2Vcb3pCJ89x+BXVKHXynS9rjxH+2b3qQ2xmmkVL4V2MOuF
qXC8oNc6pc+inXPAEIOqsPqLi41QI1sqEtJrCoy59IHe+k6IYkJD44rc0qE+
ZHRskhpAIi7nsmCI/8iYjyxMVAFank0bjOhiQ7GARltADsUNghKWNgW+YdNt
Hen+YrrRIFsbA+DVkRgiprOMoEUZJECpRbhpN5CIlAlUGxibdABNO1t4UdVo
qw2x3SIzfb23XEv5TQEZYjyTVXQTzI6yI+FNrJXnCJNNGlG50sP9xPkRzONS
SDXN9ostDDTwoDMOvXYW54SN5D0wXuU2/ob6C/OxFtWo5Yos5XHg/WQMr1Wz
/frzmJUE4vlMxuJWm8R2XMUZKy/pumNV2oLOImtGY4a/lgWVRgHMtX+uH6fd
t4aUtYd23OgB01u2iTEsVBwuRHmp3KBTH/WJF0z4mpuuiSTd0+mTSzT2Mwh8
I+XSHHGAvI/memAC0BQgNBB5lYB+D0tTzxNLQsMvif6VrmkFZqmOhCU4bkaG
OafJWCdLb7Mnrac52pzWULPDqMt4RzaZJr028z2wLLmF52MID8VjA1GOsD4/
MW6aECsoW4kWCd+SIHJQzwu8x3f6EZEvNA8nPBWiW/gkjOzP/K0avpaKAVW+
WqQLhvXr+YbpWs+l3n0egSjFZIrqyt3hXlHN2ueD2M1HpeL7Xl7p3lgaY07S
iFvzV+za5doN6nXHnkuzvced4lwTxYNQFGQ3XmcwCvtvvevptso4WPZ1fLL5
Maenh4QFir6mGKIT7o27f1XcCxDyCaKgxi13BOOO+XB2MVFZuk2QoZTRf+TM
kt9/qTKvAF6/lN5g6uqDiOfUUgVmz3FC2N6MBFuSFTIEbeYePR43PMEA8JI5
/XxUKHd6mRrx2GTGfeYbsv+aiC/fd5vmxkk2BaLHDc/4VrSFtcLJ/Q4k0z50
04xPaiW9hq3F9zBza76f65CJ/yLWGMAIofEsx4wHgS22R4A7M2nEy3kiqhaG
CjlerNJbJ9xVBv668/iBattCV0XVyijbKgIh5pWPX3gkqwK6VBQLbNeWqj8M
h64DkhA+knD0gWNKEuZgTHnp8jNWz5um8eYMF/UZLAu+3Q/S3wNhNfQpQUWN
AuCKIQ+H5D+tTda91OqOAGbv0Svpxc8l0Rum3Sy+j9AH3YjK7G3K9coCVtCY
ugE7aCelKQxKce+VnO+tl6Ppd1e0i6BURL3oOY1gFkdkz6MsHBDfd7uWBD31
uTR/lexCNM1aQQb6MTVEoj0NZo4jNG8WD8SnVfWXqHcfcRwvlFZBCqtoB7rd
w65ryebRNz2r2CJ4FVFh40s84K4UsC6dq9hKiKJBiDAeJocepIq/sjv7BaM2
qZR+mSaerXp0ky8O8WEpHaRBM9OyfAGNmi0BW8AQoaz5Z92u/xG08feK/uLk
WI7GQEajUKHgCaDTWJqVnrRZr4JzqWi5wJnTCd7KgpkpnHe2NlhUzV9HzyAj
j4xoIv/o4ACZtrh/8HFxvIV08XDp7ZkR68D7ry6LJ5ThQH+OVgiUChDkEn2C
IIJRvjHYaWbeYcZ6aZfixThhJJIg+YAp6yHhvKW9mMiSF3/PU+0lG3tr7aSE
/A5LJzUC1imP5h4KnLsSniNL8/br6W35ND3I+L6e0akidpFnvVVScbZS7sQ6
nWRc/IVNUlFJAyElQDC5f85D3icE0wzWIZ7AgboDY8G0XYZvrPl0SLCO70AR
EcJkFizJFdAgb1/vmR7vT2dYj35/iTDUV6sAtkIYxjDKuH5xduqbUtA/kYeW
JdZiaUZH5eMMxRzzLlZx+guGyegs8l2EY69/R3vfIpsFiSmjjrrwqIJOD64E
l2QMGwAv+jzWwfR0yWbtJZhmDQun5ofJRHM/wUjcC35Mw6KL+AsT3jDSd+J/
z6wHi/WkNgn2lpmJxlEZL6rSHYOhDWTwYEjqDqWMgDJlQXqgt7f9xvPnclbi
d2TEBjNDOKGkzDeKOKMEz/zXMgcWEAzylVOTOnd6gNBzzuuPEVABq54VZl/j
jli9tUZBLS0+INbwkYtdkx0v+aAA6N5PUXcL9QaUGh35tl/Wh/cAl02lRsEQ
MazRHObHld6fhCUi+a40KcbkKMe5g6n/M8ho7LT7NzfTqwp4ecn76TY7ndB4
yii5BhA5pAIqbMd41TdZxMx/UQmQbhBks9PDnxhxv+p3Z/YVr4HiAo7J/sR6
W+k64MzxdpCxSa2M8SNs2zZD7SrnmGw/NZXHAwa7LjLthynp7nQEeztcLwOh
i/CMfPA6tHLlqGhtQkbV0wYY/Igrk/MgjCKydQTjWfol8aijfZhrwZsLyMYE
vblQRiB2frLBNVM95h/1vpXZkGKCxijOpvQXHWfq7tmeqAetmcYxQLwMS59Y
JTs8JXMp57xoSeLyHnMOOAtqK/xSGwpgm0kX3wG69A0zOQw5xIPYVImzX3Yj
Y2BLx/zJkjLGyw4UyOS7gnq4UVcQRzlNhzxm4oaHe4XH/Hu3E71p/4rMXKDM
6ODfzqQDOmrW/H9YjqmHLExChMN2GB0p4xH0K6QB8EgFKKyJd+FiuL2Dz9yr
Viuu/a13frwhviy95QvEFNZn1wjDhfzQ92MtrmZln3IGh4uAnCNQdDYw4nMD
RdIq716NNuokUY5nWHoj60YLCSf/QFQvyIOLsdWGM7do6WjSmdzM4D3PtMhj
nqsuGJfqzMtMtpK084hxqGnPwSGq+Ql3StOLz0rFjmAbOKP8eH0oUjXbqdBC
Rr63IaeUGebcRoV0/Nhaic1ndnPgD6VtYz71Dk5KdbJ4RSmzjpJUp7z8b+j2
Wb95i7GbIHO6iEfHqX+YnWmp4IpdonkCMO9AvdAa8j3FV98jBBzG4qBezNI7
4otTdkBM3CxhHMna4ew2ye+saRiiL2kq3AGMdrl3Gjb0qM6E04K3rq0HyV27
st+bOwPYejL33D8wMZXu8gndGmyiwgih0SERICQhNWT2nAEFi8gStTDtByWD
1wrROFIJOfmH3QtibHMpAiOrjCS5y2ptZJVpeJWc1b9MmUuTwQKkL1mdRPjA
X7mcZsJhqm/E0i8lJWwIKdhiQrn0Mp+mSGqi0D/oMidlxe8N+ZxmmpIwtqTY
qu9083q2evFidb2UeDfEofUERJ5LBkYjFXqqmHEITusCFyGsxGLm3SyT0Ji4
TkTxYkWm5dTggGntx4qs5nXVc1bUmee3tILiWa4RQfnaRaaISZzYL/mC9Ix5
YuhtBk7QMwVXOS0S9QBJjBvdNlhKLo+WJ2sRENN8lttY25TrzxljXWwTKViy
QsLZ96TbwHheY8EQFhdDKMi8W2wI769DFESpQ0koPBXMCWvpUCGKh0JKt9/p
rE3WWh6MjThaU5+UFZWOev6Yf334WpefrzT/O4tqZx7JK3+LxAks3N0/Ln2q
Ng+NM8FNqsrLl6A4DaaKYUzz7Mk9btbTYF+8Eiauu5VSlMSTdvE2rsoadLUv
Q+pV6+P7kAC6wdt1De0kjEeJ6UV4+ksi1XMGBwGGNnArfSb0J1r4L7oIB5MT
wLA3/S4hBmdUc39rsElr2sVC3NTUcqiHemxpnFTQiw+9iw2qIB2tiueEL7JZ
rPb/OHj6VRAenjxEvkvPJaOGuxr6ZB82iOffdvovmf/V82dtKAoSg4UwfueY
ics9I2KdkFU/cbhDPFU3eQrEx0ml9BqqjCXQ2i1bqjCadz3fVSjw87kV2A68
p12QFzBSnVNez3XQM7UuE44gbP6APpPICsOqqvSUV/lHObOf+MVB1hJgN6cx
ymC+tY9YdDkCJ4e9DlJAiALK2C+pYM3jmaqGDUcQGNYU9kmmheVFb8bwM24C
BZyNs9nT4GPTOJZ92WkKyi9pHKTj91qkvo9EP6aprx6n5A5WjMuPmQ4SkgnH
Mz+re9TnU++Xhj5cfEQSWty9BUnCpmSs8VW1yjQEplXzmWEqqUaB7nkAOSN1
m8ABSbaIkjLIzQ/3nKlT97j4KoQLtJtT52HVoUPpypbr3XHV/0tsnHaJ1kdV
NvtLXm/3sRJxa88/QtmGsqKlTshIG7O/pppJ4SVhYG8W+erNV6ehJeyOzMgK
QpDTYOLNeF/VdWPjew3kishNLBRvaILkXn945YpxzrPD2o0dwCBG0EVDJxqn
0CLf5hWCNy3tfBzA226yppcysOk0dxosyFBrux0f8UZMb9f/X8Wr7so6DeGb
86+6BX3079xX2KCK4TTi/3L4Oz/+KjkUj8P498CMpKknaDH8KfcpZ3+25+L3
YKSE4h7+CXnOjqBGW55auOFEaRRqzWLIU0gGbMBFbpMLMqiNeHQfY6taEQ14
+05yL62mH0f+qvY0oVg4jiFOyOtjvKUHj+CejTqdIccA653OD2LEUC3K+OMS
wVL+7ua9xTLbnw4vEi47p0ViXvyO21+zSJ27DDBF5RsmOe02UuS+0zNmgPe7
wLLoGRt6YQ3JLxbj85NxR/bVkOTraxRbwy/JEFxaqnN42vkrnHw64g9e/UCv
y3J0MD0OSIlSHht2WBwfQ3ho58u4BjAuVRTEyaLFEjhmol8sBkPLbTrD5Z8k
aCe08qNU0LcpRF4Lui6VyBAC6cdVZT0ApiG58+Uz/bSZJ7scYwea/BaIrRHQ
MbdMVKqcUqgFZRcU8OeZn3STyGsFu7IBzVsfF5qx5vicYpuVevhJ6rdA/l20
sQfaqvMb9WfqlmU+AWlK4d/ZoNNbm4YWNHRvsDdsVHQemLQwDC/gH/Aw15R6
qkumo1qzkyW/S8GWZKpwDwps/A/wuLDMKUDciUAUoIjHagyzVLkmYq8BZ8FK
kyNDEsKWCD+BzutK1Hrd1Gl/NNkAYEvKMoO5sJdo17Xtuk526esCvBpKnF/1
6fGg12EbCPV2keENAuvsSoQ4GiqTqKGE4VzlNFQaENnl2/f1F5E+dYW7Ibu8
BWAiF9l6ZOqO26JjyS6PiTuZQnkINfeJKM7NxylarpZctesJI7An5lJh55Zy
b4CDpb11fBovBFwyMbXKNQD3r0peNMVT4hbGQgiVCCeE5mvdWWHWvovdGMPc
ifKR2OR/3Ws2gmkwygYMv86xeXaGj6jXmEOlZJloXo74cLf42qRDvRMbkYic
Vke7EjrWiu8OiNY2Jm9/P+WJCI4rYODxo+qxOEP0Ubkk1LwTmtoW3LNSq8gF
+YMsheE4zMEMWHQdoxauLHMpc9I5GeqxGUPNndHksWV5p0H9Bm8oGoqZmL+M
3o6jQCubMjgnXcykt4u7sBJJRyGQ6mpANavdXoR4PlEts3Xea/4q75H4Wf/X
hYwSaZrkfkjP96nFkDQRXwgwTIfWB06WmgLX3jQucodVoAJ1FUfOl9QUUO5C
fxwr1rIJ3x+HGB3aigIqo1OBliHfOaSdt1MEPHicOaxtpeF0kR1N4LnYq1zU
iUeDE0YFa7gl/5zqADyPNSSMEsBadajS3KD9fNJuoAV1KpUXJexmOy4I6L9v
wPuipl7KB3vHqUzPIhGDaDVjN5rTYlQ6hhA3ik7OygKi9Ph1hwrPh2jrCort
UAcuQ7fz9ZheqnIN5qeRn0j82PVMkBmpEqSagjjzjLEumnBiymI9EDSXra4B
puGHBL+/Ek65b8PRIpWMmldYeBtGWDtABEGndfbqyywAGDBdqHgN8K0iBMcm
7djHo6Y5vLeguB5RiFZXktLfYs02BMs1EnSDva4IRt7rzcztE/NtR7Ea8UQP
6iol9E9sC3Hd9rk9O4svlj67Ids6fwc/h3SNfombxPzEsNmk+yxVwVxTDeQ9
IUcxBsQcM0BeXr5nDFbgdwexECBLEOv6GP7QZq8aR7KJEbFOd88oSDqUKcHi
GNbinS1JAc5c8EUWezOWdK+2kvC7K88X8UXkuC/72KV6sZ8uB47YcSCVVBhO
59Cfj2bj8av4cWMExmxcTQpn23K/LJwetsuSVqgXkZUX/DAua/4Sk5GmWAiD
+qISXGod9ZN2PDSU84ojXkKQo1YCLs5suCjB3fRPG9gc94BO+sULA1VdDU62
DoIcQGtRwhxV5QDPONPtemJe/nkVy/kc4eWab0LTV3qa/l2emLMvPsEMDDQv
NWIMgsYl5S04+gytwVliHEl9TQ7tDPjbixK3syVAQcy6CMzngzuCd6EUuxhm
xY4LWtFudbdcMuwDRLlUh1S4HbjqI8smTbqHmrllFggLryrvtxiLMDCqxImG
P/wZU8bUcStZ16PUbeXYMhPtiCmbQLZNfXsmPBx5+g45GLSnkk3LVXV0ssHU
wsRbD+bUjByylZgJQhyEb5X5AGm0JPdXYTOr5Ccjd136sHT9Jj8ugslhnP6G
U1dkWgpSKZpvNMOu/l58Z1aLUfcTF+VMHMMRXbmZFneVrfosSKyeeqM4rWMo
Bd6bYOHIWvykGMClJjcK5+nRnZS4Fyx+gq8QbCM7XMih1n/RCDW+t471Pnbv
mFKlUmfD1HFFhClYTN+D45e0Di8fYVePNevV8k7dtXLSVEQEL4p4eP6LJBZ/
RJ/ampXz3m8ZrHBb335fTJhGESOJ5chnr9Zy5JwJnSjuixtJTCGTW0pEfX/R
3U5laRa6NOcNUMz7ze1b9vKv6pCf/yFL+RaM6AITsTPJKslfOC5BScf4WQvR
pP72P995Pah4mFrgv2mFnyGHWxmGReWzXHYllXBwqmt5YEyBjHmToQLtXKru
TMPXPteA5pDubcmU/dwiFPpPmxI/+KNkShVVdNh0/+dgE4YEM8CNp9U8guTe
cf0DfXN7yFpo9YE1e57kbsvLvIyfu88clKQSYd5Mq6os8Z8ezNaDF5Mg5BAT
0drcqWysdY/ZQq+Q3usrWSTXFXmR4B9BSyYjtaR4Q8Rsw+LZCXP8beuS4YHq
NtNSNa4vIXjS05hpsJ4vqVCcG4IVJYx58D9nl8E6pku2ct1nRpP1G0UqHiB2
iYHNQXZXrmdLAWNAFisVBkujIk9yVT8oL9Kmw+vXchnGlwCBmI/XZ//7JBkq
KDbW7Jbw70rfuEtgq8Bl5t/RWmM18hvFrtDf6bGZG80JD/F4VT4z36KLDaL/
PC8gm4reNl3K5ILx8lflifaOaXlXaaL7caZkNE7UyG4HGzF3YHBM6n56tDN7
hsVrvKTBJdg16p42anNLOSohmih4SGBwdSdPa/PQwH2JSFqPL+SZduhu2Q4z
yerD/Lu48hX4pKp5BZYqis2UKFMBUWdYEgzEdZ2VVK0Eyd9zRl1v3dr7N4eR
GuAfZMDf4s8tpbo3qVfdrfCpQ9sLUkZxLHMdig0TR+9ab6PqNA6jDk/nCQrs
0s4ByY/fqTrCu6IRsE4vZZThhDNNKnPzHJpbHVPiJaH4v7sf9jkYUG6uXobQ
Z1Fo9elmODBz6uCS565AlSFR+gSHf2hBsRGEqp1k+bq+OLpcXcHKFCdxugFp
rdSiRweoihVtLBmgnxgR0+4RC3RKu7UVU8yYQz5OkFXAfzEXWqCM3tATKwUI
3XzBwqZWBwlL0oRRfbzMxSfJ1pN7uk/LaSWwwclXHjKl4LHoDwGsD7n/2nF2
UHxeReE6QFrYJxiyJbl2qfqLoFRGBLvNbhXcG+M9GY2CnCSQ7c+/EQhlZi7C
qJVdJ6HE1xgE+fMuyvHKYbg2uMN2nukspo7e8MOw0u0GU2Qh0Ys22Rqn8U2V
PobAUMyq0oPsAWXZN5LZB+62nsauLroN8BZgTzKl8eQfrCP8ZyL3gHclZaRd
JjEZeEU5rOIp4i2ibRvzMxfMPCr8c/vqLQet58og5CohMgrp+dvfUk3h27J1
yy0evauSIfmFAaOBnY+idfUc9gv8PMGLDFQrFEkxJrWiVGDBnkXlNh6lhTwR
KH9x3CLFr/TnQ0HwXrYBV4ixI+dHO0I2FFom2iBx37sBOlma4aPJYi8/Pmsi
AUdr7CmGYPtB0viwnoZBxycGWRQm+xJ+k1e+RhWKu+okjNI0qQ8nbxLROaIz
Jufn7ePWmCmYCG5atAqFBvQkcYbEbAjEPangAnhQlTM/4d0OadSzoT6ASIW3
ljO7apikv/Jy5llD8BRMrJcwlVGZ0sMef5weayg0RKjQRhnLUxxNZrl75VsF
7x009aIQsgOeClPCpRrwzjsTvCl3MIV6hbjzERH2S8PDrjTIZuAJZvX3cFEh
AdRowbfRd9Saog2B8/lL3vbJMgeo6xornD0ZqKfbiS2l2xW2+/eafvQJ3MIq
jk/Tk1pe9GMXOuElUbQILKKf73AQNIJSKTPG6yTjuvH2qR2cGd94a7dhaNhX
Mk7qioxq93mQ3GgHbNqyd4P31HQNLWUq1PagDVZ+JgVPVNwgMoiSFpSQJC/a
SH66hBDFgPgZBF9Zas3olIgJpiYLeL63efA6vTqH2d6ceaor4sBVHS7z16ic
DPr8giUxz404iDYrSOyC0g3XiIWMYT1+0UhLSJS5oufIE4ioq2Hmo4kkmimW
qKyFkEQEAtXSngEtXKfYxZqBnjZlEql/yAvkN3hIkLCPiCfKDgeOaGvD9RSa
vxiHkenWlK7PRQKGHbh7ILYXGfGcldVlrsB5+QZlB/223X6AEVk4E5LLtkAJ
Gk2hgaAhXBgjByNgnGHKnLpeLXxVGEdSX8ADa+IKr7uxXb/19cplI8Wt+IZr
tc2id7QnlZ+2MkdYrzk3zs2AVN/NbCWWb+is5gfOpQ7qr+glQghiMzbYkGvq
OqRmMqor5Znf0TYkNUEJmNzKod2F1wbbh/isXsNSkl8tWZHK0OrJaRjFE2Sz
DN1IcFFpsW3Mm6y1yqaHBMWQzof+tmM7XAoCmosv8gZ9mVGhOpsSrbG+6gQs
SebBOzwpnhsddO0uvyBSLwriwjotK7p30iNdUDbMMAA4dSrljaPEMhfwQ9FM
DTU8DZIKhTr5jxNYNNhj54oJZm3+IO82BekgGwfqdhPmGU0Wr0k83agx8bRc
vXYI96JyL75vS1MWLmN+ZXC/qi2rZSDGiXLIkWXbhHvmTheR5N+U7lYjuKuR
QGzK7cB4+zqh18cqP2MuD+ZC+12Fj17AxVMwoyOcY8Kkh9qEwFk2W0up6kAD
zUyRXVm6IYpLUwOmECCNhFCKL7ZpuPhFAzKnzptGpiayl9PqA06OPqlC5g5S
PVwmB1fkovLDcMrGOcCwQLt+/59KHkwBy9dqQQlV4/0os1EKYA3WOjlJRR9A
rE2JVj0XtI8jxPq/coQm4jT0VKd/m5ORchfwsxjqKMm/WolpjtIDwsJwcAMG
EqqfBQ9FPQSeq2BSqLkmDZehfBOUEMNfO/7ogC70bVo0d0SWILPSLI2dC/zf
03Ta3JWFdwngSz2VbtnlyPvKswJC3tOlSd+lfQIsV83/NF/iPJdheQciE1Yk
c6qwe0Pm9qVpu1FvEag5d20UESAfsrE/Gmfcta6e3kcbOaqbW+qWkUEBgwgi
n4OVYMq1eqdYDVDRO0t98Jiiql6nXlndKW/Wy+SVcKlPcdTOsbIiKQk06LC4
nRefPvxyh5t6kth/KL3jpEjQ0N1XqjDtZnN6s8nvz0aDYau9Jv+cr4dpnRo3
0JO8K2iD/Ykv75X3RqxDjomCfyRkfUNEsxKNtTCXQsc21ToFx9G3Hy+muv4Q
mouenFdTfznWoTfuKc78Xunt4g4sbEzSkkKCF0r1y0fNoaklRewcSFasoWr5
9XX6HAxYtpWadnV607jl/7hk7k6j8SCWEVUNwkFL98obGiVSppDy7oa2XN1h
eyqMs3PVMNcqAsD6oC1K02pcdWTxVvx4oNiqLckCmNcIeYmvJQ5JwLd7znUA
JpaXGhTxHD4IrbMsIoDvzq94qwnjNFjUwIpyiNMjetoyAheic61cT15ol72E
GZGRVn7qiCQ8v73BF86gOIVvnrBpEX9xmok3Y4CvIFQgygHMvFme1NluRBaR
hbP5cZ3jyJylRzDYZciXhlJJnbQGy84TRjZO/+aSFOmdAxdaU1JvnYDGTvFE
lhPyuM7rWsT9sxKQMCw7UFAVxAkaqoeZk4N5JOvvCXjobyXGAn8+Vo39K4Q4
vorSKtPqlCL1iwBdyv28Tw6Zl8MXm577Vkgk9zo8D9deXrtDOGydgRTWc997
klxryZwwzQU7d7GaYXFqjAr9kj9AAiDeXmjdvKSwbtAbC55rsCWGgoTiflE4
Lki5E2xkKIKadhpXRuMQplGAaPTjmLSFtDUtn2NW7LJIL6C7VViehZfWEEhj
7GWtpgPNmW+joXdfbK3axvotM6dOGrOQtQ1wgit2tUlPeQ6y6m59Je5cazdo
0ZTECxcj3Kuy7RffbTz+y7fwhVFQsC05rzEKxjGQnlGKVXLJMd016nBMnd3Q
TAbkt5AONjd/P+zliiuWRRXrnDdMk0dzFhqJL6ejM4qHrP+Sf6StSxvZA00U
n9pOlP4dT1mDKfBPLb0ARwptszjcxUZHXrus0yFxPKRNP/C6mXkWCkAJwjlS
78EGHB3cXaPpSzPle8KMOhXAHx0ciBl0Yz1EsbfOX9icP/ZQksdUvJYtJhF8
INOdrDg2a49oC4bysOpvliZ6tyMMmLDUbDmejAs///DbUKbDneOKLqG7tHR5
aOofJhQGbKHnZuDl7/QQEPChjs4KV0CkKrQbYXTpZ4spUy0EcB0KR11jKdUg
MAqQAv99DPBk6URiYHnQSmJo+3/ehbAqHRSZBo3S5kc6rLUBzmqClDWHy/4F
onqY7Y305Am9Ki1nN8Eb07kMUriWG8TFUeNINeC0S1mFuauBz/gi4/huvDKP
yolAsHmjZE74PUFq9R4NvsUZYzioXgVKsn/AEtiCRrd9jkV9sBkPQB4s6w/z
jy0MDzl44PZ0zthJy8zmsCI8YoaKyd0x6nPbg/UlGbc3qdAlUQgAJgOXudmC
Ml7TcgLQ2cpAg8qAun2Td7SkYGX/5ETPOKiul05Q3x43PjVxsv91T7liHFnP
TtuzeavdAkUjD0lXCxLssty+SgulshI/yrJXjcoS0bPCcuxqJ+x+O3fINpCF
taaNFVpdvcF4btrS8KmGIQVkRw6X3xy5BfP8+g2pG61oHbKZZARMMyMWdAGh
Wp/yvU42ZzLy8n2a4nuQRXOEJjydyxZEljF+HqVDNS/6Xc6Vs28nZhK1bttU
u+GiGqV3KyROsKXzVyniZn1LGIEUhbPjcZNpAEvlxuHR8rzkdTSL73EQHInl
txQ1r+fie0w3l2RgmwBF4u1yrLL/2nV2EAjRH1Sq1mudgdY3ITYPZMTWDHzE
Wms2UuzFWLGSzVeP6IW2Rje2+K8WlTNfIUTreuKjANBRrJ3h2XdyLs7Wpi7D
QOWXCZ9OJnmA5Wu61fMFJwPftVj0W3nYJsZu000GjqNoHqEnh4zeBTz3VCZe
ozDRtJZCgjvG3KrmrN4Iel91I/I4Z02y1PQMFltZ1kYrknyTevsfWDQLnzJj
b7yd6RgeCtl8JFENiQv+Y40MV4rqphd3b9IvZ8uiF6K14sH/g2dvJFnrFcNh
dJrNMHoA8Xfo3mB2wZwyOsvuaMZmhmV6DNfEpunB0t8X0sGAoRGFOhtNxK+G
cioFVT6PtMDUI/aMQ7KcmaLGf7bXp0/61rJNP3reR/TneC96i+k42mq3HngR
gK/WI7eVoeOQyk0wmGob79RUYAw865Oww2abR0MVw5v78m57F1Z7sF2+otks
2lTiQnpgH6MUitlAWCa0DEIJX0QzHbZze0jIn0L2Vww6CGZ9i4n5fXkDek2r
SntSloOsy0XXvYXsf+G3Kp1NOOWsfT5eG7gQvMLVMteaEeI1xB8aruCDLc/n
GmSZs79x6BUnP7YULkKXtYzZPhLiLPyzYuvHUffRIuuffl2OcT8iPi6aXprE
ZH+bmNAMjhL8Nq9YdSNIQbBiw7lW7Yg+r7ep8WcXcx8Ycogi0r3FrUb26IRd
eo5iF4fZZT1vySMF/5lsmvPxocR3qmD0YoqlI510RjW/KxuOAgirH+9ZXNRi
/WDNKWtYw3YXzKvg8Y14D33Q/Ni00lLbxUpsFigqonjrtRDd94yr/MbSn2vI
lE4r0uNza6GI4l/xGHezeJaSzBb2iRpJg+yTOr4njeCUDACxtxAV1XtafI0g
1bCogrfCTLGxwD7OA2/r3TYHjpH0apFXTgwGY1LlpQEGezV4uEMxznvTvXRG
5/YQ7wA53z/jtfEVhS7/fQINsX4jjAqFodAYC/STRDrAua1KQ17JF+eCcEDj
h/hbLRzJ0Lc+M4XAS7OvPn/HKpkmj1vlk4/ApU/+yiEQuVgdGeVY3xdP79d3
pxtjzqDAk0sujzdlJN5nSV/lYdOvhFgGA3RTv+uUK0V8mfyASDNW4LaVmvle
Mii7M8JxVV0mWebUwtKR/nOgms0ktVn7LihLGda3GBeAMoFYUPBY4OZsfnQB
2T9lgNI/zEgiDXK1vLgQbbLf/cQpALVkS7PQJFIx6FvaSZrhkdstYdybKm5s
BCZYbDoj0SOGmsU6kbJwn6ity5KqKggQbFPaSe819hlpbnkGa3fXAHEjDnH6
jNTD0SFKZLepRKZ2fxpBSVAH21WVlgwQbdj9b517qCLSVpo1q1ugNxAdWlVZ
jW3rR68uUArkNHHq3Zh0npYtHJE+EnxKWOjxyZ4LaIkX18IUyVZM6N/DBWRc
JlIPckeNoBYfeuIlaMvXxBcZSKkfCeysgQojiVyLj3sI6kNrLg1e7Gkw05SO
/gArOZ66SXC5IQA5M7jwCbJBkQv2ITkOXQqFoapRkBsTz+xkT7OAKoSzVEsG
4npHpNoupwvX5dL6Lu2GkpmrK0CqVxEBBAGe2ORXt/eT3lcK2yv62xT0yzER
70GWVi30eo9uOHsUd4hvp02SAh+lPIv1TiZF7h7nuVHT21xvBouQfmNLImpb
i2zlgY0z3+XJHO3qiDSx32r5PZKGSs96tMzzLvwkNSKt6ccjS3VmcWBnktKy
yk2BGfbeiZ6pglzopqj6gQ3GbwIi8fTeZ2bxJAJkelb8YNWHjGQOz1auY9VW
acUr/rgefQrYdKIlrAwnRZpfxLfbei3GInQ0tAg2gBaYqDYUAX4JvIxScG/F
xolI05ryJIBjlmSpqixzAvbAEOpoCBl971mdjrTcov2N1UAoPusfQ50o/gyN
si9fwJ+9pjqJ4GoEdLhOZUZgnNu4wCKVAOwNwhrI4EPN1AtWb5llV/NbPBCc
CPhSoteC/jgXAFtYl/554+Aym0NFqzOG47f2UE4x7DW5DwNaHHPE1MmWCXEa
fOoJgucZsE0AlQ/zK0belf6LWsq7cQk2tMNFCEn0Jlxhrbpg6fCybVzdyS0W
4d5dPvrIPx2iqVoMVLqe48NJpadKrXsqj5q/zFQr+UxsPm7WbjbksTqox0TN
EaYQ08Dyw335z+BhqrfcYw5t3ewPfE26zlbKDeDhidRzz3x+Ri3B6Xp3+nbs
i/GCLTdBSp2oDpHGXvKHMxLsdirlfr0IIFFjwD1P434u2y2zKmM0LUbkjKB/
xErqA3bB+ONwCiDI9XZBQN2orRpfCJ9pTHJFqr/UOEbpVqkR3E7692S0SSO6
E3XTGBXtEuhMoJtWaaN419C+MZNHJq10B0qcuzE6kveOhfku/3jfnLVrEjhc
EaPhN3Me1h2cPSjlt+IvoNgmpLylOIq+hGy28Ou+HGjIrpxXm1LoC2D081Y5
CQarD62gEF2EIJIbAmogkwmaMClNPoePm5+dn/voNoxdos1fO3DLvVfJvNGN
zvhYbuh1anxNt3awJgZbs7r9t0vNtCgfDU3lkw7WHtJq7xi0tPc2VTYhTBTW
IoFZ73auRM7Srxh9BVOXXYXluEczdObxNFy9jrcyKYWE59civf0gXWQvnTvZ
XJQJX0hoLqT79lX2VWUViWurgyN2tbFvaJxYUkx+uK0upiBcynNikLi8E++c
BuOmejhbAxGqLndD3u3zKO9Xi0h2xxYAO5v1BMS+SNX9rRLJp35rFl/wUtzv
fIqBurmFLFa2V5A/OzfWAPU3EH5vZ06YlF0Lu83B2Qhjzx33LT7Flgg3KAuM
p/1Cbmzl1bOdY9nmSnVES8YM3UB/viqVeY2VVi1Sozd2KQAwEiaOJNmnM6w3
867CTx4h/wD0Uq/cZgyFn50M6tfPdes+J5/EnAeEbPmAYuZCm+rcobLVDs35
SvHLa7RGg3f1NxoNvGBW7tcPVMl69Iif74/DeYFo5+LEDaQnQvE+//NeJOBq
QF1v40yX3jAwdsInKMWTiJ7ZE8wdeIKQVWWNJnl7Z6wWpi1HDibLlfwKMt/E
XKXB80DtOQ4R0XueTEtsRm3s77kEWOWPBWh/ZMvptIjDuU7X3qO3oJFPlFo/
ukXcijm0YxqCiZw1mB0Wkvp3BGEpTVf3UzYeAxMYb77gTIXDvqivE4wtVM3n
CYDJBkvlhsQ37Rz+Ekn6JkYWywJlGBYSLBplhdxCj0S1D+k/IYkP9Dp7HKKb
gt3FNbJBUApPOEdH3KvpJdlfihdlZzmXWqXrrikRkyINml8WN91bUT3ydRuu
GDkvq0omtexY4s97NsdBWP7CrHtPZ4rFiDCPmwVJIfriIqirL1D6s2k+ZZgJ
LCcchhMfIIHGT3s7C7yuC0ZMwALq4spclvyyM6X6LHCL+ik+45ps9EJwdsi1
8sHr9sR563JR1MbUxvyUpMeLOHJGfLp4l4++z0xtVn1OPmU+ZD9TAl9pg+To
MmpNoAc2GFmHFg9iSZGaE852DOqoIMXMiFSBc7Rho93ZpeWFxhY91WqSJXK6
dNja0AbP9VckFiJzIFVK07LsOUCehlU3iY6Z/xV0zJZi6NEwBIzFZ9WPCEAc
slsQBxEX53OHRUd0gYcjgFggIyGna1EeDs5o9leUcwhs/uafHmFYywf/Mo93
usVMAizPQ3B/fOEq5MvVI8wLBVVDzZanRvzTotXtNa1jS6uuS6nRgzt8Zix7
F4MIS+1GV1PC4ZD7Z2TWC3gLY87hI26WgK+XV+xqwXECPUQ9k+Qzmad8iWIu
9GDzKJNg19BzZYR5W1AtoxaTaDddic1inMiG4s/28kIrBLuYmUwORLwXZJhr
8PEMQdgZ8qMSC/ESvbz7tErweJ2/yQWmA11RbIw5WOLxJOFaB7je89/Q8KSa
O/qXA8N9LJaipaRnJwc+IEokwxbjJi7DD4Zb5boBdpeKDlEaNuPvbWfOX2+3
/OjZNdYrkBZGwp2gDtuP1l/DUlkP6HkP9T4CE/cQkqj8idqE7jd26nHMBSKT
OW6VAflQSjxTdIgDqJRqkxrDuuyD1EfmFedpbOlte9XkZSIJ7+LDjwIFj8hH
1V6fw/XYlfyT6WuUh4O0TyjOmKJ4kj6DnHZQ+cQnaf+qL0GsNDligVsMjG9o
u0OPw0ALVuD8NG9I4s1bLqYwtdZ9Fz/W/OK8NmpuZNeo83lDjznMgE6R+Mor
E1OlMQklCZXlU3PIjnpn3Bnri1eHgwqx4+1QvIhsCA3InK+EWKq7a4kyOiia
64ggazsfXUbB8JgaiGcFpBHRJ+4EAJwmWpoEewv5xyCP3ECekcFyl513Ub+Q
QNcDuMfmWtBhOO80GWOD+sqzouij99iIL38/2Av01v7veW2VkwUy/C51xIT8
A45l5rCVpIjQceu/h3ZMmTiwPMLov6rkrC0rsF9PVwQRtGnOJUGzocajlJuD
1BBPRTxRdaAMhAB0Mi/exfAZEIEKBZHF4Rl6SFzH9VRnRsmo1jytcZEmAvcF
0di+hh22tKu2EM8qD1EpotaH0q0gzkXfXvaZFp610RPTJAvs75LL83jLVhIQ
XJ7bYied4ns6Kz0G7u+/5nNAvmvurz7KtbD1JOo489qzNSbD2pCeY93wk+ld
adXbNH/Bt0eDWu+88RU64rJCxVj0U6CT7WoEW6bdtXv5LgbG2uoLtUd5v1Qy
F4xbw7GFZKMpS8HQoD8vfwrqNIjOt8FVfwtLe5iLue3XA4P/G1VVO4lcVC+M
Ll5QCvrkagG12h4Gt4SKa/YT0x0ePGWtqYRiRnfw8WIhWX5heIowuWFwr6Vi
abmYdRedKTiNknssX2qBCsHqBHVVRVV5eOZJ5c7koE5s1MJTQ8y6pI8YPgXG
r2wpvR3xxqlDP/nD3UupZ/TWSjGborw+1cBFHiZw6mHeZx1WLPo0yXRs6xnA
c+5bZab44LGNip0rmBzxbKU2KUZszDntHx49/NEZXaUv8dlHHvZtqfkgmjrZ
LcrA558YtCTkiM7xO1e6YFc0bmevG0ukFbshxNTh82X9k5dC/v+A4bBvIMIi
/373NIW4JpQ0Va3GyH4y1k+MAFKPid4qp1g9tRpHqSTSuYnUmwxfLF6iLNt6
oepwioRgkFFwsTPnqr2aQvSv/vo13qrJtJ1U6GZEuwUxiLOjlXWKD8P5hhLf
r245JMXlhow/1VBehJzVrICW+9qiN9FoHxtt+kYPgYiWMAD3g12RTEEEevKe
iUzoBuHCm76mcfAnArPI8Zy3zdFOyy/MnPgGcMujRvCafSyyaZmGJg3pwq1N
an35q8kPNFid/RW/Q8aCXvFSiqKTWS336gho5NI8t9OFSsX50M2X9AXaGWEI
nTn6wapsZv8vi/c7FIiDGN3FLr6OAXNQF8ZefsSPEXtCjK+BK8S3eUxKL8Gs
jn/Z7ZvwqGVUSnCEj6Y2aGRmW4caaqVb8pbUd/2G2T8ninkLjsNtHu30BKPn
2s5/IwoApsvNdfS0hahQJH4ZqiuTr0T+/ia9zfM+7FGgPz7LETDKBj3RyT9T
+tgwdJW8RzHMDa+ZGhV0FHrLARGix2rChyJqwHuWVfm1BfyjYAP62bc7lEEC
6+56pYN8aigMcduI9fsKNeuer1MLTogUErHICmg664xIJgmH8pG4y/872vvm
6uud7GOr4Oh8Clpp/XjAgSt3dd6U4kdPw0vnDyIHQ8Wf3yJKIN9orh+Ui3rM
znOkLTFaWRFI6bmbWo/eDEsfRVLieQKd91UmZOZ8O/EF6fSaXOmhaQXkA4nt
fm9Mgy8ARe23lk1BgYhbvDrqNVoAnukQatfHFD14UlHQNRVdj+8OlDZfyj28
xh5NDbXQLHg368uWH+7of1aHJZ14tkF3yLDzfiU5NosuCCZ2FLGmH9s6IZDU
U+3NoIyVZ3KespMr92hCH1qm6hXXCS9ysvgejzYZMzht3o7C8UpkFhRZ/Bhv
VC5yYukjz+BWayteSd7C9D2SfNfW7fyXYfC34d3+X8zX3UL3bAvsQIvxPWCn
pI3klDw7vp5dITWjLx19dE8K6btphXKk8su2UiYmCPdZWiBQaVD98PP09fCx
f2CBQByy9ImWk2+2XpEP381ElIhUDasZy37AwscZJh1D4pofU7hTa68apiNF
63VTCI+jvfR3lm0PXVcb4MVVDgBh/Usi9h+/igiITI7CzKq8l2Fgmi4LNvOU
Gy42nShtwvo60nvxO9HZZGWVNeaca2flEaj29skZk/Iz0aYdXBzE0asXyXlp
q4017DP/AyFdBm8v6+G/f1aRR1X3sexJbMAi85tcFIZ3k3wmyaG9Bz3NFu9t
gp/1sXBg1sZhJy3yHcNEe7+ieqvu9PAUmNr4M0hGFxV3sjIXE9uw/etBAMi0
te5UxZUt17F91lHFOH3AsOKCzYo5gOexQgTOiFp3Z915VrbLTvabncilkQOr
jMBkK9wCrtv6Q2LSneS31qkzi3JGHxvskiZQlqNxFgItu05E0ermF2X0fJzD
z4VYTZ6nYZ+osJE7B/Nh9zJXWRgd+KYA4AzfKry7I7oiL55Jl3248D5GbBpC
/Y50+bSIR5aZNRjdjU/OZB1csDEmwanEDXIO2xfOn/387PHkoM627pMz0CEB
m8ugYWZLt1g1be36morMvv3297PZ5KwQpl/+kAQnbM4CIocM4RlAdfSjlDy2
E8z9SC80HkY9NKlN9fk2qIeXk0cpYxy8WhJPjs4Iz/97Pf+02eaonMCnLgY/
xGLJbb9B4qaz0VezzOHEDTmU+KJU7wTPzpFok6mQNurlGeGZB4uh8AXD67Zo
2J9yunr/xkG+XZLrMJ47b6IkoRfBTxMzVZLTJydIMq1kyRUliCnp/Mj4l/RQ
d/tLz9lJoWS0y+B2XXeuXz6RwdAc6zzDXF4oydh8c+OPXauNvtcdLJxQyoPD
qW5Hnt5bfoCcTeF3D/hjTE9t38KFGitxK+kTGzu6bBun9XaM3fQxVXjLB4fw
h2L/La3qsNq+i9wLzEREYWg2l+JCCmU5Syi+kdFP+voWx5dyJUlyfhrqhtF5
QdpQlKjcvGYEBoVfR93jnROlxyN7ZA0V601l+fWDRCBSEsRN+KZlHmJYRqso
DnnnzYYjlSiXp6qNjpjWtB5P2DsUbS4tq6LYnq42s1oRnG7p4PLVWgAu9Zo4
ojDK4HEy5ImCUbHOkwQ1pYfnThcCntQSaK+iNK1SlGtwdZBdOMfQYDDueM2u
LXgj9tNTYIs7Fg1ZwdDkDAJ4g/gg/fl3pmI0jBqMeD6CZHlmr/uF3VFgaNuA
NvdcCniZDKCdBy5n2tg5RcN2X3MsAFz/0g51zgz/+oemVuq3GkJMf3wlXmDd
aHCw1dqRYRmpcmM+z+rh1IpSZsfG5HQwoqsBdDDniWrcFJX2Jog2IN09PegR
3P8eNUJWPxplMiQgMQfPDuxtQ90l1rCq3hi8gyxDLWWYizCXe2GVvZg4UNmW
kIUu6h1NsOXrSbJTtofjUimMyzcKTFxK8Jg98B1haqCc4SRpAbuzK4INt/bh
OsjVNb7yNagizRv/K3Zj0Iun1mdjRqDmy64tkZyQajJ+cDk+Mr+2scfPpLJx
vGQg5HV9b41pHN3TYRzBS+udIIW2xHXsR5+Zld1QRjqWw7uDniRgKUoj0ZrG
F/I6MQArx9LW7dYSVpj1pzoWh0JbT1zZlIKrA7yUlOo7hdkjpFoQuSjN6f+c
7ZRlKLzQGkAKJTo3YKusHAzzP/HQEX+5z5jOGXkfzClkIiX2pcYJ+sYrH82F
jNdwbWmAaAG2O3ppKAObF5u40QXIwPyZH2gR0Smwm/V3TyyDjluPm+wv+9dA
IuBIjQ4gOBSlsc+DHAdIexrs5XPY5Thz/JE+t8VCkyekhOx3ZsjNivxRwKwQ
lHPZ+zUuAzxX7litJ6kcnGtSakgpg0bIL5PJkajKaV714r1n/I0WGVr9g6Rz
QlAoJNkQR4k8DfYUG0mYM1Nx8jANXi3rTBjR4Bxeeb/QDFWTMLHl5nEGoxRf
OkE+artE35cMF1RGL2OBB6g4+xvGItGkr9ouKXm+ElRGg5Aj9uc1xQvVduCh
5uVTOLJYPxEIDur7rj9p6GaD5M+ihEmy79hD54o0uDn1rVTaOGMwKo/Dut/r
Cl38coMzvVEzzFEivvEcwBD1K+Wz7M+zI58jJBTF1m9SYuU2Aoa0eU63cxYE
sOlV17knZ6UMGErDBT5zB8ZnUqVK37No5hxS3hNibPYPcKTUOw5dGYkJxQMY
9Cy40FVCRISdnJgo+b8AwuzN7Ex9YpWmlEchEdjOvvHaC1ryOSgyl6gVYtBg
IHvGlvo87PbE2lcRUh3f2x79q/yxbm7mAax/95tviKYscD4iYaxi7RaPQDFk
7sk0C02YWN4bV3gdOYzucYdowFUtQ7sA+idsVj7QgdWnRIGEFeQt1wbcU0U0
Y8Sn2y4hnDVMueMeZmnJH7dFwRjm2zPbF7VljHM0rFYyENMhoiPJjG2fBdWw
IkU6mVC16pFso8bv/YFm76lvKb30ZHHAbjUJ6FLPphTBB2WYqPgRffBPFeqh
HPas7j/awvs7Z5V+Bxe/fxqIifIRdZhfy0Hy/Xbkob2QK8CQR8aBKhvx6Ntf
KP5IvX0KPZSNw/IUeiuemGT67QAgdtPkaQIB4wm0XYYc3F5B4n8jtUTt+kj1
2yj9trqIB8Y+IXQB6PWYV3fOMP2bvLJf0I8qk6eC3MTToLKTmYCRk6e+PpGv
4kvI1qgBYbz7uOUf5YpGf2eut3RVeNi135cf+vKQfuEocoYGDXcSHDzJgXEN
Btrnk8l9J5RLHAZEluLUXQZNyDXrVkJ2Bhnx/joeEay9UA1yjBQKDUanL5Ii
YlPFrXFV64+l0gzgzN2OSyW+aeyWhF56gfTTjkoP2iBUJEYorH6S3gVgXU8f
JPswerAPL69mi5/2cAlpl4CmMBKXay7bCdNWwisEN6m0Ehkm7pyCWAL9sZi/
jt+/eg+USMbtTrVWJIV+r8TEmGhNUtl5SZZ91vyxiGDvJ2bY7wvGgNE6KUdA
zPP6PnlM1tg8wjDjcysf90lwjznL+dha8NPR8YPlCjQp5xRz9Jn4+x7xxjEv
hYvSMa0ichKWZPyMVy5nDQHYkKRnjrHtteLXUBiFsVglf7PJDn8ANdLGF/L1
d6bjcM6Ee/ppdzUXe+tAFsf7wTduh2kwSa4JivKJJSVzuc6ykK0hdIFZblqR
QPEp9dfm1q0dnBnDIg8alQGriXpYJy2ejtlvuqQkgs0QJgn1Bn8zCcZEnGUZ
bi3bizn4RomvbkiZ46NwH7bYOGh2AWb2mvAJV3NJA2x70HiQ02kGM2xE6N2I
5DF/7h2+dSlZEDlOcDEvK+FrGhGzMpLQ3V+5LFmtbvOSRGUnAtRf5+5aSyxT
Cw5S3uJnRw8pP/pToPP6E/J3/RV1IANJyNWKWRzWeifIiLYW0VJ9TELn4CWi
UWfzO6azQxNXIhfVrKDrf+IFZYTwqsro5Vz38srG7KtBknFcb++jqbk0m6be
wOiIdhknZnmH27YyOxIlzeuFitYXWpJ36S7TxJag1Vy8HWyeYQqMUnTQVK5N
P1N4eq0AbEOr5lrvlFZ1pCEhG+DYTo5v00OMquo+eOCaQdF5o82ONzYXenbZ
fwl/TPc+fjK4xqbJ809Tluo+/EKmbpbRUWuDXrYsc+NPNiLt6Z80JlKW/JXW
lfFodMd4w1faZ9lTE7z3TY01/vUsk7XFdjThaBXTC3bgCMiI+L2HPNtHIh2l
xEvqCFkld7kQxU7hdV/Cxb3dj5vdRsQe5PqNw31WMOUKhe8O8LMePFDOkCra
mzp4t+5VV/bzg5MhwdHkp4zMbooVunS/q4eHN86PzMatOiqgcdSOmptoPc1v
bCrcUv4BBfdZ13EepzYkNY4TKiHxm9Ufl9s6UapVC40cqX8H4fEVOjwjuCZW
78tzVukkJQK+yS/h8x3ODeLiM/XJLnCHTpp8dbGf7hPTVaDIkLERrcuEYWYO
P304vci2EGnGG2T2ScfEodxEGAUV3t3+RBwuSv0JEnb0r8Wwll6LI5k6+4kh
2UE+pUpwUklFggJM//CxgfcHra+RB5K+L77LX9qozzpCEeSpEoeksnt0eFyR
GkEqi+aUi4EbeHMXuchyDtlFEPC52QoLacGH9EuUHb7mmKLKwH+wh953Pyu/
PBG/ICcS+9/5oCy87Ca4QEGFNx9ymhKFLxIMHlRxaO9SJ9WLh97nAPUYFvAT
HgbzTg+ZXsvUzJPBQGdW3vWbNQO1j+Zbhc2ndL/ZgUugyFXGkWjo1URNh1fg
Qe6apPs/dZtesVgxf6smXDQr83rfW6yIb95pR8UUInwr/Z6FR+YCIMuif/VO
gGLy5CbzkqRTUvgIx0Dk3R8REaCxmeVjTd/OgNUgpKhKVv3kzAlHhligwXMp
KLtU5Himw06zVNBV191sZQwogwS5eJziHdCo/DgG9Gve1mB58083PzS6kJ6j
riIMgBlCQ7gIsp4nlm9j0N1kG0TF0eXsJqYX3jQ/cGV+MfMjYUXcsnnfGn6v
Jhmb1NdXbdtQ+FMgO1kQ+SeB9M/tZfPXJ3fd6TIYfxQPV9H/53LSceTKLIg0
zVZ7/mlhqABKs9p++1FQ3eQ0feMxahk8Xfr33Y6Nrl8yUEqpq773ixYvBIyR
OKE7f8wakXD1Uy4Nv3dLrfL/+dHlTUAbnTrAxWc5PXhkoE64E66dSFv24zNs
4DbGoxXewdER+0sgTR6FJZ/V29UNbbeKPeECw1c98S5vivztvP9cPWJEQfdW
5eisNffrvbHP7KhHp6g44QT2+Z8m0lHyYxbwz8ITBZ6zk1r0Pg9R5YU9013d
txa5eXrk1/rQfZt6f7AJ9rhXfUo7VAHRw518FzKYAQx3rN0DDwhvtdQKtk92
3Zta7FljwS9Sz3TfagdZM8isQdC0aL2NozMKOW2DWzrcbK+TnMi1CVtoao40
YEf8xoQYb2BrJfkUUjVW1EnZMYZTXkX4gtApww1EPdfn/dv8XFb1kXHoI2II
QeM4MMTBaoxL4gpVwzXEH9gaqeE8EegwS2LNCPfRnzlbnUmg7CHeU0ZAuam6
CmSb0XBwEeRcT5SzN/r24GEVBdCqJtSEzd1DB8XHNh0mQ+eL8Nui3SD1VxrJ
utQfNpmr5k1hZHi/eQ8HtshuV8KHPPWr2S8eiM6DZbJLLJZ46BUlwSP+X99B
3XIhJH6b53THhCfwqoB40VOLqMimMNBme3BU+xeoXXykXfJrCie4tTjyybyB
RqO45F+lZtZJ+giDpsK3aqfhgg7lJUa7Fnq5D7P6rGrLfidXcy8V4c/MspSa
rxYbILIujTlY/bZ0j55/H54oRUFFwfnm48bAYVW6EXfGnl3dGU7Igd7XdVjT
QmSszcu0tFJYk5P/JxgnRcMkrheoF4+ZbWzoA1WQhLLoyB8uvNW9M2SDSFJJ
WJxFSVIa/7/nF+GS/Mn8qiMjAYcyfDVXs++wRrw89+gcCjucXz6nvqjeJLVe
ddmgjHXapZ95EZP7vMXMluabD+1d8bN9HN2LmQLvW2HrB8620OPH9xCIM4n9
brL2aWrITCWNGySpUTlee0AuHzF0Sr7dzxW3voIQCB5KmRXg0btGnpCgwfBn
TC1czBMMdvQ0e4K3SQxxvjqYHyV1g+dH508vYBwScOr9nQYnNab07LTAWuuh
zuzQ5X+gcFF2Z2E5HoOHnDY2Guuz24GG+sIsVQ5eyAktDJM56zGfLp9Lf3bO
tMJT08WiKyJ/xEIMIbgiCluV8qKRcKp/bRcazTngNC8Ys4s6VRVT0ihrceb+
mhW3agx+iA8PgSOPmf+9OyLtHNKbmWe7vGCIktxyHCglK/oNJegY6WhAyPVW
jTbQJ2TOWfLGT/G7Zk3v3lHXOXtCmC+K/hqnPnADQku7EpuCyMPhbNGTyvea
9/tGjuS7HfgO+pv2qhQi895eygvM6Zo/El8+lw1Ya/egJrWB+OlCvGpuejXM
S9jDhCmRcCsO1JXc4MIo5fexCWGfTIf0ZKpZhz/rwjUxGLA4ANWLO4a8z5j6
/R0VO4aRGE2T3PqNexK6L4r7NJDMtdCh8qFXSvEzb4X0G7BzpBXn4qtfAeNS
ijozgdQ4BEcLXItE4DWAlX18FWapl87i3f0QaNsNrKm/Vi1ckqwkLNJCVtBz
FtCeOVDefTv0GhOTnTWCIbDqrTKMZuJcERqHLQz9DFZph/YYyP4vkqswErpD
UH72ApEzLMBHts1rZccvoN2lFVaucceWOgZQwsaYpsEzyRN6+suRSWVBKeFQ
aASkeA4BcmVQWkbmFhtyd//LJ21kCQMlVhddDYLXm7B2uhwDk3ERY1RmSxLz
Mha0AMTuMp77gU0Im4wzSGTXvnYnsxjOv7zRIH4ep4hTKwH0TmZ2urVhb4TX
V0/0mFCrlUBbj9oSZ8wCJq5P+BjY7IsREZNymrxXgGpWtqIYc+M+zbjWbyeQ
PQNN4bQvWBUJ7dyBQaeRgXY0RfiXnq747RZg09+gs57MBZwqsLNwaevzx5SI
lnAjZXjxTn5dXu3e3mbTDg+q36V9ss/C0KOmRCpRhI4bq229JhGqRKvO4FD3
ut99ge6Mou2NwJDyWzcl5GcAMtxozSQXRU8lBwEn+KhJVVdMcMpA88NiVYSJ
Z20Ezr4ZBC37tbCKt+nrFRvecTKanwu2TLaTu+ttKU2Np1KeMpbkgYdZCHWw
YUnjA89YUFH5poL4XvVI6XC9c5MpdyrMkm6YlX/tBR6ilqh+YGV+zcqozdlQ
6IVsdXSu4Id73SJEtSZxXKtb024PIENxNXd0vNWX8685NHgQPSUNvF+Uy2O7
luVz0nDkfV/aUQQe/ImDa+lXNuVHaI5m1uTIIFZqTG7/x9oUZwdjXP89Rhlt
y4ZeK5InFHfTk+n4PwElnSO/hFOrxzCI0OfCMn+1osOWHpW8rgqOrMlCaaOe
0qbj6zU3pSHSAgY/GglaH2mu65jjG4k21DmRyovW70IKoL/5ruoTwzOnnIoU
jgHgrYg7mTIuwNMawwP9/7JGteOiNQgk9qPDM5hKTvLBMPeDcz5m9kOGux+Z
bs8/N1Aj3HknJxoHHblcWZA5NN/Qh4ODEx8weaLVzMhuaSByPMlQ0ii4ykdF
9LutaCwTsSgK8QRiE+27OdHVv6LNoQzJBPBoV1PF3HXz6h0tU9ODO6mpMIgf
mRhymjZpGGVFO7vwJgQBHzrOFg5NTvpvAmaGc+qq1errHPrTfXjneFUHLo/5
lkf6msNOCakl7TOninT7HqV9yYr0fRvubDJp6xQ54+1jirsSuPwjSWldyxqy
n2e4yEq0XFpUmWqOZTNrb2uGfzcMX4IGldcF/SKoH5wKryiQGxm2Hh4R2iwf
JUdvRrgL209Pl//J7+aIKZ5lj0Vkajcp94e+/HinBX2059rNA8rUujYRaTqq
CeJd7q+ihIUTRjfGf2+R0berizmkta1fCyv6WUeAwQPcMTCe2WVnFhNnwhnQ
HPPzoM65KwlDb9zd3Lc65VSMCyw/osdAgPVHEt7STj0aJdPAVV09DK0uimyR
ba8804yvLWW5j2VCz/GR1sfWcnXmKHzOOzdqENC3yavLjBl5cEr3iYA7qqwy
h4TC6uU9vHzY4AL9YeLqmHOY8h6BsE2iMtvI5hjbopyboaTzKf9f1jCxt4NQ
H//IkZYw/L2mFJrTG5re7far3VXijjQOzOBAmyK8bk8VHqBgjRQxwc+zrMMK
ktu/ks3YozRgl5xvjrPIL6E4lRrAo5B0ksCC+C32ZB11CBnGfQai9lJoOwcY
4apQ2wVZ937be3Zy2HGwFTXv9AN1rXRICMnwCW4Q62zqhSlx5ksJPPboO2rQ
uJysti8TQ5xiOkKefXO0iPxAG6EMTolUZO2WdMBbda5ad1c+SgkllB3CEcGk
nBnXFiQmSSCclRD3Y/COmPAY7dzKhUjogtZQr7yCgqVfPjSjynu3H34IHst5
d7u0tPKWafbgsdlgtbY6fxE3g5N073l6fyJjwiZpdn7outDHFMR+i2dxK1vO
cMzYJz40eQ+wzdUiPe78sQjqLLf15CAYz0ncnivD5UDORIwNbzOe9SiQoU9V
FWhGSCKxL9XrhL8uL2Vx6iw5wngyChsZMQug2C7JsVWzLVOTCaH+sTYFmcC8
Na0nXzHb71mPi8wHAhhOVjKzz6E1vKhtDPcrBzGZgcqBC5tIUiPvGP+5TDci
8uUTmvL7+hvf8MAphd6ELmx5wfDtNYs8mfuOTAl2qTLTeDcFXWHQWu3c/zEW
sholggoE7zXEsZxuJjJm9HDHD66kD3/k7bfWRdCVMLgw5A/esuNr0caci8yl
L2NEQYOLniVsa1leEHzkoCFMyZ1aVEfD5XhyEyJW2W6RIMkhNLJFpcpqD/ht
10FBVSelHXBQSLrJJolw7qBoR7iGceeIeC1p4Jx3XRQmKrlZqXvcOtmi7cxe
yS6DO188AQQAuq2FbPuOePc3PIuZOruKFTPgJReGlFKeQ6+23iiHWkqdP8Vh
NFPDlNZjaQI9A0GPfmCs68B1/CKsY2zxXgsu4tBdsttqSD9GR5doR4Shi8j0
3ZCuOGl6Smd4waozJtS/sFKWoAZRPBW5yA9FFWYscc0K/WP/KVBI7Gm58j0Y
XyGsKWJxkN8NABUmhJKwUHWjG2OjBfbydO+usmjNhFCfTqYVqi09S8/RU3yq
0tIScMU+K1Wi1xDhyqzjqalN9aQ1zTCZ2gMBJHZb3aIFNqXcQHYOPLKxUZ+T
hos6xaD+b3av17lc3X+EYpfojJosUZDuFo7CurAtwh7AYKnZv6gxNIXAySvd
WxjJo4cMjKSUHqOyh05D+LCbet6Ozq84s6pc0ttGI83McSuKxTLrKMTJmL/p
vBEG1+Ci7R2V7tGD4ssG/u6s9x41kRZ36jtF6z1wtHjrVHwrrFMUCizgQdPE
ahnplNDSekmnRcoUhM6S2QCtj1Gq+pbp61uGm0PRuYZJ0BmFk3SvN9GvdcJl
qYko4gz8MbqcOXcz1Y56qTVom8aXx9pOlboenJcfmspDN5AU9ACWfvsTgobk
b2hrrhVwnvIbLIYQulBKGXTz0BbTk7N+7IqMgZWFQ7zv90H6IHQkIi958m60
qTtsjmmnZCs8B1Ymur3ZLoDehKQv+eBcjeIttMMdZ4m+9tEEf+CeOehPrsZc
MoYoSVVaY6LNk0et09e8VLS2hy45oeFWDzYHiI7CcGcPKJmNS2/cZh8Iq1IC
QzOa1cXadAPnsnhFC/6huw/8XgG0qC3z4UwLUxkUCgiIK0feyOi1AXepVmAO
Wl6K2M9D9GWYTTXnQLd+Q3W/yFjEpbA8oZyr4C3lWU1IQam5FuitFtux1b6n
zRUDkEjk69CosJ0zfV6rw3ZYMB4ZGqeAsy3QGHE/nhzTWh2FABF0RW0l0lLd
kZTRwIH2Vlogg7a9rlnSU5Fb7EMA/WhYQKLJ0wFB74pB5kuCQqFjifxc6+lP
b9jZCuhFmWaE71q0xaDz/H6WNKewHSAaiw6Dfpx/3Oay7sZNaUSL4jfqNw67
hO1MeyYch7rztWFmwHunu5cKNmizSx5Z8L/cKi9v//C2qsvfBG/uhOV2wjDj
BcmqwYZExx0k5gZ5qky3J2psVmr8+bVToUBChdqQ47oGrE0y44jWYQ53Uptx
kN5gd7OB/Mr6SX2oR04zFEcsjQ4xrvTOn7A30/CwpSprCOPzNAlpLPH2Xeai
hRqlvDM3D5vEWAt/t3liiM0MU/NNpHhf2EoTM+H29VxiS3WcPuFYwbO2lBel
l8Qf78i98ZLkBTIe7+vn6t99NtXLAdC2Av+j0M/hoVisMFx8ujNrCurv+TvY
tvtJJ7iPOlMwPwTmjFbvJuu6zE4UTnckIEH0kyhMseKTnGDyPRz4giO15DJf
CNg5nIVxLx1uVaEAnL8hahIMuEOEVhjyF/sHIp5HsgBRTHWATsvkqMT9jAl1
4n3JdEexNgiturYbpZlSNSYdBe21Etp4dD97/d5w/QIv7ZdW9t8+XmjspXJ8
h8MkiVwmeFpaMTcbCDBIKb1dtmwcWkyDVH9jA7cl2nKiIjNKR5d6F+R1CvlT
7sOZFk/Mxy97R8VxO4dc0xnBTSxfzErZs4kFKb2e+TTEsNspDVv5nXqr3Dj2
YnR4CypyhDttNok2VA0/rZYYt31gdILaa4XQ4axb3kwJUIQMOaTWLiArjQrX
RL/NRG0pL6BkesagYPGTi3LAEyS+8H43S1MDAtghFBy2RR3lqmLnl8p5DGRC
vs8Vtj01HJGce2Rckb5sLit4/3KyIF/Eqele68BmYYjiuj8FDthGVeXuXjZ3
qUK12oGrGz3cFEorHDPIB/6LmyLoeE7pjZvlQeaL1givbsEeUs56U8Mstt3I
hRFwO4kl/1lGVuRz9bcVA2wwHTnYlCFi7EfrMzV6LI6FV/KjRVjEiCAQKkSf
H8cRmZmMCL42lBC3P4/IJGHVIlp/hccg87U59y9NkPyuoB4o+4aWlUTZkurW
DZLw+lPUCNVt/NrBtOiprvLWsDmzMrXX/cMBI3CLho1cLZ+kUBrBRRO6SuXg
M6fCfhtW69NwMfiRZrNKTbcxawEeIbP7l6rE7pq9NI5QRx3V4tZbkcGHqc8i
YoXJrgD1HAJdatl2WfyPuuz2+8qBkI2nip8DDm+1Zail+1Ow0ECaLD5CiRXw
ydo4Hl/eFgegPUJhIO0ifW5CTIOFqcPQjFxeyl1mG86tV2236WEUtjymqQrU
pJnD4x2/0aAp4utXgEtJ9aznh2DkL6ZQKb8qBQvKjFUHYZwsg5LmP6Mk1/uG
01EsJ0Jvu7WG7qC/DstzElQ9q2ouNluPuXeIxn1ipTzDKDVi7aXehHwCxXnx
tnh0otsgfu3M/NM2K8lFaKovMJ0etrV3/XYHtbFW6qqOHb6cZOItsRVQygdu
A0YyDWRVPYlQhkNF1RZqVJloU29/ac6Q1EYGmlkzg7wz8K6dTZML/0oIw/9R
wYX2kJn8N25JSd2uM9z7Z3enB4LjZKC8PYgweQbaP0K/17F12ZjL/Oy1DPAj
qB5RSpqukVQY9PNNYmb+rIFOjRFpY/gz2Kd+NrUQn+S7XwgGmNJjZvD1d5hx
Ccht29VlEsCDsNYiuuRi8qzufoRpuzjMgMXfTuzJ8ehBMhW3oAGLI4Q56TBe
PCdS8Z00Eclk0sKceFf5nm8gNFJgYxWDnzxCt1r9juyq2Na4h7OKQ9Q08bMA
vtVGOXaaOHTd9AuofXjFEhgfjYg49xT1NQEljQXElSl5v5e0q2Ev+waKgc36
4t5OGKydcVyvq9VwvoUvdGRUTHYBM0K+aEiHR5lxSsP0JCh+x/iOHycTd33U
ayVT7L28QQEwQ4hVDMToh1aB/33yxlVmmeVOpkHDN6Q9HTx7f8MiaHt277Ha
w8zf/cgurz6FZEwaq2UkKFJ4PsenVChrruK6Kk3Vqnu2cr0ZGt0lo7ljjVJ8
eL9MpL5HARtyIMjvXlWNcBMNSQzQDFoPWRrLsXD3xILFIGnoeGpp1TUarKE7
CVU28GUUHIZ/6SVVwnxLkJ8WlYTAfFfOyDxe9aOZassCynmRt6KJjCdt4qn7
3iK0SzOPfUEHAm5QnvBk761GSLhXn0y6La07vLnF2xEDdSTQ/QHc7Lt0AxER
1rA3O9iwhCfEG6DnMOnsmep9ncW4WOnQ+D88//ZMxWFGzgtgso0z5Bg0xDCi
sKJr4RLk/6Lk/GXre0p+2a28KNcH7uLVGBWhfv87LhhOGSSL7l7aprT3D2ug
Oa7bUhYMXZzGWXShvxk8ixDqpZZu1DX70OspHA+n5qL7dR62Y7O6gRXvXrrk
EjjsNiA6gQDBY/5Q77qPu4E8a60Xp0KxJSAT0SI8j3oaTiqWEq3p4bXu7MT1
VSUcG2aeLXf2SnxR6B1Ua3MZCh7OpP5M5YXQHw+eYJFl8uLuZ2F/wDVBUQQJ
M1qPTJaUkc1NEh1h1IVkQj9rt8CGqyuZa628CmFAONt7VxJ8+QaQkzqiKaJU
+P3Fuy95Mlc3UuT/WIIdAIRONii0U5yh6EqXkBBlJZ6X7GM1hdd/5u5twONb
H4NfpdA5j2mRLFYnzbqNrFaBn2zfpSGtFu2zfhcO7Unmg+wSCAxQPmdtAn8y
Zz6aOZB9oK8UmqX6l7IxZZzEuF704kEN0WeW3co1RcUdyR5+b3L/vQhStDvE
lJZj0NIrbC8xgvGJsZ1CBsEcVzqRsZCoUnZexiXbMvIxivaUYjl9eHBEr2Wc
yFTHIV+ALBZE2R/TVOGbTwWIG+LqyF9hpcHScVfjJ0nFE2JeDdS+lZ9b0Or7
gumC8aJB9XOjp2hOT7/mnkWw0B7Qy+iWKjZwk9uAUioFasL7eP1b0iPEUYTX
iH6U0Q14K/8ond5FqhzHPYxEl4qCFPAlY3qwe+2qXdHfGrjtprsxcc8D10Wq
iyG6Sv6bE/sc3+tOsOc/1MFObxvUtqIRMpIHuj0/qN86JArNuazj+bQ1XEtG
OQVs0kHWEorPWr1V7QT39+hpcqfHyTlgjji/mnEYlMlZ7E2FDpiP3V9P+xaA
yOn7ElHg2exo/71VIhfkBykAvXzdnF/vmveq5t3cKbVrFob2m/TBFGTzuwqd
56pjlcsXKXy7exN7NhlSKwz1ATAUDefHNn1h+rB1wPZdUoLnhA0GH16md/qO
nmZlSeCxCDZfZxeRmYntPi17Frb/aXE5+W64eYOtxthVTHk65IYrvPvXbEzb
VQwBikLCurq9hCCwgrxOPLUZUCChPJ6mgLZa13RXU6Kgp+n5SGtrE42HEbHT
SYTt4WDCdQfSpyS2RllKJCCqdsJgivY5lwnVOCaet4NU9VfkKw8GTjV+IB9E
3q8PDp9A/P8fBiX4CuDtSilK71xVuwezRzn+THjGCfgiTOgkqg8Jt2MOQNv8
dW2e8r7kUCqi63HMBLxlzbOrW4fhB66UKiefBJx7YXBZ2ZqcjDr6ZCGVB1rU
YTil78YfKieyohpOfnwDLs4nuVzuzdxPnDWrLpa8mgdduEY3Tl0rLNMduUqH
VJYUOPO1JrMhFMkd8ad5uLlD/16NX6js860uHWtAba1Ms0ylOvkx13TyHV+l
IDqABDHsY1JW3b1quzyodv31nqLIaXomS0i2TALWwgGBAxErACPexxjQu4Ks
y7P4XFSmz3hn2BQe56SfRkFttJGkdl/Z2qHb4MIbUrfvSKxwcs3D2RqpTKRY
4+EoUZklwJl2BY/UYQDJufidr/eL7hahMxXdOxgi17IP5tb2OVdItBg4Fbls
kYTOuh/1T5NR36IOb1xVfs3MovtB1i00ae8++ZjRzNcUT1WVyy9wkrjdTyxN
+RlrWxZGvy1hhit2iEhbEtEGhZLY44IySc4iv08Xaxy/AGAyVwc7afJPLh6z
+WrUY+iS3wvm8ZjwaxxAF0cG9OHXOSJ8n6i60OF6rRQAa+KMOxGeBQR59Xew
CkcX8PbY6E/Tw7UNrjJ4RHIVUiHHpA0kJ7hQFcF/NrUPf1yzoRnzwjBmrd6J
SUNET2lHqVxSjt8sfVd8SpuXSpJR40JLNcOpYjmRYcVLP94UbLCJx0m/9V33
zTGNTKI2OSvOz1Z4WUQSWouU9eGufbirEecw6ZovxRiWCw2OJ6G6Mf/GUtwZ
fuHklFTxYHO24t41IhDhB9dgkQiHQ+kPCr/XetrmjdcXCO035sfTwLIqQy4T
s2I/upotzkjqV+5xzZyF6ZrQTi4RrYdcC/qmQvXQeVsNAxhSd7BcCv6GgNND
6mYYkukL5R6SYX7kerW9dyRAZm9zg0DVCL4FW0AICwvOoIEQokMaETeRtVab
DyAvzhhhAE+IzelMKvQ52q0zlUvYqEwa5XelYokwaUknOvCXc3EGbtKlPaRm
wIPSTih9KG8fq905gHu/3A0rQTOUeNOEVcduoSPg6lVv0UkBBfKK4vobPorL
v9IfLLTBRxOUj1xd2d5CWstE+H+QgqngUXQWUMtf1CsBztiCFJxC+0ewyxpU
vfr4scuaDlKVBt38W8pKVRqdGbNKxWWtLOCkBSY9tNb+8SMH1V6qEFgms5PF
ILxF2HJf1OBhPhE9ZpfJbyPJeTZThFHkZeKis8kRYxqN/ESBUF1KXRwHAyaL
hE6Oy8QWkxWnrEz1GIzHWiZDl0Z+jzRYAj+sk8z8DHFxNVqEP4PNQ15T5meM
Cwirs4zmB2J2+SKL9BKfjafteNLtJt0HVHJdXR91YqzBn0X7De1AJKx4tNjJ
xY+0EfDk3VsdxGSPmyK8bABWid438peJFAc36VxBeg6+3oLh4f+084JPN23U
BHjtluFa7i7K8zDpQe9YqmZ8T1PoCg55W12IPP1aV/ddupv0cnc9PPFwSs2T
4C++Opoi5V+78fgkuAu914tMDx+gFjXLnJMUzJ/hBmOjOx2uyU3fdoV9iPCW
BToQta6DnuGBMXcvpfhC2prEsUjyMEMfo4UjBTM2WAXGJGr6aFKgu3i6DXHk
7jo49rdn29dD3l+wU+/Ost1MqLYhnZ7Pk28NjgT/dck+0YA0bB0eccz5crRk
LJwb/cc/RxQ9Cr59qFO5LXXPO6uBxzM2Pf/5Eb0T9G1P2GZIpd5U5jMSmBft
txqBo96tdREuPnSYCrzUMzgEfGoeh8z2rZ8K01Cx8Qx9eqofix/oM4nPBM/5
rfYnZ7ML3wvUj73SuzAeR2GuOU0GGm3t/Eh0vgtVxv+CBlguEUOkQpVGLwAX
oxJsxQ4lYFpz3IdWSPA3h8C4PGEtq42hg8gXkVVdG5v8ocM/RPaYHKKVA6QJ
t6FlTeBn1s0y9PmjjP5SmKEJSVdD4+MfOmBX1f8DAqG2SCEyC7ro3Y7/9tRy
jUSV1nmJrMNJXS2A3fmFWWxPumWkDE7b+Wh2tJeKDsok+pGvySfuwfo86tzV
0kWobmncjjnThsZ1HRdXqIgvS9C5mgsbpQh0oLVG339aN9GyUzw3j/NKopuZ
VlgoP3WTvAOmNVoheLxzZ5YINrCY+K4p0HIhIlVXK4XKcR5FuP2WcQkkWXU4
hJSZnJYKJxgFBJSINtcu4PezQaky8DS3g7STOUT5xSTqDd92G2zyRAywZIzh
76Wf1twMN+j48DkIvwtE8frd3Cd0nJ2ipkW+SgKerpQTmE8I6e0py0us1G/u
1fBsPSSRsdKdVVp3mu8mMEesbwvlhWNzc8lp5q+xHTIK096BxYQ+VU9gqNqv
XsUawkIcrcIkz6fS4SwcKcvlDUOcakNIlC2a4fwIBS/noPPXWiTFQjOWYfSc
Uhu0f2YLq+u9x/oXkC9jN0qaOet4UByeQjgY6Kl6I40/72EUYROaEtF4rbdY
OLcw0xMvPK7a3aa/3y2iVokWoVfat8UDaK1g1X7rzN/17yJjFQpposPfOaam
nS1PJN3siTk9jeh5XhwYXrTvbmBcnWjjpG6NrGxE7YkZUF6LxPXiwxAxxBi6
F66sJudMlpr3NgFhSAXYMTNGxNe1qC75hF/383sTqGjER2JgSV0dMCfeZa0W
jEk5cUaCrVqqc0pCG/uhnHcdrr/nImkZyJXvy7lWdVc1/nVSPNXF1nhvM/16
wdIYPqBYBnW2NeFD1v3kZgb1jx6p3ulxdFu/sItRWV4K8ZuNgLHMqhP+gEHq
CTD3u/E+QcZkfiHGc9kAXez/SOxf6oIBX0ODL8J+8mar5r2Nb/dIgWz0pUL1
YNlkWPb5jbY52Gl0jeKWAUgi8DV47dR/NY9j/nwEW7yOBAmgdoXpRgnB7qIH
fTromi9nXmn5U7moIGoJZmUaA/y3AJDr5uE0/GXE8ESvFuOb3kRpcx1lMCSH
vFkBHXtWQt+3olgGyGN4+gkXBK+fZzV2CKRp/qjx7qIXMw+R5WcOQWpPhjlT
sQxW5Kudua1Xhc7R11zhxvYjC67h4Xk1N2xogofBzqELDZSTTpy0Lz0BnNoi
nzpRMd7se+KgRAmI0EMlFWGzghqqo/yK5Eds7W6FQKFEaOcTpSy7s06JUjmL
gHRMhhcw4UzcVJ56Qb9S7E1oBEbycXQ46TwAPLO9ucCA6J4kvZuazfMXjPmQ
f2OPMuqk87/8e9SYAwpN6gRlWMM5E9vnIxVHPxfEGmKuEppBp1DFwtTUlkIR
eT3ibYChrrZED6ih1quMmF0yGVrKUH+jDj1SrKJ7lIsUeoFldvL+ftX9y3lt
p1LU0PnhqyU63NQRp0VhsLhC8sJLjRokWS/9mTkFvUfAM/SXUP0EVXqQ/VsW
8F5oJdgxJUNfsbBd/nU1dFt24RBE+iEAEP8P9h8FuEQhcf4YuAN8+QZZguHG
F8ohUGUYUJY5PxxJnEKj0v//Sq0NOcgIi3Hbj1WT/NaYD43YKa2mGYCpZOR/
If4KwadnpbFddHL0WYpO70hvlaLmRCr7sCOFzbHjHaA3roX1kbf+NjSltKCo
29QG0lDap15MvjsRZ47D3Vxwd9LkAvwlzLB0Gm8z9TE7msM+VD8pVfLyuxT0
v67ceO3KvUVgRmo5XKz/DrqEzNw5x/8fzAE+nkT/74gD/luYMYABiG4Z1U6W
MS4eH3V4FNFOA3HGQv5SbGBWHJ1q1/+Jzx9ELf2Zdp+LwUnm4lYnoupTAXDc
v0yusUGH/sM9Qz6kGJQ4H+Tt4rIGHssOmE+11qa3nfrYMUWZvElYgz7kv5Oz
avezftDmdrkyr/LEih0zY8DO0bkcjXdCdoGTqEdzmlJ/p8aQ1Yd6ULlxapqQ
E/sB3iZV0oLkF3Mi9bSxxjK3l2huTHtU0EJElXK28JYUr/YFhIziyL1zthB/
yeiuwgjH010wodZqapXz8ldkEriui9mamy3Wd3U/oMhj3PfG8JLnYMPUAtNi
KH8hTjwKEUEnf9rWuVbL/eFJWQVqbSUJMXmgYEl4s2e3lmhhJTHxWeUBP1U0
CXNAdzbtbYRh4S31a19jr6jzmesa/teG/R1FUyfgePYDuS1i4ErgfhNHvkCH
9gxZ7BjfdeXvHkedLnmLqzXQgSJW9zOjfpaUShsLFpQgxS86uyxrDZkEFpMl
qRm9jk+In7coMG9sGXP1L8cLHzDpNtYvVbE/yq8CaA6Elzu1tGpT7Lt/2NRD
Xg35MIj89cG5Jx+FZ2O/zU9QB7oO2+KJEP0FNKCPeRh6FZQ+wUgLKVPjY0CA
QNsk0opifv59SIYAP2B7TAb9LSEmX74NDz4dxBz0NKAFg+Q08QwpYuqKKSoT
MiqfA4cFD9UQXSPQAk72i8pCF5qN+JjGZmw9d/AoCSkWk+16HpHMCX3gmrIT
woNxMFoo+UUuTXVj93uu27h8xMaVMEPcYhybAdCvtW1mKblRnlW+T47uNWhb
y1JSNS4t0WCMkXBANRlPkVFspy2oe3x8nwL9tbPM6X4Zk+QnMJHQrT8bkbSR
tVGrQ8VGCx6XFay3yNVxLPF/RxotZ42gX+/z0i/L61na9xwkdDNyeTbFn+ld
exmi4kggpNMeLjnEvNWCWuMYY0VdbMT3INrYCJTx3xWXEaYjY2E4P82jy0gK
XyKCFIxnkVEYLYZ4CBSdNmxjhTNpA2cysX5a+XfbwqOMhr0yfeS9TsKLMcIE
WCbnycZNA81TBCaQFLg2zVb0KpTBYKkOb7BnkRfTJIpptTRrIXwtUkXmTFOS
+QoOPJ1wTGN1JUjn8hJXfBUYJq6rb9w+0qJ9mwg1wKxiAYd7TBBNvByIi/dR
qaQRMBdFBc2o/kg+EgYE77I2On1dOwfo6pWbQP9OhVo776hb4mcxZqGz1wJE
yW2FlzjwvH/KUsr3I1KD/Y5UYTtQUj9x+20uKfmUSy18SrWAjrePnUp/5JZC
zAXNupBNQCvuS0pDD8pnKIPp+LucCCDKUWvpbQtGsDTH25JnQ6IUZ2Yd9+LN
xDN/0DLr1IQpBpFfmiuE9gwEm5TVstR35a+498H+aeDmew0Rg94Sh/CKA88f
6pGfm1CQ1bUhnzFtEX+Ymjx8T9USdvdFCq0Lg8F80kWoJE987/jg4+dG3ezZ
L5V3EBsLaQRgX4v1XdIy8MpZT2CuGwQgHfpoEfFqTNKZrBCwZwbQ7raB8u3p
bD5qniQw7YEfHdY2zkE2r8m69kQJnRX4aVuILWPk9G6+mqYfbXiYM2clO/Zp
4JjHfIP3rCEhqCZikP6+pe9SNCIqPh3kKmO9WvsnT1dpGwdnqx3EooofzZlX
Ws60FABUi35RzBPJOfroZEGcYF9sy35alF82CexwuxRWEJv46cmu6NULBwKK
6yJW7Dyq8c+YtjN7ADsoB0N1pK1u94sGina8loPpjh8ECsJeLTP+PPGZQo0v
1tqLhRpRBqrbb2xf+oXKJPpq7EZlltAa7vHU6fgDewpxr2wE7qcmDzdAhTI1
dDCLeZeUot5iSvrwI73wG9L0nt+y3ETULscvKUWdOxMDacpQbgNNhoSgRd1e
Us3I+3hpaU973LTFT+K2HOj5bNje+lA3iPZ9QCZ7mpDJoGIBzmZOCRLnHCDO
gYUjmjnPNeOGzePsQ7ynDR3cGa93E3nSQDaVXyOpXqiEF2yythtpSs59s6KB
BQ3DlDcQGTeVYzFJQR6+zFxGbniMwgGa+AiCORqm60K3npIDGPTn5VTuPqBx
GGStbaRVjS/Q5HJG2As8x+QCqdxeFGA7kg2WMA75v8s++RrVgH3s+yOvio+p
heWvS5SblCuFaHQZFNzXFV4GPCcZVw1kCvSO+FAX9rxkYlJ2oQIS9rQr5f8L
GYWUe50j3cJvUNkkQOK4WLEOMG/RrVwfMF3hBX9vKo7Lpq+oFvppMgEoCgd6
58D+dl5W/JrQd9AQhJArIysyBOEzwqjL1T+dPAXpG0h+2PaqcMExVvTsabxY
KOm8AYNrtG4/ODcQEQTaVHpvbo02pGy3/3ZvJ2hALhx5s6LtZBKQpj5Pvbsz
Y9DAQ1FZNYeSnTcCGlK6VW927Hp7lf1RteG9Hq945deqCk4ZqX4Z+Mks7IzJ
WclSiBzplJauX+/J/HePbpTx6HaXRWn/U5fXM6/jodC9+zLXO3G3wkzFumR+
z0IM1polmUyFmOQlBHVi3D/0shKWYWFHDaKmzFkdPJ9eJP04z5mEKXQtWiDV
lKRDcddHWbYWJKS5CgWmJKISS3mB+5zffg1oAfcYUZNciqqqZ6HUSroSusam
d88Uqs6FVZHIyprSfF7iJ2mVVNUlrexEIx98Rn87COofKYwOCZE3Komw8KHn
VcF2LNJdUvwNVykx5GRa206zqAp2CaN0eWMZag87j9mkCXaCF/a+54znJTVz
YqXXq3up5WQr6psiN+skKiIRWBYzoo+6Y499g5IO5+NV2DE48ekzApLMSmIc
5oZgdfOHu5i+tOG9o2hDyTQrNGGVM/lN2IIpGxxid/x+4S6Dl//tFngvB3DZ
NE3VhpO3NdpB/rYl9sO4uOQbcNFoeseSJQIcR89YCFELJG6gWcEHR/lsL/09
vV85QIB4plIMWS+pc+oQ6M0040AJszI5Iof5yJdK0nCnnhAixaUCRcFnp+ps
itkCz4HDkGkJKmV1AULrob9x0Q/jfIoiPC5gVagK4oLqytLd5bPCGaUEs7q6
icRmRy2CfLC0dvk5JB9GfoNIwNt9A+gc88NVr7NDLq1XTV9cVYy/MF4BPOWV
6E3eS1hPDao+2+tWuEBjRAL2Zc+oyrqUQp3zrRcrFXIbts7QFvhXIZ4Pj5O4
59KidgyhcoVnhWBYE2gRRvdTrOHAEgSeEo7Gc89gbKlEDttR/4jCV6JdhWhx
Umo1xg4X1r8CCNYpAz3sqgUyewS87q7NdlKVwCvcM2+mPgfy+1AnapgT2sYY
B+a1dJ4owa1H+rJTzk/KLx2Z5BDesSHxXU8P8uW6Hs/6EgqCPzYVwfF/HGe8
o8cqKs/2rRNw4NwB4aOgeT2IHCSdtIxoBGzlkqNg9vzGpI8Fc7OwERqlwFg5
EjbLcKisOlUvIT5rn2n2pEvpaOH3Uh9xzuJzU0YTrJnlMbnWL16EnPXMjEyl
Pd8YS35n/TrMb1O95+Y8x6B6Y/O3GKwidX6ADwSTLW61+h+eRWslKH2Mv8ad
vW0aFMtJ1BvnbgeJshnC4XZYWIg2anYThFKO8fTHV/LhPYXfsf4Jy3ssrMIi
6gRT/emY2AV1GXc0RNPPtgknPX2qYUW0nW2YTh8/ywKbJk/TZ6of97Taou3Z
WnfsxtF7VeDlyPl/iDnN9WHg9YKkGNMV+T+/n1XrmUghbHwkHPSfFUwXqvjf
Ef/6osSbx5PwYVwIx+Lx599y0J1YyFYvFf0TrMTFeGyAM2I7nN2wYOEcqS69
U2dLbAgr7mLDKLZFmiqdmcDCoVpUWJkAC43GBE9EnjN7soeBAJNRkjF+Fr8S
lttOALTF1X0j/hmu0Jmq5kPQr8hUxQeuQ09/d7MzGMVQ027gP3m9CJEgj6K0
a5G/2vIdqM74vdSN6GpttTo6HTaUnvuR83xellfLyQ2apNma8ojZ33nxhnFS
ZjW7rme/CGZo6IESzWJXUKDRcjd2+b+GtmQQoPQ9WC+1tAu+e6e/98W7n72a
w53riq13XJ3SpnX08yHOVvfskqMacc8RT5GKPpByFYqP+Imf6fjFkUWH2YqO
p5yXafwtgLsdpNSuvQ3Lha9oTMNHF40fMrwjPlSsdw+23+NgG9pbiFrp/Uz2
FiPlvcekGfsu6uuzRgBy3Vq/T+r2Iu1pqK2A5IoyjhZ7lF4cs0vCQWy9gf1k
9Mqb2dCKLZT1NU1jIFmjofT7Tv0JAbODoOLH3ndS8kJfyLwOzRG5nxwI9F5K
keQVln8i6EzxUJGWvatVfZRuG3sGjHWLD4HnHnDAnt80YZ0COOqvTRxvDkhh
av3Ys1DMJouhImdujoW5aFNEPMzP1qtlQBtp4fHKTW5NwevKIq15VeM6bp+v
w/gV7+4Xvj2XRtp9KF/oWmOAjzVT7xLUZnhxm2VxWVVRZkGFWmc9oOf/AHWM
27GKl7xBo6qPsZNM7zYRg5iKXBani+w7Roon8SG/NgMKIoY86RfXZMl8IBkC
YCXaIpyIGjpDS7iOgASksHj2Bx9BwRlQmEJmwWQ+ZLCrn/Z2s2TqXXghWy+N
IBi6XKsyBR5IiS6ceuAlt30YybLNxcwXOTen28HZDb521wpUHWoAmQ5wwv3t
+YFImBgaXZUNYhOJS8xYii979gKfXelxOpcFSZeFOK0hysT0wn8+ztg8MmvZ
/IMm7ZEmzRhbzsdrGqqE8oiUMP5f1n/VsMWSlpcYJo3bfZjMV4xaneVax0Le
gQFBBr03u++HkD8xQpz46CnNgEpCLdWe18kgfLzp4P+m03LVCDdkU1l8YtfU
c1TI6Bpppa8NzseXLgJD+5ioTZu77Hm/bDvRaREeut8saSLMbllEmNd55fnh
eoLIYKLWli/xMGjSFWQl1wowkkW56u+Ise4CydQCYENZYS5mNWywTtzyeGhq
p3ghW4v0kSLKeaAL+IxMEfAiZARCAgNUpJ+PpTdpRf6PdeXWwJxCjOsDJp41
rq+T6jtZFtY5S+dOoBIZBuvkdeBXPjRi8TjQGT0/wQf8Ky9tYTohRgwTzfww
G+vPhZRA6iL8JMftVWShHS/Cl1f2WVq5WgHuXx0IEGjBB5lovmSUmkvnsO1s
oImsVTaTsBQGuoeXnknswTJjLoDoiVbpvv0d/sjRkt59K63CnF1ygCHcUKTv
AOS092zIS6SHQyUtRtESXugB3YgVFJIZpNVti0TEAVPILssZhesB86ZDkDPg
mAIEWAetUXxuQ+w/ANtCyvzDhV6uRHH8vFEBfkX8DQtRFHNpxtsHOQyMx9JV
gUo/AtRRMFJr+FL8wAcUY6KSZBVLsWF7AeMEsExkd+ahWfymkDnJlKBoSpVb
KP+c6ij15w0hTg6aCDDB4pDW9IgboKU5eU1zj9FaHThiZ8offHNJG1fXSjW7
BXSp4b4XDZQWnwgPS1+VL+yFteBCaeeJ5+GQPh0/sigYgF+7vNhMYOiF65J5
DetfQOEQHsf7ajzA33eRJAHEBcqnt6uGxUZqvIuyZE7xDhFsAx4oILGjrMp0
xY+1JdW1vP50vhiJVvdQAyg/YBZbEHLkH3Z7Wb/qPdeOw1Krl+oWjbUk+C5v
VhjLrARrQEtoiCf0yVtzON0jyYmSm4A7WFYJF9VGS3XyQSq90QB+Ipzn4sXz
xgFkZfh58jbutHr/YslChUZ/B1usNywbm3GJ6o0YPaBdnH/OG6Wvf//HBi4a
6P1dgIZnYgsNhfbwYfie7jp2N+KnARLyi/BOoPy53rCmIvFMhc0v9jh7JNmP
XnfPloKv0ppR0s3DlcX7+pfAZKOi+LSth5aLhFf/6z2HXQZM6DoWlknBg8ZP
rx3Wy3UdBBr3kH6N3knx7j0paWdK6WiJx7bmdxEWxktk1cb6S0f4cY3Haxjv
LaCxUhGA4N6VGBZRHnCXuhWFaGUJAmQuiQJNebb74i3tBUsH7b2yVgZbnPSl
olqhjte6XwludxhP2VPqQKf7gx1+1m2L68VHq9upA2hXVsl6jytfpDYaDodC
hXqwf1zBn8JinZKiDNx0tzaym8Jn39LW5hcpv4GNHqfJf5zF3IuTqeehIFcm
kGtPsByHeD3e985mF+QvJOONLN4IetgBb3fvNt2g4qJlftA+FAQK+gsz/1ND
bBoOlUB+9z5GSc8ks6ISZeYMH7W/ZRHvSKyNjKq1C6OhtkuPYimxLFuawpk+
ckUtSIkGDvbxwG2TSFhbIYwe0v4rWXrGKXHkCqOSiBJCdwrDPAq+hXx04yo0
7OLFnorUQ8aYqnpH46C2sFlB6UBDovnhbld6hJqinLXbww920/Twai6KiA1E
tKaBgGT/R+R8HD1dHi9YGt13yupe6qpzLzB7SZE6OA4NiqsaKnfqjJmvMYMy
9hQmrwaLkjQd9KyFbabxmHSOuUNZBN5eXM1stYyCOr85YbCDU/dYSCu3NVuj
ZPaEQDzIH0UNb77h4NtMF3Thxkrr6KkyZZUGH8zZpvL4J/eunur3YNMBf1oT
VrsJbHwZICd4bUr55fIUQY3j8cvIYYoxv0O+wwl2v+CTGCcnQVxgy/C9CjIc
R4OuiUsCNwl2XkW9Vt+0228EKH4pmzF7iA4l2JpUWnIo8n5xMVXTGNuC18hu
w2tYvyGorz/RMOcn6Mow5226EMI9mvfhehm4xry0860dLdE5rmQRmX7yI0JF
fCiGkfjfSEFYxOt1I2VhQmCAx9VnAtlGsYW3POJEVdUz9sGi1Vgc4A39caqM
vm8e7/h0rGhMVSiMCmzUhKd0IvS5M4A4jD66n14/bh/8Q8BdxmCBk4cGVJyS
+kimcNv5n/Hw0NHzkwIdNARGUExRPdrICRg1n6nLZbAnPoU1QIcpYJRPsBNb
RAHb5npfLfLi3CpB23fv2f9Ib9oxBfZDmY0Ogqj89BVykcGPWhAGFmfZY1yV
gPsCfVUAze2nG5DAHDro4cOGaKTLsiBJT1aGwRwoPorT7sF4PGILT00P7ZdX
eoUS39qqbN2UJMchj6TcJcf6GxxlkvZqElUzG8MXZQeN+ENtjaGUEHrDlifU
63IRvA3WzhXBvb/7HzoRnu0TYJFe+lNV25UI9EnclQCFLQYe3MNuOHJpdSno
mh5RQ0kkvr1VshEki/8V4y0AQLC4QPrUPRno06sF4IHx79J22vrXD7WM95Mw
9gCJZQhClz/9fqP0/MC6AuzQ7+SHGWjod+ECzxBIyF2B4K4TM+nme5edBErl
D4yunilvb+smfRGzOYFh4+y+qn4Ig8+PAmc/vX7YWmlpiq9BfeRyzPf7k0y0
48uMha3OsSSr96qcO3QTm9sWNGnVYDfEP0tiandPXUateUMVYfAP8FQK4Gm5
OQ+vKedWDgI7QRp4w+G1XgvUAnlIsmo0QHLbGrfOHk4AFvOCTifj9xd1y0dA
hEoXvUjcnoQ42XZY87aeBYtW8ulboGwriOwtZGrAaEX8a8QXgpfKdhC+buIp
6aVnZXfCkOJHlvIdsYqeS4zWtSYe8sjvE9m5XzCJxQJaeghstZfKt57mAg3n
kgIG3k8zLa9kd94qLY0f3WxxTHNEJT9DaysAzkMO4FicuiramvoBVCBmeI5h
8Xfv866zOmqf7adXJO7rHwQbOz+D8DJOJ73wZ1UduKiLM48ajyLyCpjHwQKM
To4EM0f9he6qPdPk5qThDyIKYcMJkcUGk1cBCvT8IsuUBM1EtH63VNJzdC45
PbGT2IueiRYPg6EJH+PbMlkq1f3QD/snvp2KvPALx4EZTA6/BmvLhGsRVoWS
YF+oaOjYN6EqSvazkteo42k874UkW2mjjZqakzUZKgdTpv/1bEG+IWptqP5j
86CjTSJPduuMGHe9VVMubWtdBGM7mZr1xlUbr5OiYSy8dqMRSL06fk8M9Xod
eVB8yGrnisoOwAS9T5DS/EZ0zEMSEYakqKzAPmUcCLAp5c0II6us1/FiNmjl
qSWM9TusTUC34mBUcOGpEKMzTEnbf0wt16oECb3SVrxxGRzV0VZEd47Rz3Yq
4nVdhiYTdy5EKtKFcQa0hj6HJCTDVN1DVSBoWSeT4wS7z1i57tylftZ0QqsA
Nl2ik2ireWdi3lxw6jDd/d1PRszGrNdbbcVDuQJ0s727rPAx1JNPHUZiRCP3
De0vMFui/LC+9DN6sf+FyAYSoeJIhpxg34UxSm1mbROd7w8F0RpPMCC70uvZ
E2or/LxpbR+O+A/htstyGqsJg5Jtucs0WVpcdsGBXDsR3gxt/eUhOrvJzM4+
VrgKnjLwNNOelgzBjnoyCNCL4lsbWnG/FO6+/mhHO1j4VTbVZimHrBzsK6NI
GRQuZttWfcGZ6lzpoBDbICilh1KB3tror0tfpsx+K8M7XwroOu5aKwKW21Rb
yClv9GnL/6I2VR2aWkUP9ex2OEQca1uMBeWLsd2UQR5EeO9MvDf2F0EAL79+
mdK/9KhLbxepqr4vVcaB86Ffd0ZVa04TaAzE0slIiwwgKm1EXzlnsSuERVsN
1uAIB3o/lcNM8t1L3vV5OPnsinKl/nAd8J/Vyx7MEDn2yAaAmybzbJbIraM2
7BcW3dJofzDExPmwivjAyZl2G9rEx4wlRmR59Nfkeo+zkNGNDCiOXYKOYKEx
rskUktjz9m6kfTIrjnHLRa3hFsVzEqsk+s4+pfon86edKrGwUYxCbWxkWqZC
6YElqE86MP/ncGvGBswrJ2Qz3SGsojyG5DGEML96fhhxXfelu0H57/+DFt/r
SrA2CA9vmowklM8gJKQMezJnpD2Ttv0QzrR//qE6+4H3cRoMw6iGpSYTCxvz
BWSznghWz8JtBR3NiHVIvtp9oP9BZyJYkg+bX47bTBwlTkKZVeZNMoUmMOiJ
+gbt1dfnrVsMg5kIq6DduDxV7kSdA7/kH9KHDH/SvYMLe/aOe3bIKGuvA1Oj
ZhmdgvjLJ7MZGgmBkn1Ph2FG70yNMprklPas6CPFBpBGG3gbAFHxQ9Ap9dve
pj5IOBDi+eAb7bj7xRPPJXal9op94p7gC5MvHq0QI6Sm3OznO7uYsXfZ/ze1
gTvc1z5DqlJ6VzyJjXhXjWfZmWFcCY/yiC3OYQ61ICn7OqD0so7x501/uu8I
4DATot9HDfkKqD0WX1VhTFOzISru7E5EC6S0PKh6UBkXYyxXVAALCeSskL6T
vb4MAnMoipTFO9koaAv7fej3rluEu66PP3JCZ8vVCT8/Q5jujs2gJqBe4eDj
FaDGjA+8hBc8jqnlvhfiIlQuNIw4COdajkEUG9vKcY4J18Ca/HC/Hk5+PEtM
1r1IITfEAAKBKdiTd/tb/jSmQNgEKdhDZ1XkreGI2qalIallrfafORpxBgDP
NoQcz8J4sQylqA7k7RU6hVniTeN6Z5LoyV4TK7E44SRwtPluhsU/KXJim/Fc
+MkIO/ICtRvPm9598BSAMYHHr6cbjCPxrgHI3N3im0MoU52QERmQJre6fI5G
QS9eHELLevuj+dZc/8EOxTjeV+M1hntpGR5rNAhpXrMkVqJ4PyC19nBgQOiT
8iua+260di8rzb9p30Eq0k6mCUUuWPCB3lIUN7OTFY3VtwaHo//79N+LIvS1
yCPz174TqGDOmFhDq4brSl4rreqc07igBKrPvvFaADl9u/4TaGScFaHd/J57
E0A3j8A8iuT6dEWD/vb6kbT2ZNuF9E6VT0bKB/B7NMuNuVC5J/GiW37gbnQj
DDezRSbiH052Y33USFa0PqJmPC0kIIwuajZuE/arngTSJHM4ajxF1hEmpJQS
V3O0uaYGTlmaT4Yy2sH8HBH3pqG4fvjjh9BnVRXajC9ehOdYDly9ErOdEtOY
SAB/gc/xdfRWqrdQjYon5rZZdxAcK1RalmU/S5h8+MgNhFk3VECu32vdPKAW
fHbZY15lAXGfG5AqBctF7DPsPZ/Q8qQbaOaCY91NtxFskdF1mCZPPvprZjmW
8soPzqCgLrnQ9YNmnPyxdtGElUAwVIFy6sb/y4GwoXplSlnd0i2r82T8VF9h
anqujwNP8KBDKmppAgsWutKY8lEVzq+kIyXef9XJESNo/4hdr2l494H+rTKk
bHX8h15uzAWnJZ9/bef82JwuIDx0makYvDyFpRvzb/V+uJahH3iYm78GG2c1
Pmiwe8AnZ4g3+HlLsYh2uFNszMpc1zeTnLiXYBeskXpXnt83gZy1qojs2wPd
xcTWWrr7COZZmGgbBTN42dSj5vGV4oToblxAjVKj6IWJol4sg1+eE1aI8hpa
6Irv9YMEAfTl2vmKFY7l+hDIKmbDK9pZ4xqIZH1qVWVu1dJYcoJjqro+IAHH
j6LcthUj6HqVmrSZQpV2feVTi5GHSigt4MghkJ1vvQXJRXh9RHmwVB7yYreJ
BQpSjkM0jFGwMAQUVJ9Q+prhaEXAF91Ktloxa9n3hQI39IQE/mm34/whMwqs
aPmlcX+iDMqZb+pdV7a/BMk7UbMtl962E7zZ1PXnBUhOOpsYIbPK9nLOeh5Q
m02PF4FVyAReHnLYjAxbMVXU7Jb8TS8vzBQAIGRMj4be2F0fN70DPbno133C
C8CgS/jCwYXAkAiMk0dqw3amuxR41HbxYJWiC1dYGPMVzpn4GCN720i17lEr
zRYqazo5oinfTEkFaJ2xymMiv1numVPp/mGkL8OVgDDcQMo+I2GG/cxwBQ8O
0dnzLQxbWZnDcEUr6bzeuv5vzApAK8mjeL7SEQBulLOFpT6gKGDXX8Ye2XNT
2ruC/uGgoWk6wg+n2A3/BXDFXcTmWUJ9fjFw/j2xNgG9/Zrr2ixiWu/JIAIT
9O1bxGH9honaAcOMO5qNNlyimlyPkOgl4+P5rKAQsLH1f59jxFOZKO17bKmq
CH9eZcSl/KrqRiYDB/VKdYiBoCzZLMybeno0Lskk1UB7+7i5HszZthRAshrf
GpCjbAcT5LopNOyz/T/ssms4GIyisvNW3PCCh0KvrFq+NUuGhRaItdqMG67u
WlP0gMDkBXiSk1iNk5e6hUkC6yPOHFjj/ydvf5IPajbeQocNqe9q0aM1YbFW
VEfxuruDrDjH8W4HyK/yVjdBnYCKa7qH/0buCP+6pC6wCMHMggqxQbLQYaek
PcWahI2Kb0jTZjFZF8lAi5uJIf3kC9L9lmXtVc6f7/B5OsHQL0MP2/PPqOGY
wInehxMqMJAoSuGMWlMjpKNoVdif7wiY9A7f+OVGnizfXhoT+JjcTJXRmiiL
KFYcVQAxXir4yXAgCU6PirkM/x+gt65ylqsrZ/82qVSKYzCj+SaY2NF4kCEh
85qc9XVwJVSCbC+BRX90+HNgl6CBRyk8f5FpNMuZGg1P0MlH7xVvfYhq5Idt
X3YQEJH4nIUvYyghUK2rbkwKYcpLaUMs8Tyd6kZKk8C8BZbmd5UqOzpX13xa
VCN7GK533O6G+YZvhJUNXfx1eZp+AsVE9fSB2jsPDPr7B873QJW9AOUsZmsx
GRfcJ/NSyDFfemyXOOqMAPcyiNCqAoHDGMppb7ormHrPCVVeNigvY4fpWq+/
RwChHVWDIppnJBi7Qi51Nk9gcOVm6AocZ/tJAnc35Ms+9RjzN0JuEQ3TduGj
8l8I7iIIdMwInx8URkWSseMbU2XBvJy93gQdqzLdgBhCDwKmJ5ss+E5oHYuo
KKID/bsF2GHi2hxiPmNoxGsQqWk54vkhJWTpI8H1TNJxcYg1/adYNztf89MD
zQpg/OgfUKqTndMYIfujhSQM7Uj792UVjKsUMddridzVcwl09KaQfFsGO1d7
+0hw3PuUCWBVfZhVybInMlNJ563X5Ee18Owb5PqHqS2ytc+VDmc4DpnRaxoT
uZLYAZ74uOmPVy+tsgu8ciOORhtgnZVFhLc3vNG16nVl4StFCWvf5w9YJSYc
yO2vBO68dJXRUH1dK2LdNRszrsUVHseyqKmgeWrTJAvmfMTJyq8iWheeaqjm
rXW4DmOfvrc9sxtlXTRko3ECoO5zl+AIXhV0b4Hzmo7a/GpRsCpIWN5FT5yR
UWXdxVpWlphZH0wrt87e+KzYPDAGKWNCQrWr5MYaGHY9Dv7khbtNMGAVVLIr
LVDNhT4nkOy4ULR+Fv7wcfOFBb12BP2cSoVKqfqLXepbfRyPEoq0J7m15EWG
WIupOyO6kcy2hHC8x5vv+h8mu7jUncAnJT1+QGDu73e02ZwTX/yzwigUSegl
YImx/lRYd2TVQo9ZngNciaNmumdjFLcCZhslw0dW3eC43K+DK3diBxvkBaFg
wecG7DbqD49s46faSNXTzwfvw8YY5TjXb6z41ErZlkwym+7q1haVq8qQfyFM
Sk/1GsaRRXBiL1GAthjq4m8CYVvRzws+ItZIupmvPRg33dqXG5+QKEibHRsF
b3eZ+QUz2AgQy/e7iLKnZSXs6VY+sG045V3PY1ZlmF1iClGQbl0Mbe3XmUSi
LH/GFtDw/cC5wZ9duuothJFV0ulTNmBhgU49Gw2QbasofyOsquTS0K2BXA/1
8qv84dO8I1fyS+noH72KBEkBNawASpQh4S9X2RfjXwDBCjuPo2W/OueGjMBP
yuUfvChkixarawuVzwBaMnciQwo9bJzQbVK8X/K9YLBo1c0WSKH2kgb1oMvZ
kAuPU6wcezkLkd0rIG3wMaQutY4aMKLJ9VeWC9Qt4c7wrCdW2MGv9iu1osvD
aRYnTwv/VzcIaJr8xzUsUWrTDf6i76BxYD3GqKdCZqSYxMQpZ83s2YadDBZE
guxPodmWLJ+yoCtX+YyATgCtNgyDm2r8M9XgOolWnleYKli12kpmm3vfdMXE
C8wYoDbG7qufvTsTPvDETTU54Q3Zjl2iQMqczOalQaElcL+cc5bMszsarDxy
cPPOOb+Mi5atcUTzogtq6tLUfu+VsEbZU6T4onTsvSE/J4KVvuQzjpEJ+Wdo
qDAaC6nT97SXxCEJ/XxVTHGHfH8ivDNrMIbYrPPPIxZefaxgzLXkf9edF+Vz
sNc7eX8qk4nYufjsjVfDZmQ/moWrpGzH7wJPSPMwRRylqUuEAe5NcIevW2jt
Ic4DqoGsfFfZjwi20s2JtPdkOt1F7axc6NjMaJi1Wc4zzeqmCUxnu7BSp/IY
nkjzy6s5mG+SJucJaNCPQIWPmtoUGIbp45+zzMNGD7wmOUQwa/o/NGmOm/xi
0s8W6cHe19y3+PUibx6P/NcwXdchIox3i/ie47eiJfnLjAtR652cZTYPN9Jd
Y7cNq55NZsKkkE4Cec5aIHO1aGBqOqu3UEGpm7mH9Itw7Gk2PLY3T0+4V02F
dfLfaDyUyVobT79m3AhnDEOCqhrqaYrmFjFpadD4vazmRWyZ+BRoyJ8e3DBP
uqU8p6NChCIAI0A0Pm2UpDRK0IJ+2ph3vuONyUtKvexWfHOmrS17l/G6aPCo
ISFHOl8Znhv3Ftx5ydxC3WSKOijY5PfhI99xQADpH2apzPtkhQtK08//a/VA
tO//PLd4ly98Kj8rhb57uStln2UOnURXALZ38i0yfBrDIofUSUZRIVHaCC1w
nbwWVIumQmPvdfh6qvdz6DM2/NO0gCairK8lcSKhmkQCp+ACO14lkswShyFF
SPdCAnpmaKWOPeIUKE/l2FAfkixVjwQ9MVjN9nlyjQ26lwVm7/7G0S3EGBPr
fujlWsONKaD168yhbkjhkZenn/EGL0SkcqcDYTzgPGps1bmxNUPVtWMRs0QG
wxmXb44r5UVPNCrlUDEKaDHJjeXnhaMNHUyI0McgXH0Hbm0MCdPE0ps4b6lp
sibn9x3ix21h4FbUPCwIIlQLzyWBlDPD10OgfNSq13eLtlvuk7nOlWOu3EOw
u8qskycoPlGK+syLB7JBgF3NqSIC46r3orXj3sPrsd35UsZxKetEcxvqUIjB
24M2Bh2RIOJm7ump05R81lrJmIdTjPfKAOjXkiEwTTupGUdbO6pLToC1jYMD
2RewTxTn41/fRj8Tq25VIgU0iK5KhvDOb4uhkIvMp8t/auBymNb6NehIKPTj
trPXnEZGP4GX0wetRFJ/VwD10C9ISV9yvzdWrJ60rp9ofiuwv7TzoYx8RvaW
eH4OwaN3upCk6jco8BNeSxPkDUDd2dRe6AqAt1/Xe1FVB3PO2RQ5EJ7u7VSF
6R4D3STocehu/OAb7qfD0ckYgV5J4oR33a5y5bn1ltLDioHKB4L4+7St1UMh
aaaRXB9QD569PWkM5hOR8uH6KFNHs/ylch33cszMnQx/o/plNtJQxx7b2k5K
fSFDkKG3NCAnXJnhYxZEkA6vhBJftivoA8XoFRRgVeT9XAFmzc3zLVsgij4v
c7/oyoQfKxqZAJnpf+cRwEY6zuKL6Ha4vQDnGSMquC/T70xh2zLCiX+t+xQl
S1Y8OpN0PMyy88FYy3wwbJch7g1M0QansyvoWNo+XguCduNiK8q299CbLY11
yRNGqm4ma0dGgpC0egoYWXrFXCwqbxtGKP5lv2o8zFqJ1W0a/7+13M8lJQZQ
3adNVlPExbLvudRXeriXiKYuaKc1KYkrO0B2itr6e4i9E2LYw58C8lv3/P5P
LIpNId3KZBSS17N3RFzTKMLfHyBLhR3SpEhdE4RQxmX00nh46O+udzT0PHsB
k88slISgX9+DgvW54vS9ViB/FtIBUD4IG9FsYv/y254qRhb1mIKm7grRT2Uv
72kyQhVS0pl5D4XqoC0nTbyyT9nsx/YsseRWwLDLkcpSGP0iDtDKFF9sNTmd
Qg5xdYfpdOOOjVTVS8ZEBmJ5gNzAj6O8g9EHLG1ikYnTLGYx4D1xbf5bGcAV
TPS/AD+JpqKGRfV6a04D9ebiRgDw//uL+IX4wORl1x68nLMjZIhi7v0zSy4j
r4zC/BMX15fGz5N/OeNOtOIqNwFkCGY1VDvDdV67vzIAH45zVn0s5g0HGKjN
3M1p6ftDWNvBWSY7/HVgWkY0HKpk2qfWGpWZV/EJrQJCy66Jkwgq7MBxHDO1
/ro6YKZdnCkGKYNLf9KE4H4+h1SmRTUiaYASiXvebh9kQfKG9yUsX8qDFqXb
iHaMZ7oAWBgMq8rsrtstms5XOh0HiAn3QsjUdGDO3/DMj69ZFXOCvRfcRZF4
xqJiNeLJxNKnT0NVaAOnWZg7VO7YMFOYNoNJ8VUDGjBPCj/yPk+jxinKF3vV
Aim66SyY382qcV3xuyMuSCm7yPvkFjaA513jqF6dqC5WzDEHuoxGS9CUdYYk
Zbh7md3ks+0kegQCh3C/xn4Wa/kmtrvbuRXcReKB9BWYD13rwmkjYqbLgZGt
cKlkIY5F2GBZxuBVOxYOK7ISD0lQKNSS5Yko7WiguIvVmiaJoP6lSxokZVAg
UGFEFevOxjlG3R2cztAXqqOeL3sQz5ZW6sEwnB01F0SAOhqfrx+JVYQAChP+
z6HqEjlLLylq73iqCxhJQNrn69l8SnBm72XXucLidqPH+RsE28VWtt+QA7/J
oAj48wBkVGlIg/toILIFDYDhoh3YOe0r/qfjMT8M7TrxYSDxhq5N0mA0+Fj9
LTdrHSkZ06UMPGSDwYBkp0JI+9ICwRnwpBvAIryytWPsu6t1POWYPp5fH320
9V/iGvg/CcXn1FkPMPDmRQri+xnHLHcQrrTpcBXAoytRVOXCzecacgVD39V9
HfTdjKNTFKREAPxX99h0NmiEF8vAbbmspSsMnyBmlKV0FT09J33eSKw3hEWn
40stlDwLvaAY4ZxF+QkVdXAZbm+SbZPev5POewWmeZa8x9VN/cxnA5Qu06n/
Lpw1x/KklB7dCkt7n+FvC+f43eeecPKyCikMCohTXHb4dzjo+MaDU/QXfFkW
VqZ0KB8QnNNC8THtsR3eXD5RhuOEplR0tQUcDYlriUKGHxFcoPbMtXJcQEKX
hYjdYCOczlO6rZrM+VQTL+OkBU4Y5fNsEL79Ws1+n3Eqc8UqyzQpW2XRHq6A
3r4mmm0qf6HeHPru5gABrHiGhLg02lj/PJTnfPz0TSMD/+FcUvRcsWAu1klh
RER891BNH/84K9V4TlEqvKsBkioJB8n462YWMAF5UZwdFe/x4GB60V5HnXVu
YBhfTK0RBGMK/1OEn4HUA/lBuK3roq2KTsKwuc2WNQCANWEVQssMbUMJx1mj
W+mk4FHS2jh2wDNDkQ9qbSKR8lMhgrxbDxuKg5pHm9gbbxZgGgHmr0hmYvbG
jX+NxBa12Hajjm/tXv24PaMz3CZpr1tHq+6lrFgVfjw00J6UHqommD5xnjCY
nTQqHGqilCvnF3Izv6RwrjX5RSJiindLkjiJH704+QSZl/Ek0iu/zM1kr6Iu
BMbnD+tBDHd+jh43PkBo/pdcnf1VoFIlkpMc5Np+MP7fE6jPLxakPMACSN0W
ECK3VwVgVyX3GMjEMALkxgbkxIHRY089QQjTXmyCTpbp1Iv4SeR55p4mIgr6
EfXWOwWsI65Td3baOZQKmpeZI60Mz0ocCxTYKMzCvAqpKI9lKfgjtS4Nhwvd
0VYDIHIOvISo79XI7LXnGQwv9j9mhRYMyQnajDa6eLl1Ju9voxsc7y6pUFd3
dphxcrfRdXsKAKUjXwXalPF0A8V14HcZWT34hFhLKMm3Nawyao+/1ugY873M
NrK7qCvxsB5UsT++eFT822mWRIyJF2Lwm2FI+bhqbvFwwD6Yyc41UT/43ecf
5pKnT+DxJ6Ak5vno4vxrmLRtF5BgPCpTG4Dl9bSKCzgWG3t3OiaJpqttaC0+
HAiP4r1fG73abP7QaVO8JleMx+NSxDaTmz1r2uLDXzCKqijoULCvDpICP0DT
hMs1sYJA66aNK7pRx7zghFpFbSGofavWhjXRJLXJtPVrSjVpPD0yIAREi5cj
rrp2RWu7/BEcWuvUhfyQYzp7PPH3Ex89zEI+/gOYJm2+cn7IF3r8wsmzP3x1
+F4yQXwSvwKqhIHidzF0WdX/E6I9sK/+c9e5tiwFlbiQmfw8yB3/M0dj9kpJ
ma71xihoOCSBVVJXB3jzrwdNTwnPNctnMZrbXC4ctTetK5kczdVUHxUKw4s0
lf2V/l/fTi6DqbJY6IX7K7Gny5/S3vWTJHxKattT8iCbVQZ9ZmyLhnIxzvTH
s45NTdx8l8js9/wsiKfEZjYOt6KgH8MIjDLd3ROWy5MRdS3cFKBcOmfUrC4G
nCpFIj1BSk6mhlmrrNCynPB0sXXFD16GpxY8O7PsZ2KWH2LhwvvcKK+pAmBA
nnR1ygIlUZ5vE0gTnn+fef5Z46s+1m+IUWMiDWOCi0SQs/SZUiW70lE6vsO4
xS09zD2x0N2w2qc9ggbILfRZ+4RaDYlmZeWyAPBDd8OyNYJLmrI71h4/PRLh
z0VxtPiJDEp+jRG9dY5lOzorSXOGpZepeXdaTnmaYzBIfuRm2QHGKdlb8XAI
Id7+e7yDrRlTq8ni3cqSUR072YdD4Vsu6+4SGO+qgGtCZuEfPx4/UYuxaOwP
I5R+dwT1t6Ghg3+lHJ7eGyNUxibrqg691I/AxCllNCXu/qYO0yHGKI1jDvQl
tQC3fiHZWWzU64es1ell8tB472/eQDpTfRBpckgoNze+yZq9fcvk6Km6GB7U
ratsz2nx9/3hEVRhNE/OvgbQjXM4Q1QoH4KI6QAkpZC/KyDAwPhWgAxihEwt
w6CiOMJA+iw8/MBl2NcmfwkvhwUoafLRlG6uudPJvMvyrxmHWy53cS19KFPR
oHYqmGq74cQWeZElMkLwnHoCvRNeYHJydda+qBvxDjXh4fXMLg+uVha9SnJa
d235b666g8DYtrQWSqfJ9fXa2XZlFxIiuWzbiCzh6N5qz3gHTzF2daXnOH82
LtcAVQTYlpEFSW772fHVAnmmYOgt/3vFFxLvqyNkFQ47hM8koTh2gGEjvl9e
CLMcoEaKKveav9AnzzOLRDMrDiUFBip3Jr/zjoQ/LxisDkaZMAdIebGdGwCY
MrvHtC+MMjdlUow8CdIps4zqqgyEDTWN63MEIdqGnNd6SBqIYiH5Oy3L8PsD
o5F6rhpZ6gw4XbrYZjuOvpviEJmwFaNoDVA3Vg5STb/91LrLiNJWSKTLf5MK
3hA3+zIM1BhnF0C9XpGcLkuN42/IpmtU5ZoQlSbNG3M1DPn+g1JUiPiNAHXE
PoRn7uXM0xmqTi+cQDgdGJvvKiwkLg2kY4D5yNDCjH0+tD0W/q9gMu2Q177m
kFSUIoUOtFhA017F9eF+8uL/V/bRudxAQWbI9nF8UtY9apR6avSJrN/pi/l6
j3wzV3V7AnmYhce/wosIu44hXPkEbsUJDRIsYpMAA8wmjMHMUYwlbHwypey6
kG2OiqbAtS2UPE6LdkuDdwvZJRUiy4QkUpqzEk8h/+ErZPgBHpCfVVShMpXq
lj2+YrJIPVjnFm5DP8tlcr7UML/j51GuPpl1TdGfUJt48QQNlfcy/LnCoQ7B
MN+LAW5s3gMoelCy7o0eyos/tYb+k1qgF3PKsKp2wdLOeEwTHtp5CimBWWzT
KmnappbBNOxWjgE7ET1CPirtao29ZMsnShzL0esKwAvR1qInGNO87wRk7yPh
e2x1YsaYY84Q4DiN0/9JJq9piuuEMBQ/22tL/qrciEsd7XgchQvDn/mQtus5
I14/Ciz67mUofWp2C9JpjiV7D2KDrAlpuTPetver1HA+tVyouqV71Yz9s3m0
itOIK03Gb0Nlyo/U5unEBqEqJYg9R67jT/bfGVQj7Aw3NSQrUdqymPsOes8i
04YRyj2+ujAth1H7IzBidPnVYojQNkbhxBmclSOc9C95h6Yupt75NGy64cF9
3seIiOB2uIhL17KGpguvuK1tI6Jdr4SvQVubV+uJbOr8z74imBLUQdLX4XDB
hOicihOmvQq3N7gBd7649aZBr/SnyHTePZRBT5XbdVydEkzO4mrmYbWgkqBr
iiLa+TqAelWsWLIZcXg8ZpgMWgxr9sLcc4t1w6wNSdXq/gkMieeqM0DCtS8R
oeZhdDmvjBDP715Z/wgBbXXIIK3lZPupQNE2osVLrUEjZPzVxOPQos7jDR7B
x9pKUT08ax77e3qI7S5/QTC9K1jcf8AD44l2zaU50fTmkKAFt0SPepKtL0IT
yYrqRy533cmEmKwRLENfWpBSUE+9oitT+iiT8Y1Y+MpPDDxfhFN47uA5OuL4
C62ZTztAaFNH4wHNTMWdSOYJf2q+XivlQfmXV/dIHQMCqNOks1Qmdlp4gmtV
ZQ9Al4kipOkwQH2w7kOAwg0BicPXLtML34ksHskta+wbhErtyk9S9l+u3uRW
vWhArUyHQLW0CAjF+1sILLlCjlffRrB5YsO+8nBdWekIBLb+1t3VbYsliuqB
0/U2gb8CFfksRsiSE+ecoYOvXPSuVqCHFTx3GLIDm66xJhO0W7LrztMrOULu
pkjj6rH75B9it0894qbqWo+btyzOLTJfp2oXPWSnYGwBkJr+hvufIIqfQGgx
BhFqPUtcUn9Eok/9gPsO8Ey8LiymKlUBqByd5luBkRODgly/skE4YnLYqrQE
DpcpIkZ9+yYOMVIsj41bJDEgVSvFxzzR+G2RcbPxoOvz3MwoqVgOH4XwhGtD
XKe5jYmMf7iUsn8sgA1kHxK1gQwgrvvRdUIZvxJ8zeKKzx54N6gz4t7otuD9
69q5rEJVuWQMtWwbLPJqO9dJvV5UT5O8XWtqkPKkxz2V76g02uUoYIlI5aZt
TjJwbtAtVjE4hrOiRmf/rLuaKMUkM+YJPOmCMfrD7ji7ftznEqC95zv6l3t9
JSBtmB23CvCGHCvNWirih03E3aBnknsEPU3nVYxVMVXKrKW2T3rMMn5ZEx6D
45pXDQhz/LzwkdrzucLUhW8vzeBMy80knTwNfd5r/dV757QKtMiwofyhodjj
2mWxD9re3+SQecWL37AmZw5uw0gXjBDV7OC0f+ZIenA3N8jmYQNQjQAgJ7TH
1WSuAbPJK2+JpAJbyDteHRZuNpeXCEEkfyNKupa1Dic0q7fGiaQWzWS+fYPp
YBHCUehKyHxq90FqVR8Q2mfpI0LLZiISNfl6oYQIyfDFuBFlXnq1lH1Fjlms
gXmb4sJAFQKZvi7GPTdu78Qo5U2uQ/YMs/MRMEoS/MQjHtbDSwVklqMg+Rz2
IxRJ7U01lPCPW3C4RMUcRnA/J4ZzvDjoMDvV9lUbtmksGH4uj6t93G4uUq8S
+dD64CUbNwT9pgXxOExIP9ClFOpY6mJir7GPn96u+XGMzvRaUyVTdzw3HztM
/4oTgei8Qx9cRooiSmV9rZp1S+WvKDhRBorWNU+zOT5RAHSp7jifEoc0PwEV
1bN3gLpyVUnLnS4yQezNwxzkf4VEicM1fy0r3leyjoWg41GvmxuDN5/FLCqD
x1buHoKpVHwsNtPNWLSJavJldwET3cMN7ku2N/5N+ZHe7mFZ370nPh4Ljyyt
tfJCp8WLqL8VVJpDMm1srF/3YzrtgblLnPIpe7JKZaOX73FPoC2AAKXGTpwO
Kxm+1ZFQHsmTHkODlb3LFF2jIS9lVlRQpvvT+JxNoR2WPuKwjF2Ym7B3gI8o
g4sY0FjTIWD8sDnIPDLMlGvQK/zG6PnNq8TMfxp3XBs5MCSzYpnM48Lw1vho
z7RSeO2unfYxgbkoq9Y+lT47MDyU4Yy5F9Rl0QkEkhHuw85xlufZtpizrCEE
m3bcQg14N4NVd7wn8HIdRTopsEYWja7zRnhP0Exy6/YeEATmP091FeSsoLa5
UtiCNl++XWLvGhyDCaVxyiot1nMeSkBNF74UcjtsW7OcnZTrpoXpy9Akzsx0
V6IdWpJKER2pqQyZn46etKFjQ27cj+EKhjP1RaySMwr0heqpgVnIElxY5eaf
aCtXOKgxxDT/rwiY0t4h+lA5YF2PhI6HdgbgLJvIYo8ydHkh/vPQFLOTFqCb
lW0xtKXjbMt4ehCwvDRtAA2oN5D5J42gQ3XgdX0Uo6Jyx7RJ83XnAJdF9KpZ
6mwrYUXwP4w2wVw2Ie+IiSZnBlkNimNTj7nrJhr/rNNqGhP7OJp+V8q1FJ9/
4m/r3UY0AXnS9oqgxFg1r82wkRMUSjt7oTR3XKtinGkt+RC0zBYSeW9gvNqb
A9+zTb8l65eLIQHY0Bc7zJcKR4AFAz6vxdmPQDkSv75a5jnpV5iVG9mLXoMR
crF5hm54SHv15Tbn0M1AmxvzIEWoS3eQ49ctqJPdQneOKzzhIkHCNqnrZSLo
xvrbF0WgdV5WAJyeecYrGFrCLoOzpqJSIsrOOTtHSVq2o8BQTndiZYPBeJVT
P+tpPEtgjf9SyxSzCZcnbw5t/spvLNJSabf9VKKgBL3+N4l29w0uSbI5HSPP
I5uiAmY1PVvePzmKES04TWmXT6xzfafy1hXAuHRgT5no/htahars3WYAYw5m
0t1LRW5pyOrkuGUavX0WDYrgXLXlRVB2ubgJxNpGxjNjcI5Mb+ed663HU7f/
VtAJzLVqaliO1dou+s07tWLXJ2ivOjdNRY3/ZSCYw0Gvylr+UtSnlWrlMRqg
qyUeJLCqaI0qjPSKLr02uvgLjtCjIAeXkpEXqLd6Qh9zdK4FaEAnQzCq6d03
hg2sFQBcB33lnH5M7AxtdFNtZewk5NJK5dmbS3DjZScyOii+dcsJQ1txQ3fF
MmUKtHUh4Xy7eG4Aq11TxygjKNqOeG378F+vLlpVSnz35dBYb82f6Qk48GuI
/0qCUpahuy3gXwaNdhGItaxo8VDyWrp3bMD23YQtDY3AIeg5HG6ouch1pAif
Hxq2xheguVoRj5eWh1amFANmWr6RY0F3zzo0O8m7e6LrZghxrEGSsxtBUrdS
DYw3Uj4BlBTGE364ZaSkNtqGqNZTAseKvw7MDWKVhAhFtYAhPicdRh5RlS9X
M/rZkcOdC8HcIfwDzqZRrryX1mzJH+wF59Am8v1a5D62+NQ06WXp6mCwFiw7
L0KiNcX/iG+F6SKMt/lgt+BZHdwUDho71ufzDQQ5CkR1T1bQ+O8yZkIbb3tr
eVhLYsc0lD3eHxuT0ecFPc8yigDu979ShmdbmXeov7C7SrlKgRN0y0gGgWpG
I+brNlg3Pu9nPnVjlHbThMipqtFIkZqqbG5rGQincz/rQHMMVFesxHSfVy0a
N5yJGd2GPnzEWTmF/YSR8fE/RuwVpbFBOTMxBAzQ1qUnTRTjg21q6fu+zNpe
uyL/J2G0CCbTQJMKXujidOerKu7cCjE5tAy8dZS09enAHAuhKUmb5frqM5mK
dHn7DUp5YL1BJq7BBsF4DBgPQt/KvfR8/GTrYxgymDe3VwIh5vg3Q95mo/po
HwejBcUb5JUtACXt633J1ejMEiArPfyIqtaUk4DL7FPh7D7SVVhRPC2JXgTt
SDmhsZuHp4aOPONpW3a3eeMDGMEowhs/TtFSqUdg1v8OWcVi9s1EFOhDrEQ8
xNx3yU8waDdxQ6cTdDYtONq7bDY6bfrl32acwIv5pf9mpPGQEqGyT337o5J0
kamKzkvJYLc0dhaiVrWRXA25EQfLjz4pidxIx3CHeXEXclnZYsfxRNt81IS9
5DmoKFeJagdrC2IidoVQVoBFbeYnuXX1yYu8N4r82bFnfwSXQLFuJvJciGX/
f1ciQ4pk6WHDLT3pbBUK+wiTaWCb+vmImJlxG2mefBt1pVf2cMxek97nSanO
Ho9N9y5T/mKF4yqjADrxAUczaSlsp9qrz/c49C6utNwHvhwqp0U9CvQFe022
z7ufTG2/QdezrrJwlcwzJf3dr+jDWpfxh3duVkNvIsmrUaAZKQaW8fCSqd6+
3Q93AekdYI9liII1Cnb4AiY9LwqBz/9ZX+HwvJY7IPTDmZYlotcr/mjkc49m
LJvNRe/avt1+7p0+03LfusOC5DbCAaA01uRWB6o41GvhsTLH7+0w5WPotQoQ
lZ8NDhVLeBBtgRjdJ8/6OcwX7gT8Bzwi//EkzT42rJzDA/wDTB3GVqzSHtgA
jGELo1lYFLMW86wVgvdZ4Zwk5fchfA3jjE/02YZbd4NoLAqPPfpc+95hoPUH
f/a6w0qWkfUODvsISYckZkUKdjQSPVTeJfpZi/vX8+z+Qw4P7Hlb6czuvgWk
Sa6OcQBiRhamen16ImnnM7S4UteFAwLWHDVA28Sk3qp08DuolPnFbOlozDme
EfMsBttCV1L8xBOzcSJ9oYpenD9jVdhv2aEk4IzNMuDv8DZcbgQbimEHGPvd
SvQJS/Oi+CtQis4qgUwX+vooydKId/g0RSE2oGdf5sLCqHiNouTmsqmoocAp
QrV5+enw+vSLDZLRriqdwCX1A0lVSeQ9p7JwZCZ/FUlnm2pkZ3+pSKcSUXoD
0QibEjQ+5KW/tUrBrkNquwDUn6b+Ha+hUx/JTWLdRF/G7+TH+nc8/QobJ+1j
KE1aiaeBTq0PHfDk3FfNseL365M64+9bEVwR0V8p/gzK5hP5Ut1StxMLBbbK
pFzhddWDNUWmIZyEeQOVFyuL9ejqhH1g2IYqYsVyKe4Ht92o21XTnC2v1QYu
alPV3u7yi75Xgx+syNjOU06+yek/iaxami4ZulOvzo9tMP4bPGFB6qSlXLzK
xDEZGQS2rN3qhB8cLb4Q142TX1qFWa+rzMExMyK6ZnxxAJx+Z0yxPZjoKmOX
8PlvHs54b+vtf84lrg550HTOPHy7xLRUN4YcSm5hrYQ32CzFaEDjh7axdUwb
2WPoWvHW8xreIlHXpCC6vZCn+cK8d3mtlmSP1lD5OWmEM44jYUoyuEThZven
LF+rCK0Y9E3L6I7EGbBinjw248NzOTy+Kwj37YM8Cv640EyOP/xmBqSSnhCX
UZNqz8Uc9S7nMiDvLtCWlDGMiK6Zn/6rCVSU1OsV5ZwrKz1S3hOVE7qFg7TH
pFlxH1O9PpNUcgcieZ7Dv0HsDAXenQGbfVgfonJBQtfB0suIvERBSrxinhy4
HomjauyH94MHbxtY+3q3dDa0gGE36YeYW0o5m89n+KbjqBy7OlrvNorCuNKY
M7BA1siazhg+UaYoV20CWWGA3kgsBSEU0Dzlxp3YjMiAOZztiefywEq8IWan
8OGYuB7bbmbzty6VhZkawjK3mGINDjc1gOZfAxkSIY6jX+DCNUg98vA8++Hm
Wt24wnqgyWixCFrZxGivugDt3tNoP6RWMXTYnjtdoCqLIPAKeQ0ntrcHnX2W
ytdEVFQn35H8PP06+aYUuvMshBOhE/uFRoNfQcSlZh7gAyhPkbUoLgQgg2E7
SdeV/BhTxtzhHmEyDz5t5Ys/lXEuGNU7982VJOQidhjPrs3QcLegnjobSTop
HhDY0vrk2UOPpyCho7ZZJnKqkiixN3CH5SJv7i3s3nFN5AO0HFkc7cQ2Fj7x
3U7RF0ePLUWJ48UYHEXHs28AoGHNv8evT9cHuF0Q0l+OFZM1Z6MQ4IqpZd/L
ip+9PtQ/RZ65y2tX/WsTZUqDmYesKVh12R0Evl1vkP1VCVJjhvoddbdEDoCh
dDTu/RCMWxwY6VNYR2UCANCBvb9cb3jk4JzjXP1PN1stThzNZOqyBa7sA75y
dhHCWLQoEh1uL+vunWBjvGi/VlJggprRsRrL+TzbkHfhVDlaFEBMwEK46AD7
eOMY6zmTNNMVNWuHgsMjRpbaKSsniUuXeSH0pluNVBLgYOKdrhdea+wrGA3H
OI17+lrXj7TbjUvcj65p1C6Ksgil/LvKAgIUK0GoH3gPjQFjSfKucySujVka
xbnnjr9tI9Wu+RuyXBwmaV77GUTCAUVSaShB8W8zz137F6cBPpX3o/GrXAym
OBoq5l1ZoA/YYft51zgLlirRUNwZXrc4Qf0dw3kRyMdvjF85hfeDt9t3ya22
qBn7oqaHk1IqejerVeNB625m2P5JNB7BsHcfLeDzm+l5dVEAYjUv/3TaO8mB
25RB3q3J6T0ovhTzq32rbYetHiiyl/a9X+Oq3RCnRoCYPUreEEeMXWDWAyux
ctBIr8OB+tBlNXdWU5bnatKiQFf8HvQya9Gbm4EENZxjmZ6f2SC7kr4zzkD3
QGNxaRNPTaasLa7pfxkROVVnQORdfyFp3a3ED8KmmzlU3VFp6Wi1vbnKgIfL
59Rez4K1DEBigDEXhW/1zLWy1KF+jwMpC3TLcoJFhXKp50txMzv1/zgjOhFX
N71HK9AjVLnqre5h+uC+h7oHbclHb6GJWFeAes36bmEc8nJ6x+Y+GnIONUN1
s2J/nsWZoRDOu3umMbWerQ76vT2boDA+kMICH6qVQnvkJxo9teBN88n1mwyP
YyEoxW/9Nrfx91r4/tEToy13E1Fyvpk9hNFLzSDPCQ2kNoBpheJpe7uoaaKk
iah638qmfzCkAl6DTMxIMuIr20IvmzyhSJUo/tzPUjx/0BuPmJBjxhAF212c
9NAD1mrArteUdg12jZt1e21sIpcYfrdeGdg+y1bBaWErIZeVGCW9eBk7fAII
ZdTGEHJO/0/75V+WhJWmV33NT7WOYwwPCSO4In6rMaMLYjuO2ZLFwVfqHmj0
cGWM1r9har/PMfRvNcXBHLweDmpuZ4SdBJwni17cslgZMUpBRZR2e/nRiMrs
6N5hQbEufsALU2QG4ynIbx+z1IatsAfMSjgKLFbSyABDNAVI6oqFJ4giRy8F
leC1o+jCbyx7jfK69n/p6xaKiBsp8eyeFpu4YbcnTI8UN+eugr379Od+zuDz
iuII6ujp4MVmAxYWyg1S+4YoQ8prUKLi7lv4MueQeMf7An8SW2Bnm+bhF/gg
129hhb7J0GtoyGfHcFOLT9roPaGvXksi8Clc3M5r74o043KwWYtpOfTd4rIx
IZQdvVQBueJEbRdn4xk0mcOQp6+dEI6HImZUhfCsXcHK1xugtyc7aBwTAigH
jZIXZOIBzQLHEMh8CRIDMy4tH/jCuCftwD3eRNU+Hkx9d3jASSLLtSVjvKtO
DlWRCLB+y1jt6uB45sDQtuAIehQYDWZD/7+oSSlCOPh0e8rvmSR4UWfgpBM3
Pe7G4x5GvnA8tpGATSV6gMKitqOQIJNZndqh5KCexVa1PuEietf4jRTCmzUW
dp4vMPObJ5XTu0hUjilnfk98j5yAqoEyaHHp5sbMMx1+XBYZhQ2rGPyE9nzh
DrG7MOdlrz9a/wtKhcxlXEhCX3BzfwfZrqMncdtwNJ/Kd3QSq3uTtfVaRGj/
YTx8h4FBrYY3A2xkp8kTTHQXi2FqQ4Lmmup4ozFfItOJX/D3G0n+vRY5pJj+
dg+iqT8LKejtykq2vOJL1TjdPqsaglMVdN2wIV+mfSjNxwpKy6o8vMwn5+TI
itrm0p3NhodqaXbv4hD1oeGKmRt7yG3NCc/KOSf9uQhSBhrgmNo6CfoSRN3p
i/W3beRHLaRecXp5mu7B1E+ZPqdkAlRrUpzQQjRwBDATKPBnmyaYRbKQAyac
hyJW68IKaBdmX3cfZ9YHjPZtNQ62CWAoeTydLy+GXJhFabgLsKG32npMXQiD
2CrRi99exZ6ArKOdG1z3yYF0Jf041qYP/1Qe78dYeJZ+WIm9s6GzlNBuaewz
Optm/uvmIo/7Zur7X9lT1HPZJMQonYzx8+dW7IE0+/uhKXWgZxtPA2+qHeq8
4KzvRa6ZiAfvH1XverT1SEAGgvDo6iEAyGTfDNhBYupusPbu4d7fMs2+keWY
Eb0Z8rv8CqFMzlWbRr7cduScXp5lHnPMxAXVjGgq7Z5jNhpbV6sP6LOEeQAX
Bg39u4dwlwYut9ggoX44kQ1Zssz/iXCoJiZlXfFg7nIdjOkczoZ9UrDqUQYn
zLPc9LpjhpghIy830EBvxwlUaUdD3bTd0GoV88twU4t5OgJx3R4Z9L2Rubji
l9Yv9DB5nbNgqPCkogPKcWENYdVs2gftYsp4JsFZl5UetTeXYzF/4TtCkVL2
K38Ewph2K9wujsUnLfbf0zUECU4nmSwS0Vq/xrrg40bHQ/XxDfFl0JQ+6vOy
dTDWbzJzCaT46K+Cv2jfm8xenCOSB+cvEA3QwcSwYe6CN1XHBF2kclsIBwRr
zyOppCv11WHz23jIRUeu8e1gNkZGKq9xaEboxyfd2PbM3TkI0T+FF3DiVCxC
WP7Vaaj/y9zb8SnfHt7eeTpfrcQv4IYQhMsu9DI=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "tU6WtkcxFJ0jFmLCJ7jDUCiC2A/5Rm5vWQSKz2zOUauWhLEyzXxKzTI0LaoSralhk2tD1j7QPW6zmJ6FZfKQzhgm7Tat0M1tCURYe6BQcX8R0O+oEBw3DzloynXgFPXHEx5tkfHDg27HGbgR+EEs2JVtJMu0aU14QI2OFZnO8p9xZ4CQ7dCvVWjKQjFOkpAqIWDTvYqEB1RpNTcqnva5ry8QiM3VVvAC3dtx4/aDkG0eIByQ+jDukOHv3/RthYmdgWT/0apnmoJt+BcWmkCYBZCf9P1jZzP+V4MuBdwx2XzS46qEoDXrIJSGkVfSg/VntBmf44ohCKejuhcSyaRUTNmDL7ZjL33s2ATSYYWI05vERPQ2KVfEOHDMDzF1xFThx1yBgKIA956RG1ouR+f8ftrVC/jIhPp0lVDBUJ1N0vkXi865zVkkUxrnLk1zbYGOqLlWi4yvN2QijOvD36H4KakuTVNyo7QwtceT6/8MiTT8CUjnjUr1cCwIXzEA5+m8saFMWwGO21qIl+lSOTz6gVld8tPYhRWh2PNhQYuYCO8y5ZXTYx4Bj8TecZPD7pw8fyf8JrO8ByFVcaNnucKJ0BVgKlHW9a6eqBVt9o1X/4IeI2Om+UzQ3sfgvTxugQBxx1wzHDriFfbh2Eg23emyDvPt1sfhHjJDsplW4qe4XNDIQt1yE4jpkKJNkVzWixetJjDTcD1jhYJWFKb9OUzqYZanK+9UGg1WEqvVqqYchqKOJZHWFiFnVl7tTRTJjMigKxJ1YWMOm4ncVhv/X36hvTs5/Aqz+sE9qk8MPFQV+jSBfoVp7M9xVnPANQB1al+lzjhEYwEwOc55j0phtUdl8Z+7UxTZ3GwYzKldbuVkCs2kuAj7jrnkZ7CNvTem7HXuijqk9LyssX4Jc4k2n8OejYUGVD7GFGba3NWR18ZbTF1rDL63qy4RWexylzzCu2Qa2ROhlnWXSCt6sfCRJ3bK6R1yVkIgnd3Nv+Yeu4Ks/hx2hq/GYyJxk/aMnGXQSoQl"
`endif