// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
q6LgwiFQqFtGkkmbYcbcBWZRS2848qm7UyL+8juq2nF0wGmawsEJymgH/h9+
1H006tin92mBobJ8sqAy1VBkm9P4qcFXtgRxIXENB6yjkBxjH8jcg8dj6oQj
4lQ0IXWd2qGL5r6UNlSOInTy2L/1eb/Hfi47bHZQuiJUYe70KoNlCNdimS7M
sRcKiXdQryPyx3AiOlZTE38sdBaRXWAm0dVNc8jx1Pej7gAWTlSh4fFeAJCY
utMHGkeHYoWFW0Sn/75qFGunqJF3hId5t6H30Uj2BwF7w1NQnVERAH2J2uF8
lhfQK1m7a/+vi3BD06X7rpf7YpODDoLGCEZT1YiRnw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
OlMGPm0udO8GU0n/adb8TpUfMpRo7PsLbG5J0OYOkaiVUcHSYna8FBHQkq9o
MsHvkoPS0UtyE/WQCxxzbtMMLJbSAw4gOYy5kNYUTMKIadPOgsOBTTQFC3X0
bJRgmPJlPp1bOv0Je3yaUZ6ZC0hib8/xTY8Txfdpc7BqRa1JHTp2T/eTQLZQ
G89nRrFUyhjj/rbquoAjJ8Peq9dzkENdUCGHByOGIrFLvEfiNSZIarr5FBH5
ZvKnFYJUYj45b+/YuSoyOnq34tjV83b2g6xmvMFVWWYZgxnSjaXDZHl1ksKW
0uBlq6y8FEgNxNhefSSF3pQuTYeBo3h2Mhg+FLG0rg==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
R0ToB6VeMQYMZJ+RkPHn4ClrOqfOwumqqK3bnrSVAi7tuLYKpqK08JvZh/yq
v43M1e+piAGxHUpD3n2uF5ye5vp3kZceAEap2d60dXXS3Evg7hAmOaE+cgxQ
BYuad/8sU7gofQSytrZXHxNDxoCB2jff4DuOTs3qP/0fHuMU3k/JdckN18ds
DbaJ+wNMCCpxgHabPuwW52zqlgHXD3rD65f1zltFHPOEUly5e1ivzBWb5IYp
txZzmE2WRmDx0GN9BvHQ5v/2xS6jRO5VwdhIgNBcHB8M6K5aGxY08ULM4/pb
jiId5dU7mveRIqMrgw+m78w3yNyM143Yz9AcZ5Pvyw==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
skSQ9nQ+T44UIfKyDPZg7hWL2MyiZdgKIxbVeqWkjJ0WHQdSGMg6cZ/qh7kA
Jgq/7E8ycPmCA4aPSeKhf5SIXjUjt8IYPhpKbiIucSL9MIuRi+eli6AeRtUk
HCsfGbO8MMIKqLa/OnP8gDAB7lVDAFsP50SSSpe3bflHElIyXFI=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
cZXDZw/WQ3SoPAG9MXCdFG4XbDQQlvMtdDmX0S5KjTYJAnDC7kBVDIxdUdpw
xRq3Y9fIiTcak3BxhzfemDYNktS1SfQvWh+BJeKKNL1AF9amH+8C0kmtprzq
NqOisnuDYBoMw2518BeYWXOCEsp0Z5AQMTj7KFno8wP7Sopw/52nLsMzqljm
TpZBfKr8FG0KDiYm2l2yamPfLgCiiYqlgeO/Ycpe1ZadEOpeQXxcFCqYsAyg
/8w6OEslrxYDcdhzdhGTnXHn8f/slIPctwNqsH6UXwE15j0zCzwY2xU2TMM3
LtOgkrtbSqa6Okh54rmnyyhINThUaGr+d+W2fK2ZB7aeTSlriSc7VeoHoj3U
weKvGYIrnYl3yOnc3nbsRpCdIjZwo6/fwTCO01JfN+7rrf413vI2U88A/5HP
3Od7RkeR7ouSeRVBwjcl2OH02mjy1PuOZlfyHdP3X0dkUTnXayeh9yhLOJXj
bVmpIEqVspa+e6WPtCV4cp/EQ8Boan27


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oCiKK8FNe4EKSeTyQl5h5yj50rrSx0VImmPh2fPjnNGY0aw5dGZvribT3m2+
0SOS6O7wTKK4TVfJp55ZvRFoDrhmlCK4JLXoHI2mw1gSKQDf++77j30xQuRh
XRSp/7kzj8eWLzBrIJIQYGaXS6OF6gY0ZMMM3k1uGNXt8+zxaOI=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
L+kHy44fJD4F8Pec/D9h1Q1CpRSNIf5CqwTd6opIGRUI6WD6PbxaXeiI3UXw
sYhugKSWk5/0oFYOTSm2l6uQi8PguzB4/nff1yAsx/M8N/+XbL3+gb2HRpGk
ffJc7hpn6S7nBGxnARV0pXTLMsh7iXAi+mLbSmSckho6qe7hcUM=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 4880)
`pragma protect data_block
K82XLPbqLF0yDxqLYSW0PtlsvqiVmXH75BBxj0ftWUUhKFMN13nMsnyxpYGE
6cggzO3ppm2+tWtVP0xpGGdbiJFBa/xL/8bjY0Fb+ifxMdRDkRFiLLO5w2Iw
vReUSU1foQCwC6SU4tTDrRVMR2RaPdK4me4uan4SWGhxL/E3Ic9bhvZ1/ARK
n1par1dcMZ8L55bEGwlT14rc7ngA5f8TWOHcJxow3wsBdqd9LjNc8I4p+PaQ
rtHGDsdwn9Oyv1jSe6XbPpub5DKTBajzPCMXShxcKUKacb1op/qWw7zqSuiL
btalTG092k7v8V5+TchjIwzbiC8E0bFylIBq4aqk0AhndNfgAKOchjYIs0O9
42LHo9A135Wib0bZxJAZHtsNuBf1p80LrvDbJtqrm9PXBTprxt2o8CIn/WxX
arISvFnWOhE916c7mQo8OjyVVDYNx+AmW2Q8VGAcrl+CxnUh1Zv6snugyR+W
4LewOvxdS/MPkQdaI/lSpmzokLGdepY3wUISvgBHKOfw70jrPWgUHDK+V7N5
GjLoAbAeXWpYeDMEsBNtjm2Kwkjgop/UbJvzqwwxjLHakRWjS8ELgukP/ZdX
sh75E7dL5h6xcpsnDB9qnz9yYPiUA0xcdzUcq5rlSM7MzVInGvp86ZhTT3PT
7HoIYuGwcZqBAJfjhq1Re3Od56kifAJx2sUVuEab61l4xnoxbyGrZSk/rif0
SrSmxSiwneM85/strvZ2+HoAw+SaPlPjSWzCWmn6k54TZLvTu3FdCe/JPMtU
3WxCEBMYZfMSWTazw2L9WfaHWzbZe3OyzCxDSLf0E6K1A9k2AGYzzLOZpipD
47YbWzxvlFf2cFv4/bhx1+ceR6ZL/6IqkPTyGhAmc08zoCg3QpgEQzoCvfpy
yEkigUV4YkNHjU6xyUZa8nQfFy139eGGc4kavaeAnrvT9f4qwr+Mwh46ReC2
qGpCjw6cOogV5OtCP3rEmbyrYfmEAa1ZoJx6mWHgsdIbiF+EGRJeiQlx97Ki
bhDOiM6ifAPIzligc6wBOGeAyQ/y4j2cY+YytmAP0n07W5z8Fm3+IOmjErPz
rx/VWL0Ubv7TzPEmowfTwrKUxSdCZZEq/CyV86g/KG0acAHbqzQsahSabPBu
I53uyJkbPkdJZGtOVb4OkqvSYGqDZ2fTOCvtax0C0igln7xWr5zGqpF7pfSn
7PATH8U/UrSUrSwpxFRYtSH/8uE4zE4wOkKo3e1rDWRDJL/Ld4SK+YpnbZ1D
jLX1LvbfGI1R/VpglHerg6r5UtIsuxpeddCLQwwGChNbyYuR7fh63YZZlFrF
+FC9CDDM0gc4jZcJaHpFCkSCcRfnZCaDg37dNGU0eIkLoHTxZyy3Z6Qy4kzv
OcK8eOZ0MVkt9K73q1FPidFXnYjUAVV4cTrmcN9HZNTySdsimRP95BzL8sqC
NVgK7Q0babkmpZ9mWhHHmObgF50hq74PyhTx92RLy3RnJdOtTpffbULg7TGE
4xOxTBOxk8B8D8dzDZ1gDwm9mhPpe+RI9xbA5L6UoErsKGhAoOl4EPSLwsOK
WFCx24J9YsH/19+22L/pbzmhBjdzZEUieXPlApnHQ++fpBVjFDp0IRlpG3ea
kbxEdXC9hSKxMlfE57QYALsgaLAc9qXcwP7SHYPJewt1tRKrMgnMQpP0e4Qh
XnE5kUt24iDHuJYeGvG9fWrdp/jSgglk9lHNcM3grBSF9bj9HWiOGGetZzdO
ZKXIGh6bMbWbxFiiMuLG3XCcTJLSvkTg2XP98itIbGMK8i1vNU+Prz7mMk3Q
L3Sfao8tx3587+GGxRUhPjYIezHzSrYL9a1+rPRxNulENwB0qM8xYPMtGDam
jOfMmfKT48MmbRBt3dVs04RbPbdjsjkvZ3di1uBD/bAy/NSrcJo9z1Ww9oYQ
0skP+eEyk3oBVws4UZCc+jmyFqSfr7RlbCGxhFXLckgIosdxMIEqSxaOPa/1
SaJmX4gMppEYBUjI4oMma2ZkfB+bKGedxo4ePsOAXLXfASPsfKLPlzqGrmNL
TCB3xYmIK7Gu4YZ6KaI4riSgDijw7RKCStaIPRXJEgYu1vLfOMQkQj1DWlus
Hh7gMrh/Eq/bTV7nmzGGP2k7K8nB/nbXCmViG5r3AXlPmzSvW9JuzV9tP/yL
ejxAOsUj1mJ/RhnD3UQeI59XfQdj4xqs6nvDUUWa6BNMOSH2ukWuGu6qS+ar
GPqZCBaaVvwORdxv/yOm6c4+xyX4z6F1tSNi16F9IXaEyx8jQRjZAFR5B6cq
yE5XyV9odLpYnjGUXudU5a1ipzbTiz83Y1EjVX/JBdZqDZmW206cq2ZdPJew
jva/I5j2ul0OLzacvE7XGXlFhTYw1kQYTXd0YWWQiFwlGI2O61pUDZmZFqmD
XZDar0QJconxGkwrRO7QKxEOxxDebWOdd9yv01tWzAc8WLjQ6uAPWrpX56JX
h7Rau4m70oqKNuZAo0QB0hfNAiPNFakBt+b2lRKXh1eTOK5hJjenHH5/3D7i
uMoX+GyZOppKA1PcJNw9INSpn28h1EFh2hqYojWZ6ma46n11c849TgxWWNn2
ZJ5FmEaE9JCNwiKpiXbChFm9N96hqBBGAPD4/Vx8PxY4BhvR4aoMNUfChiUG
SdsP2rol+r1TtCIYCu9hjChea2/69zhFoKN5MNzx18/ZIXayf2gzYsKt8QU0
1tLv2fvqd9rRArK1LYUz6un1S0AwI7c5b7BG6zmHvI/8o54NomUTxM+Javlu
njHdwu1BhgpJo0keLWvL5JmsX/bQ6WiFG8Jsm2MuLZBeQ8eHOdE96YingCml
IpI8yCVWy+rE/Bm6Ie+WYW83Ncpt1BNjJf1cTLttAAQ8PzDKPnuSjs/UT80Y
mM98CtWMHCXmg5vaG+F5wUYzUG55w6+jnFY/eKfD5NZb/DUWuoI+oI1hJ0Mq
+L0sBUCTSW/T9kjJnNesTQcUaAxY6RmCg+2cgRoJ4/vQeQkfej7q9djiVrqO
wAFMGT4ZLU9n2ZeCik+hGcQiHr2JEXpZLKYEyo7NjvaaXkK7TUAqBdLeQybQ
rZTYtb9c6iN9nn/KxLb/2Cj4db8rpixHiNSYvmN9o4n+OzgRwIRX+Iz89O3v
LZNXcdaW9EL4iwEJRVYv3dvNps02P2/Yl0gjk7M8Gu1tBvVpwU1YEY28nqxG
R97C9J3DUtFmrJpLGBQhs0k8X+3+FdzSAoZtRfOWaRYKLMoALlnJ/eCcGHip
4i8Imu3TX/qG+brEjhkBNwBSf+hhqnoK6gC8k5BLaxavJkyZRTj7+66n9oHE
/XjJcKutKE8Gb9Cd01+ZYx3CObGT3IpLZnR3pVURd1vVNbHQdCicoR00mZOq
Uh6i8IDwzeI4xGUDiGgz+b3mK/oz/qGrz3DEjTktPr+q8J5GizQ0LZdMhfXL
D3/aVrD1AGf8EqXmXQA2JRsDxU0KAj367dwnd2TH+jU3cfSc7NQvdqzvti1X
r8GrDComjLzevibuSoZ/L6W6yCYJbbww3Ndj0bZqj6BCT7YCU9w4lWviPJ3Q
fgbBZY4BZ314W4g+N//oI4KUsehTdE6Mh3+ZcaO1HLUQNiHzIO8cS6oxM7cf
UaVdQOqJNXQVXLiqJw21l5J5PmxsKMKwynrhZuyx8Qk21AiTys5LgjmxEgpj
emrK19eclQ8h/iAJLw4Gp1KhYG/h6EyTr53SECuUjx9kWQXMNnLknn+QGuRg
oQAIXWSpDZWO4YjZBpdHav+9a5iAcceaVt53MnE8rcc1M1aLdI/DStEbwIq5
i6wsdQFaqQv3E4jvjNIlh+QLqdQ6hA5cR0TDRBXtHarcXqeS8dDHawHdYVNR
wOHmKOJtb3A80tcmGeGy8IGkRx54/c8HwlzexeY5urH5mmRblVUGPNaBvYKU
sas8xMu8rXO4uauxhFvt/qhEozuybmYpyL6LTkumellP5xts/VN4RvPI86rM
ZuAc82NitVJynzFld/4hnmkpjwvH0Mx4IQNhsDluvJlTL9SULQeuC81c8bi9
TjjNJbRpy0wcUuY//DhKfwilUW1087+c2Y0QBiUmKxRnlUefumYT0SBsxi97
T08tL3drsE4UjHmXyAqfyibNDZFtsAMSyzMkOTOO/oCGKWMIcKTAVcCwH+GA
5myJTyX0nn2lAvTlc4zUmhgKb/SXU/f5JU8hhzucud1tEeVEVDbshlnLe5l8
jGKbCbGKxGnkivznynZx0m9MO+Ez1dM8ghgnoRkXumw1FQKZT2OScWNJnc4I
ap52EX3CcEs/gl94LP5dTGAtRfenHhNI9NmvGQCDFLztJuPcbD8bUCt+mczU
/BJRoy9yOmYg7oiJbmrsUeq8IjVNbyMxu2hG+I4ta3UEdEIQtu0Ls6O6M0B0
1qslhceq3ZiWYqj5hmXW6218HofZzKs1drHpx/umLk1EAwnfOpFUMttc05t8
8pEwODmguoReJ2dhHKq10qyVl1JeMDsugvJ2boLsSH274fCV+NaStj5EpimB
AiKjaoc0RBvKCvobrPoNhvWthNKktLlZHssN7xOZ0LW+gCCf/InA1/AjamRe
wqldNJHgXr845Sd+H53IgMAvNCe/KHvFrRw9tLOo8Wb5Je97LID2r5G2O8Ru
JXcG2SgG6trbY7Q8iUI5uoAUYZP4geLefNem6JxTSt0xEmwaohbvIV4EbkRv
sO+HzLtu4uMFE8T7WC/cqF2wBga8QAA14yJvxrPo2/QaMWy6aj3nhksOe0ie
GBXRiJtqdNCAwY3A46sDXudILnKSSWO4v0qCfGAMsqQXmDgEFEyMBe68J+9c
8HiOf8FXnskfuINSXRJzYlY6OiBIIDQbeKV5bnQdo8fUiF2RRbJS9Dy3CUkZ
LxA6EnJhW41ga+1xauRoLdheYCjhTVbk+H8OBzqVQR1CS/HV3FrUpxhWM0yD
MPvHHcR3SjWTuUsKkTDWGq9qoa4XUb0ju5ZsWYf04L560sYXd8kkrwiWFZiW
56GoDUiCJmZFN+p3n/cEvKx1AYHqG5AkjmxQaKP/3ql6Sl4DXcWulaqnTL1w
qvU9U2pGuYGP8HasAhAbk1dISYntfIUXclwWLRefXe3aWNgLjo+zVVO5m73F
SWovZJdEVlb6Wb2f76gzNx6QxRJC81ntSsN7cYEQf5DzoIluQNgA415IIX0J
EMt4QLtfQ9rBaVFGr8Xiiq4C3Fa4GdBtly2SfBI0Q5VSff7cBrO0JvwyQvU0
hBflMhxoPmZdXfTvu/m1lU3jnEBSDhDvaej7q6cU2Ey8CVH5k/d3n2uC6eN9
2w3aEBLu+SBIsQQ+Z14xrhPiee2pjFNnXugpZSvEmrqNjU+qdLXYhdhgmK8z
yYMGJEwDFdG05if8VwfP45A0X2f0d8MHq+6elObLbp9rbPiOUs5gMPA0UalG
gBXGMB8tX3l/bl2sLkIyySFWVMQ9yQo6ijlRzZpiZzG0aDzSe5qMF+xIWOsx
H89T0zzTwHa3Q5NYbNhuxOBbwX/UdgIzeC7yhuJ6n+ZuRGnj4Q0S+xrYlPX7
bRnbq69wvAtfWHLZ1j/cilfvrQ9rQdu79Do43IDpTfDGT7OW7Vj5yDA17EI+
NtBGq/WJE6HIF7XkVRGSzgXKLjac5imDE/mBYUShCYL023CMXcBJIAmADlG8
TlDmBmSH8ZzUObpZp5zhjVtSVQIcH5IFHQDdHBe0Y+5BZB82R2gmXJ/lM1Hu
lJwZYhqEbWzRu019H+S7VUAOW0ltQhDpl8MAzhHuSH5gtfWkV/aGzfFbV8lt
62ncK5PpTVTk61Wc3cTxe/cixewf49E5Om54O4+tYhDTX99QA69cfUTPJ19c
9le3g0QpJOE6Cnx90RKZpezNoMxryiomGirnr5oU7nCa2AXvg5z5SXWcFCmv
MpPngdTkKD/bit/HXTo3FRLPXkE2reMvSpg8S7G5B4usY3cISL59fELq1S7a
WxJGmB955HDu4azLttpQLCXGU1gFnioTMN/EEuIPIvMk3yhHH2StYLkGH0w4
QhRuLSA+67g8Gs8j6rOMGl4h+ILZKFZgs2tpeNOx9d03TXdG8YvRTF/xDj7W
wVlCgytsLhPpnjLkX+WLgjNO8GhmhRXmJTpoCXoQtdYTnnwqJ80TsYYQIf6h
KGGpcD2XT1NCKK9PkFc43rpt1dmexlQiEvHC/VOTZQx0X+Zon58zXB3Sxbix
Q5L3um3/L+jfbjJk0M7kGYvapqw/Yfja6yxG2YHOVIwhPQU1ZCHXHBoVn2VZ
Wi9q4MT+X05mxqAejO1alG8lr8qSlJEh9cVHogYAWtsOnDo0sbsm6ThI7ECg
FI7pSlVVJUAQhTfCqEfruNYYHXtGwt0g7TyufPWA6YJfRwECw9XTRWAZl5+U
8zzGGNzszeT7ZslKoVtBCpwzJsVIQF78+XI1NuptvSEqMsQ1cp3jGI+StVNW
Rmh29Fws6jPzHjcry01WZDRcq3GAsaTBbDy/epYMY8hwpztIukvXsDbJyf5B
m9xCF9jb6nBUTvqjLLmnTZgS1hU=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "2U0RSECmKr/g+vxBi599t0eHMkKGl/SrfFZGSXUORX7sahXbFFcqOyrkL1unUpfL4V71MOjtVklsNd4VGn2xgkzgZr5QcuaD/9jq4FudgF46VEXXZg78UNIfhV9uICVRrIQ9RMAotACOtaCDpWoAR2eQg8/iNZM27TK2CCZP4F++NAgTKU0adb3syE7DFFuaTUDVrZhYQe2GfF1jpj1qWSQBmI9iIRn+B7MolulYp3HZZgDHyx3OaRkHgBNT7ngIvaD1B7PH+ssP3eVnrBjvbP4iMWTp5Q/AFpZ/MUnui7toGJ1ZHytvgyUP5Ac3T9FGbhA168xGdDGxhmLU4EHvjwoHWjC/NFOazFh8jdrxRffPgjVJyCGPUUaWtEoeqzF5gZNG2qvg4PATSjD2pDhNlft954Kl/hXJlGKLf2mbRhk3qGiv6cepZ7zYjZ5+bxxqcmgxeRUXfeJj0lfJkR5G94roGlqswkNoiHOjBU+tCNpPCW6pc5bqnbJBbPDhwDmcUWEYLLIPDjtc0T9Ies0ETN2slqbv6mlCD8kVKp9IhEfqve9heE6n8xLlDPcPimhaP9+4Odmhl2VKvuttQQfODoYnpVj8c4MxeuHtDW3tpa1mxfTHiOWnH+utm3iUMZ9zFVgeG9fexJoKzI7LHj+pqiGrPl6iLE353ESx9CfmVAfr3Nkvq3y4NI6spUGAFdmqqhEu7j3GGwO341njWMiFMrtLecvYlJ8K3dPOv4k8YPgwgt/Hbn1Lsvs6hrdlXvonzBG3WjiHAp24AgocRKYS6TtF1pExzozA977bqwAVX3G5MlR/zH0vG4XOGYHbZNEO12BsytImbvA21+DAnLLKtdVyRxmyWodQcB5H/Gw9X79qtOmvgaa6cbnODWIu4XP2rjthon9SQZcIrhZSFTPUClzkm1abA7P/QXcODpCshEa3GJNLkWxS0PLhF+M+uJrTZTiBAaeWRbELN6Z5wy29n2sraNgnjM5vG8u/8I0mopASRyxKRQuiIubDDRzc5cgi"
`endif