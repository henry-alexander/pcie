// (C) 2001-2024 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
YkKswfx7WumyrzcUEvkbj82bpjxp9hi7qSrE7DLSm0QSQDXQMHRGs1WdpVlx
lHc3IdEFoZBtsYkTmUx7l3htL2Cv0PPmRqJDCG5sDAJzKEEzbCLa836SqyvU
jAJ7zUsfm1YvE+LHXMPWcBEg1yE3VxJ77Vnbt9C8SjRYZfSdfMfS4r7ujIrM
XPTrmoeMdihNN5XPmzULqxuV6FXB2FtC1QAK35z0RB7DSz34DMfOO+eU84/n
Zvz/BTHfNaNIKJYZO4Rd2jIeEKg/X94x4rw4PSmJ5oECs5O4VTfiwXCuj2C6
tJ7NsgLss08NcWgEIWQgF9i3CcskDZxQlzZrHj9KRg==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
WwoqPRlxZjavtNPY0TmDSMbcrOAWq6tI80mfuKDI9kq5CUFUagvFyT6nNu6j
RQKuwg6FNNdK/HcCSS8IaCbJVHxUFEi5unwIlp36VC/K6qOwp8G6Ry8fm1b3
DgbkIJ3cocv5SuMcEv9kQNuQK1605wemBKYqafmbS+N2seGbSUaj0iLJEYf9
7dC3y81IHozQEmWAEceufGInt2jFnxX/Ex49giH7Hz1hiBk/j/dwYhMunHwX
Det0Pk3TKzlK4n/a6zSARX7co5PYZiFn69EZhuMqXj9DtEJhhu8Nq1mh8RGK
AZvbAo6VybxPTGmUHco4jFzkZzDQBgDoivOby8IXdQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
AMtIL4O9xAjDoTkCMQDuSuEwoD4N0x/06gGUWBSrYsWNSdynzCIMMP+GgOlD
+ZdlraW73mdQMI3ZarTcLqm9+8jDQxZU7I3xXWhP41uSspAt2cN+YABXn68d
fD1yKqawpVX8u2BKrxWQmgNADaHcY26z5LKAKfmTaiNjeneD+sIt2GaLvtgG
SJqYYXYVw4/QVmSlgB3saHr5MJo/rgJlSPcR1qlIrOyFBXWSQ0lpfdLWHnfE
d9NaHjumjalFrcOIOFlZ06MiMCHT/uU5dcF/SQUbMd9W0LygtsmnL4Jn8J37
/N9iJrA84ZXmvwO0TC1c95ibYYGk4LzG7Wnz9IScVQ==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
pzgxG6C/8NCO/+jDKnm1DKte/SbEvTFxPPdz4LStcPiEq2Nw9Sjbjg3IGIGE
fTdmONGvVD6yXizfEo00B+sRk3UCf8NDllZksOKIV+QZOjpzzk7MS4ssLXy6
KIYXGnUeYyfj7CckGsq0ADiVcHK8Lz9u1wKNY8lcjfRgiPismgY=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
U3JGjlhVtIndkm0zyYD2e+uIT/GPw7KzDmjyApkKBgU8uo53VchasKRmjDhD
qtBtgRa7L5Xrz2XZavGG0wieQ7v8BiH/5xfyW6JANbZiTBQeSxhvIVLSSaHH
bMRpBkXPSLiz7n/oaBuG6oDy0YjM02wDhA/Z60mFIlqfjnPItQKwY9R3YUyh
8UbV3PwNDQiKPTAuZ22LPzuLmxrw7KeIcy8WpFHfiSlqPyemVNzWJXj2lqTX
8zbcdfgStoJeofmi3u9Yz1VKbAEf/gOUVb6klbGfdlkpWlC/brV5rVf6yumH
8YCAqHt/KG50YLmbW5SSm+fHMrF5cIhT71fYYa/XP2IuExS2Ng0pL/n10COL
I++cWeKKp+e0l+K9ShqTSfcNsLh33P2p9BTcDMH3JwrpQmUSsiwRX/hqBxaY
w+nS4qdxh/mXUaJQU3ublvtOLQRJ1suEFGyjiM7oVqcSoCdTxl5DePpJs7UM
RQpuHGyNlfuhvkA0Hy94ZW3EuJZzTC55


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
aGCKMiG3T/MGihJSgzRSSKgeBp9Pq65bjaKOfuwwOoSfZBddmF/PnBtNwJ6n
RNP/zc1u4GKJkzNwlLe8PjT83iJ2uF+e7xkVHj3mw8T64QH83uu6koZPxwbE
aJ+hmpMLqPbRDlZr/pKnrc1WkzUuyMk9YP8QeK/NSSEB/jieJvQ=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
jdyS+XQohywd+DQuipkz3fK92CtPUrcpbg8GIoezK4KLFXrOJVsPd0sSkudI
c6oyKBQ3Nhn6C+sTk9LKcHDLeHiebMu7oVcVhbzvR6htjXuVkOlMvE4kwjOz
rsk6/IOZ0OUwPTvPpPrHtARH3VhTtNf8SJD5lPUa51q255SLBV8=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 76928)
`pragma protect data_block
TwgS/d+khYRCLZyWIaEN72u51yHZpftEbuT8R5cVhRCkFKwGxK7FN+xfTLSo
NgQvQ4ImnwRiIxWCMmy6wRWm+IBZU2Ms2HI9aK3Wg9KYFCWT+ZYISV5WPbM9
YY6ZNjsvdOuiWG3NjLEAUs3lqLsD1agB293FGp914WjBBjEwBbWpENewdUxL
o24nTpWOxQFSTyxbr2b/vG0e/4Tb5FpwsxfHEH7MSzjoSzqiXaU2NmgV+qGR
bfzSEC7fgRWvxF19U2ujy8LxhjzznYUm3DLeQCy3CJEtF+VNpNgDE/mp9wP8
TfJCiZFJgBBKDriz0egY6cTutrmyordE4NzQTwKtrL4PpLBlXApjWjpeVaV5
aq4PDiP5XM2jlvWAgOhD61+/9jOKHuPGqV4Uus6E9oEypBHYHR5XFPUzi0GJ
5A+ifWM4MWGfPoRABdqSdpO7EuI7LXNL6HOeVMmEKBCdTgqMRhTJfg6T2lqp
IXUBKrhG/Rg9DvaUMwbEg/xYkCse3A0yyZuF2xmr5LX9vbaqM5Ws3pvAjI7D
/sWmB7YqmmmomzY9Q0zXwQGkCwijzpUNVHKfUxWd2m2ySS7Vdr+ldJ/qbmYN
zxxQZ3IHDch8hILFNEa2Gzozi8OnAPXur9LYJeAx4shbqjaAdxKDdczEXDK7
OnVPg+YTl0UC4+iBkD8DFRnEtO5+Vw6NmcJJSoR4Qxei70vRQ1S1mCz/hkos
uRsEWkhr3J6FPM3xmMNpESr0nyO61Ph8ri/TAX/61+UyX8LXS0Z8J6+TmjfD
xkXnICSzz5cFrLU0Q5hkxAIkq8J9sOzK8hhNfZRNxC9Sj9UJVkmEFOSpv1eY
ql6GBU1uf/Z0WK5P7h9uBrPgQf62yTlZdA4gfRM3UXdP2Co9OdpRAi2YaX9V
7rX0Zk67k0Wmmjg4oALd2JtLGIvczkeKLlEXVoYkjRkngzRGXoFqnAf6tPDe
ix5+mRUIp4dgcC6LESFeJNm4J+9uDbHvkGMNN0Exzm0RQKcHgsTbjrhwWNzr
gAmjwGspoJHkU8FVCgwvMQ80qCdICxwxtd4uXGDU54vuBjb0IK5Dydt0FBiW
/wPwaiFi9pM7PxOVDDdfwb8bnGiwW+POEhQbZ7i/GiB4cIFXTnPuh9tVXF11
uHEoSok4myExiZVp8ETDbBjRePX2gkeFl69z8/lQgzFBbXq8uKuuKtwXZHAr
Oj1Vi92zyjKx/ryZWPr4dr2H5Sce1tlMKIMpeH9DXusTg0AB3NpIOLproPwI
GkwgWdck7QHbN8h9LzRMGmXSozK3jbrl9cKzkYft/aEk9f9XetxWiDlb33aD
zipuxHWa2GeAr+NW8zq4GxIcsbxPlxKzp0nh3KcucqAGkj960gM8g+XDv+qC
BkHtLb9pRowuLYyoF4/zs+rFNuQ85+u/ulWDZe+bXDd4ZKP/2wi/ojtdKzxl
9AXGiS5C20NJ33T1EVIwiFF5T38VWoTU/PFn7ey8kEB67OEgzsyLUrBlq6jo
+jF/kCECEWO1qYXA3X4FDOMCWufe0D6jRo0PBOAVc2VTZZMFVqQMN7kcDr6G
e+CjZMi66NFQjb8kp9lMkzPdPZi8uY6q8wFlwaUgkIubaKcSEflDYEhg3l3x
n4k0i8XcOYipmvd9w2+Dy7VpGrdInX8hNra0tZRRnyIsKxBVAXrt2y6FEESA
TUmDRj5Pzy8vK5rLF+R6j1vrheSsuLFJHzaTTgamg9qhT2+Qkg7wpJumq0ug
NiOXOk0FQi+0VeAhL6OFtyXdDbOoJTZSFn5durQZnve0jm8S2fYZr/Uy1VQ5
jnv3A77Lbi7Gdh7CDEvenKCnhHWQRWX3U2IeIBUvksYVSGxBbq3rOoPCUWm0
OkOPrDh2gCFpH9XkcRXquu63IK/KbyUV2oROLAkW7BCLtt+N+72i5MZEzIna
GazOOAPoDQbuMQy/IyDJgcU6bySXyDUbMeY6cbcXkDFNsOumXihUSntOiwWr
kBfobwVC9M/EMUBaSKreOAfwQcmmj32P62MpAn+B3e+hHdTc4923NDh0O5nq
0rIEyobAWsD6V8mMK7LwyHUoROAGl7kupJMzQoKnW5m0J7tD8Av6aEIf78FK
ujFE6BVfCrRrXPDPDkTbykrxpC3eMJNA9oOexRRPx1PyW7c4V9pTnZE0+3vm
BVq82flYpGYOP8ioJxm6ZVLEudfXup68UBNrnkWOX87POuBn8a+MxAWBIKvo
SuzlZdDBbgFf7AShXk5co5kzWCYYvBZOLB138SmXaYztk7sVJTu+NWMx2tli
ToG2aCxUWAZz08oBsCUfmrFYc1PJ6rC1s9yZZ9By9Ub3ghcbnl19Ad2yJ3ug
0ftYqd9Wh6AqvkgrrC88z9GLN8CR6q/MeGjZP+zWeS3BRWkHRGhOtBTBdU+U
mk62ULjiJH6kLoHw9zGTweBOeATggbK0aw5VU85phXdN59DRlGNI5sQcB8e9
qpSFowRtBFPG2v6AV6VrxQcSWKljmZxHd4sQ595gIOFi31maZH88t2OyrYRP
bBtfaVdJqC9SUdI5YKzMk+AYOgRckXXIbV9VUHbbPcZNjW3GY0EL5hzxir0J
OvFyRJOwaBELbhvqw9o4fFRCCx3/og4HOT+QrpM/Dz6RgTSKlR95UQpFFwZI
C5bY2tkbC45iZmn0LWcmetl47rlvaunbjdDqre3P3zVbrumtQ7xEdYdrtMk5
BMcCVcHNwx1YpiOfiA6IpAVCslfDB5ptgmhdRLbzshCRb5Q1card70LHeO2i
vqpPqzBEWkegEiAp806raCkQT927FRlwmYZjYtmyiWp1xZFtn7sk2nIok6+3
qrTQmul5pr0Dp5isj0vchrnHLFgELqL/27dT+IQ6U1MsruMBeLcVwI+DKZ5W
IDBu7IqUyBdtWkahfEcRtdjh0GQOIlbRqi6lOyWDjEgf3mtKgOudYI+HN6qU
/MqAHb6RshCTBWa4N3rBYstteFuJfdzGSm8sJIXcqM8BXTS9RfvlUlaihB7L
8XrJBVLAefoCXcclJbLKMWWj4o49CHKOPnCgV9rTYOCJNBrVoqMs4Yic1mPw
xwrphPxCRqQdwvTG9iyB7ZTXlD8vD/vYvXfaUdnt59aqB/tQXiA5NpSof0jo
EQGuUKhvYHBkRxI2eLZsWD+f4InT1iNXn78r21vwB0H2f73YNSUWJrYZhEKM
cx98vmx59b7zculK+VWhMQtSH4pdGzwbiLFLyQbDeoczobv4NOyz2jllo0A5
YbRgRXDENxReTI7QKavMnQE7sIN1Az3iapLAYdzW54+wgUVvO7J9PSzBKdOi
ck/d54157dF1TiFGBfjFzPCDhN/9YMwRSZpfUWqgo65cYduO9oxKT4vXUNDB
rZR27XrNFMa13KYUjEWc9uynTc5U1U3QhtYnMKddPFk+/dtA4K37vkFR37VC
+QnFZU4J0MLA+phgiUF0fPueVNSRQPtSdL9i2ZgbNMmTYPCh38/9mKVcMDQX
8+xbzg16LqWaVupOBgiyMEZ4EpdpvjjyI3NUn78ye1/vNCpFlYtJIBvt6f8C
gBGi9L9csydLy4yMtCa88NK+ZL7M1x6sEEX/5EjXxiByVj2Pf/DYVWj7uJGO
xxZ4LIXe15UL1yn1p8a1XlES0X/UjHB6uRXBBEVcs5qviaCflkmFnBQe0duU
Xx1hyVDY8nKTR+IE1vvMhSib9WHQQjPKqGZscVIS2E0quphs4vWFpvBav+K+
aKu0rXSRK3SPTyQsD7Lne9gP+H+3F3K2OWRQX6g8E3g7FIgZwqUsLuIEUp0B
Shy/BrBZt1YYU8NA8bCidmxl2roBQLYW9i6Qj+P74CN1hfonXV0A7HNXpncT
gO7Fqe5zyB432BY6S3PKDSc9XDj73jE8bucwHffrNaeD5vgM2tEkh1tGBSrz
s2eM2PBpOH/ZKWvQYBnc4wc+bAJUGdh45z5x4glm3XQjLawIgyUJxQoKC2dv
GNcEod4hg26O4KzuwbEUCRChWveh+qC9S9D3zgfdvy+CumCVcM/j0P4LdZfu
7ZPJgJV/OR8235u0WODl5ET72rMUw+WcWTe4o+knv/d9/dWTfnsaBORMRKzl
7T6mqGCml/Qt+8QzmcOsPuHIsmZ6YE2VFVVbeZyxp03x2r2uusG5ikh/GtPM
F+lWY9a3ftbnwGg72qMm7sh06nhZndvQBkn4KFmAwjhaZlnpS68E1XjTXFDD
e9fRBiId861CMVvMjxrllru95XMPyftXqSbC9XX2ZTYrc1bDyjJ08lqnwbJH
+4DtATsMnL6SB7vXe7ap/wcZMDG56mRJI+KTs6DWCqbhmgxboBpEiGQgF71z
p+ikF8FDKZCRDtcZw98qkG0ZisSdjrbAryxniISNeQetgLCJBZX38uiOCOr6
y0sy/mb8NomXB71s/v31NljcpwpZptoJdLbRj5Mi6KE2+FiF/ISShgYHPUeT
vYTPVXgPVp19NzowZ7vmR3fYSGCGoI97TCZYnWs13UtpEEIGt12l+9zmyQRB
ZwveiLt3liyBwKzVLtIYi2c/WKn5BDzzyqhmveK095PZED/YbeW+1dbfdneW
hIq7MBLsmlH4EZnk+2xCQknVVOCL3kfrkVABJWOzMyfucqh+FPZnZ2QUo8h6
/2ByYUO++o9j3r3Uo+IjoFQqSovV6xLXxOMvNGN8jaLCOzvDDdTgYGMIVHVY
ga8PwM0Qv5EAhbKE933T4opWAcg/9Zdhf7lFRmtQ3iFoRlg5XaaEh8MN4NMd
0kF/VmBD2pWel4Cuu+8a9R8GTFcZCN/lekcg5TuNC1j/rStfXejhY8SR35nJ
GJtOl016Pnd+w5zu7tLXO71cA9ZW3GpkwR2UCovolvitg+ugRyK1qZiupJzY
E5UUglz7S0sERme8M47goDbiFemtOxO6kqSxmQmkMqm2LSr/mC2RleM/oS8S
NzreHRXuKQlkTFxVhFnHmQgwD5dEZ+UehLc9QKxHRFhufTWbYWNtX89+/CUL
Sv/nAWFkopUiesfp1S/GIpSgsfFzbXXJrA9ZkSEtbN+XmXVB5A/Jf0NS9MtD
bqOl4JcJXMpbsSbI5UOXkkwifUCLeVirIHzA80KBMB+8wCPxoPsWdlmHHzfc
OyHZJ/hnwUUrqNtvjinYMadx342hCMeSrTiX0VpwxwJFC8AeCZtxlM2Nuh5r
5qwIzZesoOiV3DJoVfIeG9ttSbDVGpPRrD4kR1F2jnqKVETB47F5a8fvDq1i
sYDC+60L9LC0dCqJu+lJG7VdCAmp0Fun3Ple5Q1kTS/krvhsID1qY9kPUpuF
paDEjK2zwX1TMn0tzux+xZtvScIBU9fu1RfnDi01Jko8+Y28SQII8tKsLQtu
HGYR+tDxrEtu4esBBJOHO0aymf5aKFg+Z8yM/i3OgAIdyuoLh+uaQVmsbFdw
xQBxfiufWjC1vCYAZNaCXXlI3tIfWJlFHPps68op9ydzMmpVL8TL1i8R0YWt
UFBc57CJv6VHoPkSbHgV/Wx0J8UjJH1qr3DorozXFmeGbnKaDkoPODBz6Mhx
F+DJQy3+VIR0qs0h509DFKRqTSODiVPCs24PyA7SYy5+BaUlehJV1v9PsqCq
1kNGdaomS5G4Js6+wJfuYMSRBXZtF9pJLq6iLi0wtHZ9cpoOqICCdLlmo/rQ
Fal7DNF7ZJd+7T+bUMfb1r3ebsfWlT++4dYHJuyl1XzhEkm454CbDkOOz5Ss
nWBPZsG6FG2B4pmt3Nc8JCRdfd2nkWS0ItS7uUu14zS9e5NKliOp3gRI++AK
sjRwcRlVf6zeUncCnQ9Kp4NnRkycx6fkBE9oHtYVG758i0r7H+5JcrTLFxb3
iwCOUod7sjzkQOv8pzjMX1mgN7PWLM/2rJBy4SnE33cGDvOIVXpFF0pEyc8k
drjRW3AuHvrJkNVMnb2AKI2F1DD1Wg1zkCR91PqtWOSKcoYf+i20o5ywhNIk
6WMZatn5h0E2X+j7ESFD0RfT5KZHn8B6Qzx/4EAt6NNm1iAOZxaAxheeRcxb
S/u8THi2w0FwypUJYB2Q4a0abXw1UVUk1aflWPgwBwIGTktT/2CLie746w1C
PMTeJA/L2/hz+vn1kGyzWRFa9WdqmNsg5orPHxPFqfFNqCO68NOoa12a/Gl3
fRBxnQQfZ3PQiseHg20WmgLlE+LUmUhsO+d22pjz70ufv3lNfAto+ffa3c29
TSM0UZtkUfjNUv1Lh8nNcAyFdGK3+HQWytDOBOTuCkRJ/pmdEJA3nt7NLdr+
IqeFFWKrktpWa69DcelpjrXLSCPat77lFBr5TdUzQA7wRnIsqEsaMGKK95q4
SYMrI5Dgi+HgFRfgUreM6op+byE4TnvONuBgLpZEiE1QBdy/7zRl6R8sj3IC
2Dncc+a83WY/E4En+ensatx1zWbivxBPj6paueLNJgNwq63Qbaz/UdezDqKv
V0Ux2Ji+xRRlCQzZPBxIcC3iH4Jq81Ok9yb33BswGM+vC/3o2q2qS+m6A1Gy
jm7UV8iJx2v1+PYuXqoPVPkWA7MOselOXEhCltn+Nn0LLHES4z9P/hQXF3/M
775EEAPMiiEo2cUr6sC9zBfLYDx/nUmg9LhhmH+XkVBp9cCGfdUMnpA8Be1k
NXq1YMvbHZy109QCnHAbLWyrNTaawJ3p6kZ5WnD6HW0j0q7VJ3T4oWFyV/JT
3lz8+qu0kgQfFGO+TuaeMIkJVjv6idPwpP9Zc8bknBAvqvGIwtOf+GBVNMNJ
eebml9d+fyPs2EklATj8Wt0oJTMeRP/ii73ZVg8Ejy/pWqXuiK3VFdkYICVB
coyqEuzQNq5wbeIwZuFqWbOl8SW2+DQ63+NrALMPu8z7FbxaYcmcgGvlpoaM
TD1L3+esr/7YOhiB+Kom0j9AxVJljk5WOTtW03T471SsPAe9jDGWqF+RSHdi
vlIdgI60UlvAS2lgzKKqpEWVHyoqgQ9A/rTpNe1EFxx/ZD76pqRC9xmWQ2nj
jF/m/CnYLKsRq1EnocdWTRyydAED1NIV3rVc+/0Zr7sQumJss5GrDqvb/hVs
VXBHzrut7KP3DGaOBSOkya/FeKT4vDU8O/imTCoa03hjCXSUS8AcugmJeXSU
CjKDPT02ObJ3Yboe4JvwVJQSGNtwzbhG6ePHyBzBywvpvmZ27Tlf//lCO759
8gL03vtI85GNtahrQ/3W7wE4fZK+rilGmnlH/V9t2mWpz5F4RWrNK+J7m+ah
xvSFnML7AAsiCVsmCclvGfjeLMEgewuCM2v+nZEx/xp+nUGSdMktAHmHQL9W
+wXdPIomKbvIGuqkpY7xA+dN6vhCfG+CHL4Y4jxzhEWIDnyKEMubMVK5JKGv
omSNh8c/rkwW1QJoo0ivTHM3azgkJ2cpnH+hlYdaJZRaOQjll+Z3FjGFmocI
J0QkTaCCmi+nKWbDdTj09ZRbG5CBJ564q2KDhKxvwlEW4wEqvQIAsfSAPJiN
2BG6DP/+LYb4d+Jg0ieaChsNSBQpatsk/SxbxWpinrhdgNP0GPtNgIMLlkwf
wjwT9WEOk8H9sJd7OGT1nFj3/3nPZMnrWzQkfVLx7ChFnbG3U0EaG3kaFrxs
ejNZFApenY4CQ48QS+GbDOn0GFVSzQCQmaQE9ZtHbcjmE7H05EO5gSO5m2aD
Y9rUJbU8imZF5qUbPGJxc40pRc0CQFJfuW25/6pWpcrXSau5alI1eXK3281t
8OMmGFBpw+6XT6/B3mdhsTy/PATufslKcZ61pXAx1yuf0rqNidCDANPyh9Uz
qkMWwyEsexQO48J1TTQGxtxvYTfx35A6hpfosWXFZjlJx+IVVYevjj8vGGG+
hRCxm8+qp8d4Sm18mcA4hh8J+XYU9Ril7ZkslfXO+2TosdTYpZOLv0zJAEFW
pQyg7yUwMU01DSB9wqO0Pqwbt4GMhYinltp9DREbQRjXFvGbyovgnct3Hptz
BrXaisfTY402dr5ZlevT5jERUqdS9EyESxMc+/DMtEYqEvqgOqTTkeiCnilP
tDVkyUkbN71WyeH59lVHnOqyK6ypDzmaYB/lAs//88KfSSxvr9B8gHwBtILl
EJge97LA4CTuwo2maULW+JNr5Y+Va2zPm40/d8zvMs1UUVSlhR8gGkQQJaW+
OrSNz7mnsnNO1T7IRQkQ0wh/1ovreUQcrM8oKno3Pli9qv8qPxBtEEwOu4XJ
ttrtZN3yIQYQbXvAm+A2pCzJedJA1y/G2eyAZnHevUggJosj852F2PzUgmV7
NO57fg8D6Jl5+6DTVEzlW7F6hOE50RuOzsO/mVhcTzDKjKc9Vo7ZN2NfN5Zg
AM5+J1Pxk5NEFTUJtt/lZlYEcQ6w7eEOiwkBHffkFeifBbtr8yorGuFgrO8o
XvBQzTQzeDPtyJl1Nu5ZQxgA4GHKo25S862Phyu0+hgN0GHAP37VNEJbLme+
1r2iv9Jhm6nA4zWM11xUV8eofMwuWsTOHy8PTFtRJUscOYrtzuH5ZawhVnLy
psIpkbOa06dptmo5bpaCNhAXCeiXB3E6i3sM5uC6jHz2aai2E/RFO4Zwig4L
8xi0PrfIYEyxwZjVnYbAFuwNNwhFnTmO0jvKyRwM5af29zqz0OziIuPjlxwT
5r79pEwmEoPBwkL+3S1ZwX4JlQne/tihvGfDz/lS1rBdDFp6TisQa7HR992f
3jASEviWnSUDYJ7ZZhpUd8XOfpV7+xzOjW3mGaJbraMUSrcvp6TnrCaE81b+
7fz4PwcbSVv5zCyZ5Gr+Tivfg24o3jOLk53G7m9yJM1PJmUXu9cP6ICzpukb
93VR+NiV/8W7KSgBzw0aPNKcyN7xa0173dq6+tgUAtmcyKJFPlmK8FX8xbOA
wWIwBT8OEVFUgKYL95DRf8WCxcUmb0cM0wdsjMy6vFo/PZPIDB/5H5Z4/lsW
SvD1ujXBA+3sTemjuE9yuZXOTs/wpunrXqOwM5nfT9pxJ+khRVMijdzy8/Ob
jYB1YBdjxAlGRyjiyP9eNXlgxw1YCas6H6x9X0CEHwo+IBsdJToRBLZ/HWE/
PmHn/JosuxCqqDnkswz4pzxZt8HFtFrJcI7527oXCU+nB5brMhqNtm1AvafA
QvHVYA8+qS+MHqDeGxG2yeZK6dy2THnV2pRpAyhjSK+MnGo9Hxfov1qB6kMX
5XyvaxAIJG0AdiQKmfUVhgAXeoF0HzPuRurt6VDDbdHg7m+BYQTQ7XDGzhCs
pj6VmKL+7S1OKUUjEZc50FFyO8zhB0gW9IiDQfoMb3Os/nok9mTwBt8h4HL0
XERzMPgeLyA0tvc81nHmwUCP/RsNbChwV6YD80IC/2lcPzRT5YLt+FrcIumq
BGuOaV0rgDNivTZolmuVRoUT9h1wVC5czwkV6w//St64wkcQfN1QdxQxr7Xu
FeQnoW64vYcD1fUbHJ7TK+jp/Bd91JdYHbjgHI+oRAo4COs7yIm8yXGgAYFY
33XjXLrIt2nauMnSRTm/HOkFXYg5e+tZ8m/Pjlcl+PMXlnAPyGrTBWOW+HmO
EUFGVEeLwDlkCZqzhzps5VOgpLaSgDC9a98XNL3+XZH4FN+RMHiw60R5i9LV
blC4yKt/GqziRqXHVu0Qqp3KcLHB4txgLDenVyG+mYaQCFJ7V4DVJBXXesmQ
1+FF3XpUtOukMT4Y5OT37ojHeai+pWF9UdE3mAzwMvgJOKfVOM7YdE7pq9j7
T8hHjTVrycAPM8fw+OJ60PyFCoH2N5ozLQjOOlQfiACffyR0PbYP6cSRR0/E
pAFh6nEY6ijUCYd5ZrrJ+NqXSKm90mAlOdvlTbopw5r5PZOqoNxoZpb3+537
u5WYUlZ+0sG7ebJK/lLGIp9S0AJvGgP+BB6KAkrgO//BuSNO8GAsjBcEZPQn
MuKs4buTb1ONxWq1Cnrms/Z2AmGcE5IxakjkFmljmAXyxjaQt/KoeL963Ugh
OeCMPFMDiT2OvBaiHyMVnTmVkBHkW2SoDZKvEZxxsWKPiMjARnebwwgMIydZ
XxUq6978JqxEVOFYUulBc4a0YJ+n569rnuP+7R1AXECvV42ZORY2oFj8T4pf
UcRqkob4rZf5nfJL7GrRGIs/JwtP9TK9VAvNDdazY6615L5LYgQdvb5uI9U2
CeGJFQRqpnUr09pD8zZTy1OZTBeFAChHq+hLXw6kg1IlZWJ+4/xTmMCJWh5m
mTS0tnPKnhJztsyFMRRLAOxRyCHlPFrdD8K6qfmMse8e0oz0wYwWNSqV/pu8
LfPZeNg7n/WV130eEheR7JZnBAC8gHvVSbmapLWRIlJLG6sQKJaW6OoMZlUg
UawgWWKzzAX3RYxg1WscKf03C/kaSErIIfwVUsybfeIEp8SouiofyUHma6m4
Sg5TG1gApYF3qbKQvxFgn+7M0Zcb8O+cGQ4t8zIuUO6t2J7XG4ILwI+L2N4X
DQQTy4wvy5vADxp9knjdfwW6TX6zjh9ASreDE6E36K5+BlNqH0j5B8otKffs
JVh/YXHi6V3WuVMT3bYb8CFY5/Q4TCs1Vkp3QJolblafTk8YKbR2tK+RFBNb
RPteoCMOO3naU218yiRGwpNzyUaSUO0bP7yyn4n0SfXb2EqykUf5w7IYi9kl
fcUd0hSW8f5LX9cBpm8dPhVnnWwXxu8KrO6UV75kh0Y3y3t0dNlVIIHCwu4i
U//UfihMSxuoFhF0xACZwjoleoFPMNb0gYH8258cLkYeENu1RqFVbXMQHApv
qj97vJhJDe4makX8blR2oOyrG/0yO5afT0++V7jo9Xqah92SLUOR31wYEXmQ
+eXW2K4fB2UTY83TVrF6rwRtC6iBtZPT41HaWik6Sk0lUgRHv7S9UP68wMMh
B8rYeZgzUrl88yt5GCfKWYtvnFi5ZFjUrGBf0otuhnvFJR3dNlv28MMWVMXf
5ELSjLwVSNDaWL5pRCE0r+d5eRJJGhwe+/v2YeZxtdBX5HF4nuH/JwwuF9Zj
5ZIE/7qP4AUZe7ElidnZrfyPQQhU9MmrJnkqsX2NhjyUxtbv33tIYhCHNavL
C9gxGiYVLlmJcQ/kZmJfpH/PaxbCZu6y+nCo00gcPxtpIytg1nNCbPbBsYuS
LxQJykOAJredakawAgLNnSLl7wMcajyYCo3ahBPzEiW9RZ4Ix8vS+Ih0gQWx
NT3bgTJwXQZe9PN3Q8numCwaA86V6A/LmSaEsXD2d/5Gp9bGI46v6LCMW5Y4
s/4+aqbDYNPjrtgZlDrLFas3HIQh7fs/dD+NR0Mlmq07qJg/Eoq6bELz9M0P
zbV2kSsNZgi2vGisFooi6iXhaGGUgE/YobYJb3+UDgxXfYMO9x3w/5APW2qq
JRYLMDXYlu8iS0sdejX6Tvf7y38ydGdZuXtV29GCAQvpDOgeoWY8YuOVAKAT
yL4hGllJavvi1d+RvhjYPUfwjiWi6NhKErcVICbv5fiDrgak0nUpAb71oeZ4
p7X/RD+L2Lma2M02sFotqzafKNtuXohX+1+365prJNSxxtJruwse3ozImGHL
UWpi0mEeILq1Wii2+RRURcnNPd3gMnWXf/XNPoAnYZU83/JnweylPTxoZSWo
2rxyK99AkJ8UMbZeIpCr3Df03DVwKf15r5SNw3lJVKkbgMgRuj/IcZ22PBdw
XcUuWP4Isqu2vjfVKFzWT8xPwkTB9lnS51uFB7JWsPGAqIK18wZCToy9Hz8B
QoR8UQcMYrpTyUbOts3fILrj6m+pzQ3j8Ohh7aqu16Y6Bm1muVuNn0NTWDXl
iN5pQU5RIliw3SFvmmgiSDl/AU3upkFwigMdcunGPImcYj6ooLojO+oDSKBi
+7sCkxWRTX2wjP62u3a8P+qk0XI5nIsJf5onAgZ4NrtpeAjHExaEglZx3YWt
lWyHvye1FYDcWUMjkjdGz8STH6jrkDGBln/87jtTfVlIrqq+QbYObr4lKRET
oi2ONMYInJB9vWf0yLIhVisKZdHmlRUmWd9Oh5eWBxKe0zNV80ueJGi32a1L
Xsr7xNry9GZ8rwbnazhWgMqFZf+0q3JkZfLL0/GYeFhHS5ehva2fpor75ERV
2a6vUl8Fh1P4rp1sKwI8POGISeEms8KE0KMYfOHxf2TQ6I9pt+Uhj4etM5VX
6uDc8WXPm+intO0tvPM9leiBL0h7Nqub6Y01wozDMn2uA//K/FP9j0RQc89h
fqlMoWsFwOJtLAGRvBSbfphFw8cbnOhbJi3lddkS/iZY5Vo6QPSZs8Am7RFF
I3Dspq95OW+l8g4Yfc8bvafF8/DN4EnpBP5SHwgj1q2C/O71evb1q5C+uR6g
XVcsGmfpqJ20NcFMcApyy538Wus84sl9TUn4NK0Clnjr9kvnyJ417+ff4oDs
v47usXf2alrPAokl3HhBp/ieLhspRJ2lb/e/O2cG4m7q5d+0bOL7/uM98CW1
4SexkseAtDvktYCExQQvOtVruXQxPKyH2T0CjKJ3A7jnmfb3UQqanV00j2JN
31QzOmkmd4mRzChuAD+1zJp5n5ULHwwRebDERfd5S1wC198GzCSBE4hTjJle
AZ1GDJN2dqN+tG83dBWdmrAOCyOCmmFKv9uNoA/7rUtzYOKodSxAjmgnzVVu
lU1IeLe8RUK/ELNLXVsqOxM3QyLAFQMji4krJTAcU7sjuf/UMi1aM2aZ78qG
ZNro5VhRWlcXfncgwpMA/FjORJ/q/19GEXLEZf9fXim6x6PdIqT/vd/xEsgT
fyfz3UUHbd0nkTinTO7kdzhC/rI+U+2RJzrcNynT1Hmym8x6aZPAPdl6PJMQ
359+vj2/Otr8pfdgVEUlqsUoK07zxCB7ygl1uJerprfBTXwhzxFT+1LxPmCW
rphRSZpnwUPYCHi2qKSJv3FuAI99NN7ffn7fFP3FRplbXUdfcqGfoSETZ3m4
28v4BKp/cryIGGbYr5lz2xC3PlzfN/hMOfOa+KJNQTlyt3J4oaE94+m84PJU
iT9/T6ThcBXi8g023wKyjmX/j721JzmDNznsHScnuJNwTjrmULIPVCKErKxR
YJweaOay28sOw2Vc4m62lirz1b11HqXKiDxSoDpWh5AGm4FBFb6hdqTYsWlg
liWOq052v3gewLLHl0G7CwRpUwl3U3mtJtQUHw+ZQ44EJ3RzodbuLeySZP5E
RmAS0fijJOoXvm+TyhLcuWdUnseZPchRYtRQn6hN0pDoA+LmwmwJN5edNJ2j
aedgSRSFxiyUrAausa+WzfdBMAZQL2JBSkPf+nlDSUGaZzp6BCtw6CVP15zi
21lHXRz/pWikJrfKbChyV0CJogpABfEQbVrEesM/8RUATTXKByzxTxJm7jdU
8eB1q1Wa5R5Ev9OsuwSQ5PVbPXTUUfVw9yq7YxEyVBLEiMojUTUPQX9lmpk8
bOk3Bqba9CJaHqUwdUwZISSwwZAsWWvRZFSpKj4M1O0vGs63/IT4X+qRijYQ
sFtnn+K0p3HMFVteFawy1iJsflPtvi8HdF/tHkiy9wObPYJz8pidAe8VWcDm
LR7xFJYr9jYMgn1a+rqfrCmRQJz03OxyabbxkqYTdAtGoU191Z6Q/EwzKodq
OH9cRmbHnZBCEsC2+kkmy6grurNuCVXlpsxYi472kk+Qm2JUIPeP00BBqjYx
RKbCAzW9rJ0AvQqn0USU7zLAv3fYYv0n1iIoeOQVIrdGpSqOHWix6AgDSXvJ
U+og72017pQQfJPePdbSE2LEVBj8J9MAkUOC5wFv12THUOOPegqg3hR3Is04
moyUYO7+RRnz3R57VykE/NWreaCnc79zide4EibltpZWx2IMpluAYFbHAKw0
ALp/0OOOn9YwE6pDxw6CbDusDl+eaOahNOYIlr+9Syx48c2m3XLbPZ62X9+W
EexMJgm6m8aPmBy6Df84Zf7U5p6wK6RiPgkk+0I+5DUkzvvGYDINTno2fczT
tiVVsJnFdfm+zVdVbIHj2O2T9+b5WmYrIGRDmPrLbjj/eDZbMFOY2EQomvuv
adSuHuYC9uJ4rrldmdZw6ek2NYRqYzdpFW0DGXONnPxNENGpMBhSTK92ePZO
e6A72/n0TfNuncU8cECnBeo2GWkh6M2U6HfyXDJcvBKAJtxxGcXL0ttKrL3X
Ao50BOUfh2bZpFwQ58r1QjCSZ+ZhhRB1fXHBEemlHQCBbmzcDtzyxKii+Dvx
IH6h0fsSXZLN1Rugsdksx6zQmCN64ZcRi9O5NgtsGB8ebOTTUH/jOLscv9G9
UENRomvdlPbUE2roqNMEjVZvVkfs6ZP/tCMXpiPgsGwIuXxJhxFbGOIm+bEO
byyU0JBz0dj4zsXE0z8xkC5sXcBkLNmkxiefWnM6ERiB8WHyCUl6Ybr11pY3
fUb+7FTPCZn5AZsT8Bs0BBq31oKOAz/EiIJ5nMtoWFDEbsmZ6kcEhsGhB8qc
KTY3CpI6YX0qr1RXZ4kY+G5zrFtA4e5B0imPN5wqF6//bYjqfatYZaCg8Q0O
62JclMv3am/z1Pxbt8Ann4Nft64709jjqAuNLKpLWUNsMhGJh6sGJEhHbz4D
DUeDtOPp77AasyRvPlcxqg/X88b5aYLylya3N6190cqloJBoeB3LFAOX8AY+
BbPTrOwrKKrc+G+UQt/HJBux38DDejFBPa8YYWy5TFTpavx2aQqpLl7pamY6
3wJ7ETcV5+O57A/36EBqeFNhp9GEYNjrU/p/1JR04FCf/spUggMGZir1dhsX
2nOoJAfsPTBzPa24EYINRZcBEGb3IAIuSThPfsVADV50B5n2PpB09hNcAdrt
t32UzUPYEBQqQkXL6vE14VWYZh5lf9N6pQiU+99NYXmRRVfJUe5JVTZ6djRr
Vw2LzixrGHwwwTVTa7XBrO00vv4Z7nakvhhxJPLFwe9MuBC3dqwMp/MoWGP6
mMlRLPEdu5m3UyGEUDs+dH+XmG6YSldga+C6WErwWgKpUqKLQ9lL41ixA/Pj
DzF7rkTtk5eTb9laqOw5WRApZJp5CSJLKGKL9WK7xJSInMy1Fq9F2XsqxTPH
URc6br0bAMm2vw8SFAiByxmv4ffpG5SvXYcjHFVQY1ut4pMC1V5PQ7xgWmsM
Mfb+mWWZ/pNMRFng3jiQEutsTGRgSZVWmui98Tor0XlcZHtL+kLErvzcjqLG
2C9782aB+Zl6myzxc39POsMz+e3tl+HQh8H9x5/UwNrFONcfk0KMXxIKvqYx
MJsijqEsvEdjT85doCnRHzVKLH28geiyLqPinMNYVu3BbdkSGiXew2HXD6mK
6L6T2PQFf0r3J8RPfaWUo8RD2tfeFDivCP1ypAzInIpfXUaX6nE8Kl0QFEse
OuVgUJd23yt2+OpIO1yzkRkLnV1E6El9sHOsWcT2lio7RtEZaTkBvteF9vIN
KrgiTgDGYTFWf9f7+jAc2b4sNLODiAxBetm3h1yiDKZ+TDd97rpV3VlINmNz
cCbe2Nym566Log12+S6yUnltHqoRvp9QQ3ApXKOVxo8iGMgjRDfRf21OZSxV
AnIhKJ7/sNGOOzto9qadeRXMhj/F2g91myaEUHuSF+Jkucm+/k5e240o/lUq
0Cgd+1oAsBqjQWY/5IY482fy49G3K6oXJYh5dIp2PGc9DxIcvPryrepkOm3c
kNAPODo2aTs0waUUONsY0to6kbRM12ALmTfpDvw6VU0Bbs3G5NsDN4mv1AD5
sYnjrP2WiTOJphvPDC02s2gesl1yoldysiKkTWpLu2bEmFOAh9NdDGN4CnJl
LkXmjzmLOmIJJ5w1N68NR+azScGGKv4+ZkO+FQ/tsdRLRneXsAG5a8YD3K8M
esSs1LQEGrZAIPhPagBVEZ+Kmhxp4ZY/SXLX786h2+HbaPQzxbUwksD6boh/
Tsf4j2C1G9vjFU8vIJyuvTreZPvBCU47oE9qrbl03cuuVenwt/AtWhkznou+
z67qAMUEn6FWOggE5Jhgommn0muZ8zajo1QDKV23KVvG12SjkyOeXNDxLE7k
Bo6GA2vYj8VuN68L7o42cKxFK3pcv5706cwCzaw1DTGnGO2WN1GlQcGcvN+x
MgFnz93kZY6elSIlKe12k2abXlDtJM7ZFBLKl451Xc/0mBluW2iMO734+00N
qoWr4Q01ClD8TbdDAbY7B9esMhuc/aWz8jGYLQgZ/QQ8B5qdL2sMah8UlrmN
j0EQO3zHRJW8YO3qOKcOz72xfz3g9mZ6P5Owvf0EuLV51YfiB1NtLsyYiX0d
LGb4fhNwcTh9ITyR12wKu1cHZCRv1UKjaNHtDJmugVlLVIVr6hauyvrSnc2Z
kH0dmbxN+gCWzAiGSc3/gcunEUuMTabIVJOpyx3s9dTAfvnd20BeCgut1uSg
oXTTCUz1dUsEVU0SwS9DPnfhxyjRIDugamV9wVpSl/k5zt9L0HrylflMZ0sE
1U1QT036p/3VINlIG6w4BL8If7I99xC1Bye0YiMaErMStIQU+hsA0lCWtggI
7pZ0biIPsScerV82veC2BmI8SFISYC+mIxN8XkYpIqdtuHZhhAkh0HqQV256
+BZ0lcj6jeLxNSkXGcKwoh88kKPsmdemIGsA3q2P3hAttXSaMkGzgspIq4f2
XGAqu3EV/GoXpnu0QPq0QkP8v56/pAUyPj7/XqSkVU/pPc51tWVFxqbDCA3J
8EShOHcxwPlh4l5fGaFuRLKk3l3PW85TNwPj8pj7w5/Xv40jCDXFkDObevPQ
UCQhI/PdaIUNhgWZqhJZwt65a3CN9ht2U5hciNRLDueXwhUiMwd7XHOL3Bdm
o0nBHj45AWa5qiUyaya4NhiwXClN0t395cHmNM7BbEkNg3sWBCf5+ahS9BM5
6RI27xpVNsMtACTrVi2R8PuNwtKN6QpolpjzOLRkNixVR4yniIRGM4LErLuA
I4XG3JxjX9NZBjdo/xmX8zg3Um86IIiFAPR2E7wd44rxaOBmmqqb0M9sE9ir
HlWe/k4RqxZ3Rb4PWn9ouj31d94cGtXcfNB5GV9yv+DnHqUVcCOmF/Vayp71
4c3xAzD9BYAUlYuL1hExgODr2/IuS6lv+xs3e/QD4iWaUeI38CpEF35nplPQ
PWEldhVTHChjar7ozuil0Q6xrpUqKqDk0WwXc6aZtEHWLirzPRoUxPfv8PA7
/gdw3PYLJH1LKMtK3Ktc0z9nd7d1GPoQI3XmmFVOd9kjCChbEys6fWw47z7s
cY7Ot/tkHIa5hipbrNee38lsQaC98+55tf7et0VgILpi4bTzfqTVgRv2XLYm
u8Yabnkjgh6VaB4HmzPJ7f7RIPmodqu1TjBz+44r+5unv3s/hINa05aSrd/4
qqTMttuz0kTWNCun+pRZ9fvio0yr1oV32U294wo70R3q8MqF/ImTEulYRWWN
YJcaTTPXKyZqKLVBV82MxkOYVbEXenshXYzDC8fZVX2Ru2NR3ELL3HZwWQJb
c21Xc1PU4aACIUSUH/4ifXOTfbpXuPk2LgxFPICH1mZq0gUcGAliuTrbGLy3
TYi8PgH1ySQ3IV6mM+KZtYaeyZJ2uJ9AptECAtrZcyCyy/oQAEA6Xb/9bE4g
nApoNppmVmTZwPBiIw7SuaN72YVTExtodkD1/KomaUnpevyzsKDlp1fjv7Jh
9Q2jRvFJuYqHQ9o+34TbmJ8gLuubscqXLLUwHHWx7jPBcvAF2EGuWCeWJHTE
SFmS2vJ2eE8aopxfv6nIkQHH1g4TrsEue5tW12yT33ozaEr+5oJTCmKZ9ps/
M7ZzY7WcS+Y5xVuD6NSBKR29M943sd/AvSQXRfe69F5mkYq7o9QWv/5+Asme
0QSwN1G3koQ3ERPqCJw667pvkwVz6AtLyxqKg54uHlOd562p0wLjSFhkmVYi
S6ksf/zps7XsUt2WkUqrax6ojB1onaTfKhs2ZI/9AIrjjLIsCTeBQyJsHGHW
zseUL5aOIB/4rwBRNupDSwdqvUjRIQCsClOZeM55qMInGHX4FQzxIaUIYg9S
MgHR4cZJ1GVjcUPdeigCHDA3gaguilen15i2suY7H3dUhN17TUW6T2iwkLoD
lbgtr9XLJZ96pHNpOTfEWnsSBCL+FEmkPZlgA2Y7faLfcDNLn6JGzn9En75j
ciXfpPEzwvK2pQGwxwXEoiaYDQhlHxfX5q3dYoUWonvVXKdWLoWsY+73bVAL
Ol3EGkPzSovqTcU3U1YdIA6wBHIk7knzC8ATfsN2xr38YkMOeil8VG3vQjbr
bh7Z3vhrI90okN7VJZH4fJz8DLqmI/T28NlvYd2idcTjQBGmjj1TlE/MA/4S
YyI1IkKfKZkvIiiPpM4/VlJbnwr2c7Ehb34mKK+ht0uHSGTEXOsi5IOWuHlR
XQ+pFgaMqWd/IDfAzLQS62tbgKV+1SWjUVEZChcZ3kg7HjrqAKajEjtBqq7a
RySdb2ex/fVqvtTwsOaAc0OcBiTjvPY7jpG2UFtYeht9UTS4TJkWkOEeDvS9
wD+nblwuKdMKH3Mi8vVZVASdryKn1AFq8vgxu0VobNZf3HHdFk74NWmQ0X/Q
tZxzn495jsM56dmSPJfhOe5Xa4+eEES7iMojhZCcqvvu6O2adf3TA3XsUkvq
rExfeuzg4y8xQ6Ir4b5vbXltmeWBg5L1ssHgIbcHqkZRTDYAuHbV2E/nCuWE
tCiHzAnFOS+5O1AhP6zGtvoCa/NieskBCgH9sNbGPiCO2QTo68tdzguXgLDt
Sk+KxfMIAZulIpAR0G395jDdrY+4MdUwe+qFMTKdUn5bpJYXe5HPwTarbSlL
4Hc18CrjcEbS1MRIMmiqWaQNdygL9hvF8waP4/bumnP9U3Kq4yNNJiNv1Tuz
h00fyfET/k9LfYoNsjFqqqKpAdKl7qIjCGDipb63QVftc5qoiZ9hwCtcECmH
Mk5AcgEfyzxtp4ihlmxaWYAgD9183QfnPj0/C63EnEQMaN4Fe6LWuh4oATsd
2ereB6BmV1vYjofprsePjnj3lch6B0pKow7o6cWDk14Ljjqb7nWF47f1Di5g
NA7uw9B0nvrrtvIRuEavEpcK/8LcknL6oSTTgWhAISKHGwuRafak2KeKTuSk
ZRsvRXbLdjv/cLLPcfh3s8k6CCDChRcXcz7rGHGiIkZidvj/SmfpuqtgHan+
5glJ2z0SDdqd+kqcQJQyQV1IYSL6nxXsqB+Nllq3goDfY33wEH6ME3KeW0Xi
TrQIRpfqAwBAsQK1jRC45UcGEPs7RUugvs+T2RwoUJJX5COVMrcA28xDV7V8
2TBCxotgj5YB3MmHRrSmqwwUpujRRWoTTxbX+/soA+jgQ8Msnt52kla8DlZ5
cTYTHelP/iUng2Tb9UH6mFsTiA65vkPA7eLpegQmzRlDQMM1pYMUGQxsvNyj
HdluJBlsr5xjLX97nK1VvcdNR6XwU4ap85vNVN33gkF05F5j4mtb/DnW38vC
DgHUgTG3N9ISonvIrYF0W/xtBXxANrvR18clix/rY544QBDODMYJRSyruKc5
g+uY6riSaybkZpnYDVFTSiQBEXP0cFk1pGMRkEKC0kMUeyLXMiyqcBFDbkZQ
Lqz1USTIKs6Zlypttpr9vx8AxT11r3S5GgpnLoMhVnpL8Y1ZF/fzLJOMPHg4
kaYQvQp64bSn4QajcEXUJddo53zQ4Z0N1K/9HrorQfe6W9v2m1A/h/4OJTiV
dCRQGzL8WWHWlXP5ATbgxkl+MCcCntUGpUN24fXTT0IYht5uE5SM4Jab2IxE
azHdA/shbKPArxwaQkj2IGEx4LhTrlBqFlyOiirfxEYSR9r4owExDWrYtbkF
7El0FFtHeMWx/w9MXy4QaTWElo7VVB2QIcYY0fioVi/+CUDzJ/fjHEP9qepR
E0OEje5dX2tagXJq+/J+j+so9yQ5Y8GAGXx56a8gRyfG9SvuAAMT2yO7hFlK
BF+jB1VKLtPsBUVJ2MVErlQiZvYJym0D6PnFYM8HW+8luw0eGHNZ0QOJrOA0
EbQae5ovuSyXv1aNlcwzG7KpGD6HKigCCSk5z6Vl0gIyHPlT4lyuYr1qmiJd
yVrhwWIA9qMNznYEySIZv5aw1QTY/YUm9KfcJVWJsk0/TtMx5A0753k3/40o
oIlDxhYXYdOP+VzV/BOOb9t/Sf8vIqPLZyFcrsLKmTunzY+YfzfDBenqRweX
oENsTaf9FnUPu83rntrm5HCRtHnWgql7fX36wzEILsuf1euYFi28U9fcXQGK
AVx1ha1+MRTCkBYSx1tz+9zsTQo3lrqn5gthCCzMLHjZBsajk99qv/gInQAw
FMVRDnQoxv4+9blEG/FOVEvwmDBYcq8umlET9dQ5K8jLAXAg2FiHtAsta6rg
JWB7SVkU8AESBuplyft26pqcFOTqFEy+vbu8oA6yZ1C4ELLfQ86TxCZCcoMS
FZcAAQPgq+TDuxJXrLFxYOwUL/bTshuUsVTjzcIgQqBPE9yYWUfVq4RbWjuw
0Ylxvd8CsWBjNFag4TL9l+URnvdGYWsUnl8AgfXwZ9JNofOHEBd5EqOcA8l1
7bo8lV8NCEEOscXBo/RvXU1O0cc7crly5fFALtYMju5Zh9HNxSRwGuxNFJuU
D6B0A9o9alwLMLUpt1UUxkqyFbkSC/03etQYwd3wple3qFLdH1rlYc+Kmy6X
jFRB2s0w7tzZk/ZHYGN4aHnhDYd1I0BHl0OXTq0IVtj+p6NOrzDdXxPtg+Zw
RxGY8AQbRGf/S/CBY5332AkIDBsu0q0eAR1dSnckerNaI6DqX5Z84XWd/Iz6
CoGs45s6GHvS9x3eAqifzlDvajnP3AqTT+htaPH0oGFLwvKke57Lgs9cTQSd
IicMBUIkIjJUizD2R1wOzDz7ptkCeXX0m0l7JAtdQ7z/X5M6pSjO/3bnPY7O
ZFcsPAj3mabRWsRTmGQDY4k1lwpq3+x38zdao/WM2HWf7ddgPxtNwswmWCeE
1bINdUsQdggWhQLg+NtDFhA+vjUu0clklLOkz1cEdpNkwN60p1lUfEbfBfPy
+dLXaXiDM6yT/wBfGdjV6DjZL/6/Ah5lLdLW5MWfJD5Id3Qh+S+j8biSEkvY
fxAw2zm2C6mEt0nTMZ7nZnYpUaGjZqekiC+d8C6NmT/KLieJmRbrENAIILv/
HGyeYDN19SktPWy3uXjbXPGqDls62bKILKQzwFpPlavtHySXhdJ9AoPHePH7
drkbFszq3JNI4eTl5UDSdGOUVHrT5Q3t7Tq3qmaq0qytcZYSp2047wofBpZ6
vOHV+hKd+BZ+AaUR4rIjZ5y3IfHsMdZiHpd1J+RKtmnZ4pgJdBymXFVXdte3
/QZcK8gDatMBDRpQpUXFDiujUD409A37k6reZGW4QvWSnn7PZCMGPXOwH0TB
h6IEfIji2X0qBLYoWGP9jiMv0Cm9q9vSAfA0Ai2CtifOG1F9G6eZYxA7jVW+
hL3kBm7XcUKrCXfFTnU6PaiL5NpZYUVeyavFcuHsagNzvfoVL50/Ak3NCIWC
l+AmMbg0qWkDkhfLN0Xsa/Unb2xrcvKh4cj70KHoAjGTKVm1CTOEHzSvxFmo
43FdzVzPS1YWQWsYLZLMcQ6jbjIwugUDip8zZpI/+wojUh19Su1NAPVPKbAw
wNqqKKjnc79vTBmzHAVsz1YL0nx8z49rsh9GmFAiT6S5WV+gUwCZ1FjRGFlB
O2/CkfK0FHf1mgJDwL/jHCa6d9FpAZLUur8QcjZo3W2DFZjdnHl4tYwr9PqJ
DG5qK0w7J9HntBvuY33jjYvyPXFeoRPE6Thd2MIwnmJ2PyiLzccwjUXGaGCz
sYtjrsR3OAYqWpF6a4hNR+4rrjCpqJdvRxSUqGiFzjVnIJGg3LwQzU/ZBnGC
2WmCkTLgYaC0dccNVNP6HQw0ZE10nZsnocMiMeZzADyc4cfAooQvZ3p0WI37
4QBNt9vI3LTXYIH5fw8/Zoy6mTUSltt2nNRYS4FOJA7cPlSppsykhWN4aa3A
IF1VCjDetiLJ3+etvIc1SH3++5ExkFvhhtayITPfIDRHjmLs9iUZnrwXppMk
Owp7naS+8teFuhTsvxsaaZ/HjPAOYpwzV+zEbR58V/fx2lc2hFB8Hycvm+Ro
YfexjHk/WbQnU9eryNNWKMZg8DAJfgsIEKAtUbjnQaq4gHN1CBicnWpKcd//
fqyX8DHRROaDqNRwrmJRg9wWU5WD6xoNSErYcvQ6ZFpzkYEY4ntzvhErizA4
lL7yDrpCZsVvilRdzJjVaweavNYHjORbRGQhTQTOmqbV6E61kHCm1XOrbHMe
nybaO2frIcWJOkL1YVybxAawwMZUVC7RgaBY1UD1o53vx0UQF2LjV7FHdjYL
xQw8EoOK9tbwoRAlZFXDxfM+kDdvUKK/7OEOLMDdvE6EGyZJOCBGJi5Wyt/x
kmvD0oDKo/GraQMDub+FATKHChnz3VWqLX9o2kaB6BcvBp8pPNxCu1KvaUYc
J60MQThhz4CqohZqnggQJA6RGiNy2HYPRptYBvtBW/AzLS8S0C/e75h4H19Z
TDreQxBvPGcpCGxi1Qq/0bz+13qSAtBjwGeXB4ofYZnILBRNb66ugkcQ+Er1
91QSdk5rexq8XyhF8LvWsM8YGp6b7Jgv/rKHGpbXj6gyXvDgUbwRX1YOlrSL
htM5sbt194mfZZDg8G57jrJGtF3OcCi0lqW/uWiRD3H+9LXVTnaIj17no++T
oUsz1EK47esh27vl3AlONWLRC/QXMVkfvGWtyaEoBRAyFEq4uuyxUbIN/yQd
4o1RAOd19HPEktzdpCodQM9VDe+yVpBeKsSc7XaTdMXrxljPHK/p9JuWq+TA
joO5NUJsAVrLW6okuQiTm8kOFWrN4RIWCU1NZbO6milM7RaBnSa7My3Ufvn2
Aw5YpEJ/cxMxZp+v2TPaKASlk3oo5qOrWhp5b1C1KgXMo7/qkunlKtmuBO1q
aFg936Yva0PPlbDH1ZQqbvXJ1NC9MdYpdkKvqs5+0fA5+q9YWaKG8ZfmXFxm
w5PwCm+x+HHqrxfbnuDVrTv8PmQ+IbnllW+C6/16UtswUW0f5Dwl/Ca297A4
aXsqpGZs5lCaQ6+jXuecDYhdfnBC8wNX/svMqqQeys5D7osj/maZqr1UL4JF
35qlSGigtJbBRSFtCwkY24hlyapOeiwgi9yOUuMwQGLik4JpG90zdIr8MhWL
EA5HUtW+lX5JCkoWwQpXaWpViyMEklfq6zaAhoaRf8w742cj+YLk5DM8elcv
jNT89Z8k9S7o5rTFGN7cbBw8JzEM48X9wCaEoIsS6EJAfWW8gf+INU9bBb+1
mRK7+zwE2jdGrTlKWjX4uhX9Sx+/bOWF674kCZRF2tZ5OSdDS6ZnYcCypuCY
6qcNuhfHJTSSnSsCk7lUc/zCqE/dCdMfmLR0whCi6H1cuAFhGtbe2m8sYnFE
7im8GGQ6RhqgvJjCpSIzzZ+484aVfLaB2T+iWt2AhfTykbVAFwn4W6yuYAlR
e0mEBriSjj8CbShT9defi+e6nu7KJc3NR2BNHyqc2pjBxE43D/f9NPyAr+qn
sxMWYrSBmZxTjDSfLhXlP7fCskreHYgigh62KCAmllt30mUO7Ls3oGveZWig
euAU3YdMF08MtBg/Kf3q7fKaTc7qnbGYb3oiNxDZ0q9OV3DYaI9iUgO6c/LB
/3RCV2gL77vqObjU3oY7hIkK3PD3HmIhouORrGLUMm9WElshOTp3WOQvEtvf
asNLASbXP6d11B7VsLZxLERaNqhS+FPKem3n2x/+mMCIaLMZM8AGoNsbEBjj
JFOLFCwcAvgGa0pqVgc4fR8TFZNqhDsp2jPLl7uudcDXp0AEJbb2tBIVDvQN
gyUYOLhPrt3SU1hpCwbAptOm/RkviiREiCcBmpGPSfYcmUcUKtfwwKoslJtv
cRm7sl3FrbzmXV5hHHEeki7JGguw6kERJRC1k7VU7QnwWQXaFJsdNtg2vmj5
1aP26lIstO+iO5pdrfxZwidHyje4ytPRYZrBv2cZhAkjjXscp9XFYQYCwFQl
M2dBn4CSIzm4b8YczKXgZh4AIR4TdlcidR9xNxoGMpHGW6SRE7N98E3ERqb1
2KFWJUGY2zhp/FUPvZDOYECINP5G7sYRVjc7R0xwOOWPgoXwV70ES1AO9sq+
0tcHCWMyp9NE/8NrrKoZxKeGCklig3qXiNONHE0okVwOdHaUw9nva9ZuiiXv
k01y8hhwDzGEbXhxRVFizXM4ZYoVxtY4HcvtgCxaOYYC9dExeKMkMkPUBY48
bJ9CjHb6FlABkqk3WuW9f+4rQNYcQLfTO9TBMEFVtKLveHC7X3wP47tELDAG
Nx7ZVLti71czftr/QGYZYRF95kKb2MPvPtgdN6Q1Xs7t3RvfOkUvrE77sk65
t0gq0gNIZrnAwYDDABm1ys1y+ivZcqvrckThKpYXqOswDYVoo4VZ3NryNSxG
Ha2pF8wwFZe0njMa0w0XNS5xT7gV5+LRSBaS2R8nDuM0zhzV6LiZ4AyQrIP/
V1ljkaZXjWZsjwSlb1sjgivMPoH0w822tEYRpEOfCQ1NCabZdkfg1SUdN91K
Ez7gHaw9j42gdADZbg/MhFIxhzKJVcmL/nFOUaatVMuibFa4ebSnx9iB3TRp
bJN717Pq0gfLqjw4te/pfp/9hG4FuhlXjGXh6F7/nk7QpyWGaAg/WMHB8C8s
EBLKaLl6T7SUiwk/gBAgTL7AtDBlQAt1Nq6QAfJsBQSuyjG3KJksVncyu8MC
sc/RW7klbak4+a4j25CcnTSYcWmLjpdgRuz/9vVEBR/Ky50G9TTbLxOQxk2S
LMvXMqL7Rrgm2xuDXetvLMLnn8OTPvvoseI8S4M6Rpl7h26IkO62IikYHXXq
cUJQTMIQ6R8fLhJGDHKuf2EnFoq3peni9tIr8BeQiWu9QOpjvzhVk1nFCOrZ
3U87pAOJ5larSrQngRBxMkKD9DQSSBt5Z5K0esroAbPkP9TqttemP5FrUllD
axvCkG+yXV0dGwPTi6SPxAuP+ZVDcTIuqkbJBELWwxaSfPDpAyf1yWl3s5Lb
13d8PyCQY+dcKsOKDDCNwK032zRVyPps7w4Zm5T2WwtQilihOQnwiO8NFNeo
LQy+zFlr/qSNMLvtOQgjF0n0BIjJhiofbYT+dFTLbERnlyOlK9uQdghJQaFh
RcklCgpvlkt4tov5zrJsXLZlAKd76sXO0NCCnHfYk3xbYS8GY0ZnIcNTeEMF
kN1LhISTVgjkCRGNaTYmrzhWyP2xOd9xzqp1wd359lu1N5e3KnDdccJRpMQ5
d5uE33ci1X5w3ozISESSIuuhYhFBgVqh0gE4hjMwxpyt2S4tiXR4ANZ1F/Hm
kMgzpsT3qDOMjndqL/ECk+1LgpKgQMUdHbDYy04nYBFwlJK/6SRvMkJ2w/Q6
Iec2H1zftceAlzXLUaTyMYxyi7qG3aAgmVqHeUdPjftJInz1mt5QjeNQ+HFl
IJNVBFoWbkvQOxzOHUHMyoET5Eb15bBuFrHOf9oov3hnhZD+CHLTxDEaWO/I
2M7UC3N8VOgdrHvby4xpjHwkr9ToWYdkmNiHpP8uYqOt95tDpOxTiQU7DEBR
r+A4IYt24nmTNXhZ/3OfqAhY5/UhJrNy7BrafdNb9M+lnupH7A+sp4Lqa0Hl
14qIwVBXj4JWyfm7qqBXl7SnKKrhnAbw8rtoMwZbAFC/K+pHgLoLn1ezGmeo
YNwHDXAk8BgwCxEmxVXisOt1OoClwIVw3438NMFFAtmdawiVlSuhmxTzEWz1
beG8vnYPjx5C2pWppWOkxy77AG10qCgLeRygFbIQjOQIQTHQY6mnGBwvt+ka
/+reNjgY5V+gTdqYZB4sTHU6SBHDLndC4qQYgu4AHBHoS+JbyZjH5L3UjD2v
Bwglocrb6W3ExBBkS5WAynz4blsjtvk+lBXRYZbF0B+klt/IhB3VK4Yu0NYj
gREOkeCYdkHHTyUOHJnYE7PqPy6VCoKkJyHGNSj/4o3BlrJhkR00Z3Tqwgpt
AnX86fWhIy3xH76Guy1MgDbQ55F6gUHwyrxpLZ47Sj4ECBRFXPcbzXh9en9H
Ds+qrchp3MQ/BoQjuPm5JgmHFntP/LH9gKCLXA2WZqAyMsMaGceY0PcwVHx2
8WWZhZ2qlEVfCWBSwez0/d3PTV+D9Xny2vErKBZPEhlguItfcQh2wN1WD/YX
5hSXTri3d2ujAxH9pGHxQn4mfIt0tmAzrUb9j8eJFHkFmE62NsMFXQ+Yvt+a
LRh2uYSLTiuZGkjW8uD+p0UllRH90IHxNBdYkllCYOpSxpSEdHTtv2kyKdbP
jPsSolbIWM1PLQErO8isOLqQTyr8gZ+7kyEyTzOtCHhlerSpramnSCz+3QNF
hm4Ky3/so9vYYZMeCnYmLTdHZuE1FCRWLdT210O0dcunz1a1S6e96O54F/4B
VJIIf93wWot+eHavc5OBAALX3/PnSOEXMdTEXN1UY+/rYBif5/PSfKjsMnGX
Y5XJQm+7+7NfdmLDLnxsaYR6n6pxR05rVCIDeOCJhEXBg2Jcxb9WvfrNB6F9
ENeTH0ZP31yTs8axp2r/PCRxP4JMyVW9BjYi3OgZ0bPFQmxj2s4ceXXl/mA8
kSADQhMquw6W1W2N4xB4OH6eaIu6GRvrMjraMe3mlU6prAAqlb3agkXvPWdD
Rrw1P8lskV6z3C60lijkPkz/z2oc8SMiGJm0IpYv1tcXgXb0Q6KL1KGHCWJO
YMOkqC+YT51GZTr1othzLDzIeLVzpWdh4keKLnjKTEK7GxTTu4vTCiSsk+Ya
lQgdA9y51eiXLXPMCD8RaskeNAh4tJOpfvL17OBL6ZKgb2Udv9GdSqTNSWMw
FrwSyGrocC3JyG25+VKlqSLblrdGJ2IM6f8zmvUhrrtdNneOZqgHUneXREsd
zs5c5rhYxlc7axUkCxr/HRnCevY1acizUAWsL+wyIb8QXMl0j/alSFZHknRn
hKJwCvE0DDW3+HYgnW2sm9nNcIyRfG1o1VBiOIg8lVC7Fll9Lpy7qq0DM0Q9
2gLjC8UZ8luYy15+eNxYvBR7PxRhq5EpQGuCG7Kn8HPS5y7ELe4ghtFLE5Vo
hE329yyCBTywCQZ4p0dnSxkHlsvfdFndd9bN7wuCqv6gnWJDIefHpXy4Ivo6
BwQs7tLW3qOMo6KLQZtejzaCS6Cfhu2sqUr76O9AP+ZG4/SviRBFZTAUGNGM
IE9akfOaWTTW4e58E9Vgbouf6rvf1Ro6x+f4rKfxYGmNFNOA8TUvsIbSIR5K
ud48AUUp2uoIif9cJQhdQFDH57YiQWYYZuZR6KP8b/vjPwY0Sho6w98doxjT
xISzj+5Wz6cNmbQWODLY7L3GzgqX6VwbX1RDL1qh1Q0mvhXR+JZi0qsq2xfX
LkRbYxDD1dDv+TUCqZQ21NxtIrY4xpEcvMXCLNi8OYffdf0SWDC4rVJ+fm6x
YPEizZL+ul19xVHZR11daCcxiJxoc0JTiKLbv3ZJQceJU82XGjBaXywoB0Gm
7AVvpyqV8lepF8b4BvfJOIkGjLxu2/sXOEMMOdicqdKR4/NWhl5WoTgpYFrP
VQl/Ybi5HSv3cnQHv8nuZHFw/tmKXbVdJdMSdbY/Oy7QPYibZ7nKF4UnhLuI
HxWnsD1YfL7T2F55E3Y3XFbzi7+6nFislNWE5NPVzstK1OQZR2fTolxMimUa
NxCKKkDZl54IxHpdItmBhQXjFX8bV8krZyMZuzJ4xZC0IGaGL3pWFXx7fwbM
KqmqPXemU/JnKY+PF109Zm1D7d2v7yFHN9dHjirfVo30PSoylFwlHmA14SXI
Dxn+k9wvFs5NK0wCw7/TWuY4pe2fxwznrAp0h4L8sn7stC1l98DlvMxhQwr7
J7n7NUTjKr577muDpT0jdbvmvHj2RatuUSsoSjxZ39gUan1r4tJFjoor21Pp
8yMrlv5963Wg0KF7sH6hGmugfn8/x5woiSObxn5y7olpLzMgtfQvU3DSMBtB
UW1cSklagtowSL+/8OWb4mr/VK7avXr3A/VFXQ6juDnG47fZ+PtGNmGr4MuZ
Isu3xWYJlv4Neppd/wC+Ghtn9P1r0pyKvTGCyj8XtkMe/8N6v0y+uzjyIX05
jp7r5zC3yK9Pes5ur75FPhCyiZ0Dg8FpYXt0iDyw5cDmMAQ7TNol1DcihzZ3
9VkGFu0qBvhBccd5CZOSkivBPt7UjC0SP6R5rmVnOUTHSdHz54WillKVF/kD
A2brEeK1y42A4f1M5NFt7aTBbdLAbdNEgnYxJJ5h72piFA2LKLWvd8CVgaJC
W1hIPduUVy1JI6s+UCTkN9TcOIqfxsH9z7AgZu5k6ZVm59u4u6oD9hYy+ajt
s4DozfTXFzxkXLRQsQXrmuOowJDByylLVeF0WNlxgi/X39qjKwLV60ZIos2D
gTYsb6eHySGuhdcEjPZR/eeCg7ZEhfoYQG4jmc8/bRPgcDhtRaVMZV1mcPRY
xbfmK2vNAMn3Hq8hIsEgeT1NLfq48zu28fQPGNEKEknrBIpx865EEnu6Cbrh
F1Y+rUKyR2ycIvVVPXy6w4HlDpP2NgLulCq2A74BuVAreu5yRUAyK0oExItU
XhtfZ3I94i5YD2OeOn2tkrZsMGLBo9rPeZj1lhxRfeTH4K42p4kfR4K+Z+gS
e+NqjZuS8Xya+3EGFH2GT+Rf8BlgOpg9s1eYRBQJQKM1WhPMbzooVvPGb8ms
W9VCyspihE3WLjItKMJ9KD6T97O3AusPpRlG8KCkfN7ErTGDSmEp3gBiuGOL
NFS7fvEE+4Yl4eg9kc6lE3+KoStAPYTOMLCOQElpG4k8l6DxHQnXTgh9yFh8
Xk8GpP8PlV/Ss+wZi9iDUjk3hMOi2OPd2d30zlaMzQLlhzdzoDgAXN1bmR1r
Hj0eOctVW1vPW5i+DzmONOfiEj0nLIKqwNx6sTdJpWjp0c4r6XuXi4FeZgXK
Du3wPhqs43V0LgSaCwEIzDqwOxUU+Njtr2dxwG8zBmQqHqvq151/SE60SaNE
15Hb0VJoxU0ysnPFY28BsXFxBSL24kAruWVqaNkOZpLS94u4ncNlWTk95dax
bxokdwZTfvxUnSjiDLYwSszsLrOJWsCpg6R8o3+hd0phX+9OQCBrClQXhFbe
1t597Leo9bIEOv+M72Uzlh9dcPqKrK7RZGMGcwA9PkYrnEOjART31NiP2y88
JrDhlPrr1i60HA45PWsrZq1D5/GPNcvcFbbSTP8JMMSZCA9AGbDwkErcsSMY
xkxVwUeFGeiDPCVP4kVHvBROBNahNjgU/Ywi+zl9gMi/I1hy2vNjZ0EulvNg
SR16I30UPV8AkztBWSwO2e39tnBnH/VlPsDp8fyljR1FqD6jByvCLAo0jPts
JLXmhLmrxu6sKqyPI8IlLscYLhj1GJAfVy0E3jtbFHjZaq5kbo2z87Umi+ne
SPoEBWFrZUWE9kTzFxqraHLPhbyzFYtkmr5C2L1ykQUOs8BTKAR9rKBdXnSh
ma9NiTUPj/VfdF072O8vRWlfMzJddK2eM5KVpGg2OZqaGKG2bUORrhKn03AB
2sDJjd2o41poWjEN1RClkz0tKgJck2DooHz+4WzYwP19T1c0LM9hIwSxx7Sc
+fyCGObUmckEBzhwzol5fxdfm2VEiwVRt86KFTyA7bJDDjj6RBYUDwTenLad
gh0Ncclh8P6Zqy/mBRwrHNc5FZvvE9NTC4tXlrpEnH8VeW+yqpQhW8ycrT0+
0Gsx8tMdiATNLi+rShDw+otFsLDcbjNClIOiCD6J71TvIisF6fXUmd0z1sDn
nSHpd4xBoyhcO7O7ZN5MNu9mc9Rl4eDyjOoYNYvnA7Tv0CTgh6yBU4R6oJvw
2P+8wu2XoD9vHOnlu0S1cD82vs8w0twCwIYrMXGyLmTueIaMjst/DanxnS+0
TVpLP0gmMfCJeORqtg9Eutpbc0pKZrH22VkMxY3yFVfGMQu+jI/I9noa4Jwy
YziDdfl/4SM5q6pjHOT83uWkQ5g/S/LHyNHU6w5+ChOYlOgJ55I7+edd9991
hI+V2O9bNgmqiUJC+Q89tDChCejOaQQexxKyMoCFWdW+p1Z3bY1MOZ92GAq3
VO+fAbhMSz1xeq/wUnsO7XE3Rqpk/dgOKFZd3Cc+U4SfnOT0oFkwF9C9ThsE
hNLSMGel2a1bfQIiA/kxcbYqKK/KJGTIaCm02FNvZDxyeJL9CjGof7jS42rV
WfkAqFRQRmsXvfhwvjdurg3parJXWyh25cWaG2RxoEP3slGSLCQ5HUphc1BH
5Qh3M+i8gM0juefKlkmvpcK5zkMgIB6uW2oNPYkW5Wszy9ngoGZunCGm0Tlq
tDuRWvcc3eT7tYO2jaL2Ayp9FJwgAGwlXGziRrkaCLOMMBIzYJcf07mb6GCt
66NYDE396/U/8NtNGyNA1UQ1cZzjlTzNzTQb46988Ch4wsptUFPHBPxIvysS
q9wPUiJ662ly+7pHoYJEPJN/44+uxj6WbduKTc9PQx+tEMN489odogliCF7R
bSXrBz952wox4zL7kt31HL1lN0M2i+QZip0bX+/L4SszCyPefB2ipEdtn36W
nmkJqHxfKO8SvWXVGhFVJ3cidpKgAcxmGsSe/5UEL94DfVAkhSySqY4OGslq
WBUg9vqqV6JXZGYEeZS+dd1jKvZktIz1uNPloSjn3oi3wG3IpImmwfCMY3r5
oI89TJMK1yU+fpbvFMzgAFWjbZaGJq7FGhOpz0om1UrpMIQ8f24wIhHqHMez
Um3hifMBUacIci2pAbY34XI4f/lv256whgoOWXrLbkyePuSSEL2jfOsYgTVp
kKKMXt0/tXvyol9+YS3L1TjlHE3wHImcBOM5yWWXGPdRb7qlvVzTmaO6H/KY
8yfg+X5iaTPnvxLxnJldDUWVZO6XeKHMDUBs2aAHX+1EDD+2faWUoHq831fN
7asPzygMeCADtaQDWpQskUIu71iw5qQrohMy0hxP0nthWFBW5VOUPeQePVu8
eg7mPqaXg7whIq8eabZ62588ioODMJcSM3cq3kfRNIhCEkUy4neOfXjzi4Mc
msEFAnje5EUAPRMW0e8bzVPHY/UA10kzKl+hSOuBqWMScKarDXPL3nNdWZZq
zwoMbiZ4rooJgzzjjj2Q4ru0gm8WEJRlAgBsUWrKo5fd0M5C+ETQXZI5yqUG
OnbKaEOFSxFGOUpptDv18SQYZpsV2OTmFfqQr+pnOk5n0m/MmGKhZ7wzHtXU
XRL/fezBcM6PPuCBIcu2Fu7P3FprmKlRjzokxO3LkIDJrNbeihxAozN/IIs1
a7+txVoAzF3+E8qfE52EfdKoyv8O5aYm3EeKC4seEt+/Cu6/EENVG69O4lsh
eOtMVpZ4jiWHv9zhyfI6u8NlZGrF1KmlMGMwzpg5+CsFY9SzgFf4LzE8U9Aq
0/+VTgoePkhx80L+/6VMIy/XnCOO/jw/2v9hYetM7grPPSIr0OpiDP+GlHq1
F2WkOMmQOFGZjZsrnffBkICl7TerQ5J5rWaP17z7Ty4kzLhDQq+BIgXx8goW
/sJCUGJzHX+ivA3vGtwp1gCiqNBmoGS+pI88bin0hlGlS7GC4hVivg30UF/7
7z7MOWa5IJ2RIp0Yl6z0z7KsuCg6IsNx2quh07LiQ+7R58gtJFznxz+g88xG
tV2JJzKceoAwXYXO8DlhFtzy66mAwVMH1Cx7jYr+w8Uio8DvabrmtM4f77z/
35B8IrAn7wNnoXbph/ImijwIjw8JDYI68yLX9Tq5LTPxUr5PBZeZ7+V6EvZl
b7CAYHOLkwxLhihUq9ODUIPA2hw1BfU9mzLUG03HzaWLonnHlSdpsas672UO
Xnm0eAcT9uugB+V0PqE26nvt/jXleLhk9ebn1v9mXlyLIRXBTVuhwba4nTaD
HTceb+JagBA/31QX3FYjcL0gFj3pacDv6vtPI/ufAhN8uN8A+t46rOdHiyAj
m+89A79cagSr4/mthKoVY68R5RBzs5mcujDE2LF2jirSlu17B02zUMdDh1gr
lDCqex2/GF0mNNeUmvupQt6auZtpKa/V0/eyXoWF5RQoOt2kZLhU87eUObFL
L0OxZyN+iyLQRYVZZ+SLBU8Jls56LFBka9yvpcLESumoGi05uCXxLcxuvkf6
p2ehebjC4JVdLJSXMxAYxb7XzGCJvrEfMr0/GN5KvjLCUSZoS7xgzjEWB9ae
8FHcY+Cv0V0jLvoJY1or0YmR0NTbZtygkU1+ZikBywO3AfRDea2Qx73u0H7X
WWVvJLj53z1uCsOI6cHWw4UT/DDaCI3iJVLAbpDEOhub6cxm2fGr5P3Jb4I/
5fRmwI787zgzGctb6/V8Qr+0xEjGKwj5TYo1rwlKP5B8J3IhQcgMlGBwPa1P
o223iiBi2xTQEgzBOcUSNt82TgjpkS+AD2/UxXAZZhJY0oZUGCKMKrPFI04Y
vOdFlbvM86i9hz+imuYdG0Ab2QPstHZp7PX3qN4kkNDrhmCrTSvgN0QtLKJV
3wltNhG1IFOKhWaNJkBUFi/lVnO8fS/91sW4GgUFHoPOkiOMesrTbxBoefHK
O5Bg09sUf+IN7TvAci9YuWbnbqybj/jdcZ38x1Kx3xPzVOOKQewut8JzqKgu
oxPuLJObfLJz+agiTVocpkr5RKpEXLg7a6v8PcI3VJrcSn0c3V0P2gndnIyJ
RHYtg0wkn13/DRqrxmXtc7G8vfVNTT0HVSq3/x8Ia5fNI5csbKTBy5RbaS/r
CAxQ7ELkvo0rab7SqI9tXDpZSaTqlmC3BXCH8TnyJU3PgwMp6xyixyXMnhw6
Nh0oUNPunFEDgURzqycQDPaHP0s/tUF+i64yBx+NE5sfBHOhnO/n3rRouyIH
asov7ObQ0XaE41QSXgdrzjElutkJYxam5jfvF4AVvxUzNa28qavikyN+kd9N
VHe0J+rWwPTd6KW+xq1ax34ID/wnyu15keuylggBKkLM6sTdpd+BrUSCv1dj
EltK6JL+qCrlXbk4kN/arYVoetoiyFDwreLjRnmmk1mvZrLTbHO5UYZnVX98
/aemO7gkX4xEDEw4cJXuly33SAzDwRlrjM2KkUvdv2EVciKdY1ALFRCxfJut
mX1E+YCxhjK/vIw7S26NC8yKpFiT8Rcoql52vYfChVi/loqNWARVyCCBt/pj
pbzRAS2n/WRZUM3oDIkMd19Iw8vorOJadAkBRBNnBhygedkVwuXR5NdDc077
53ktei+X6z7tsTw8J9oVzMlW4NsOFb2cSBvMgpIGwaEAylM7sYzy7ouoDUur
FilctWMd83SSuQeOWzjgkAxDt8ggwGgPlS/g4qWD2nqkbC7uf0w9vayJlom2
G7eEFeQ+CLlxNH5o5hxAK+uU/WQG6QrKG98KfeoHMYG2cDVCTV64w3CbOn8A
fYynM2mwzNa8FIrkaRR8TYwXmsXATDiZMc6AhT+Zkk6FwGawGyWI7cC8U6Ic
AU1bF3JrXfwlnpR06mSNqoBhGnbTdFlQNKfAcsQL714MoZYHtgQCUHe8De6V
ERIMlAeYMwVznoC42pQ6qL1mOkUWK4NMrR1Q+t+1hFNtS2rnufuf30s6CAIV
x+f2jbEJvWibhOL+JMQ1ZoCxJOH+f2g7C1EJzahI1GBqG254h/GZxzRbgnZ2
QTHDK3qZPH+O0zvXUsLuFFf6mI1bo1AXT0wmOx4YG9C4whY6ur7cMqRe87mN
uj3UguKFXzSup2eJHc3oHZj/kmxNtGCMRg5SnpsLDqkj2Xuk0NG29+OHzYjz
FetUs4nEY8HpOoS31jxbfNcoWgSXc1DQ2u74p8XUQki9atBwfuaMbO0KyIQ6
rPGfBmMyWxZjcLRGrCqxPAN24RhUOb9nRzRrc632XWM7iFpOMY2dnHV4ZlTs
IQmldbsvWp02+S++W0cgtWAmzc2xiK37uv/ARHN+zqpmGJh8fKRKDMfK3nQV
5oW/lbrzf9Cvc3ilYOsIhNAW2C3WFmlS4atY6yI2fYcLLu0Tz0l29HZr4Xfe
DppBMfh4VKgH6oh4E4QNHgE7D+LKehPFa+LJidOq8RAGY3L5BZGC6pdVdYZ9
YUnBUi8oDPwIE8GHZBInwXwEOitvVf/qmReujxgKt6oXi1n0dwHiHgxbox6+
ur6eCPtl6LpXdATNo76IKb1ZILxpwZoyzKynUUCgbQUXsj3HUWz8HWfLNf/Z
L4RDfii1+VZF5xguSHLIn6d6x2tLuBURBoPz1FHWCLpa6KSpX3YkrbjMQf5b
IQ5ySrQeu2GnslfLtrVtuJ/QV0frFxJSw5LdKG6Ov19+mMgoZy2Fru6Dlbjc
elDLbNpOm7Jgv9AXTu1y0/it9R8ZcNiKPabJkDvm6kgMQfAeHJGaNEZrMWNO
mFjpVyl3Qz5M7Zz/OCz4G9y5+49acXFqiOzfbnsWHhJmZmZuw44IQ1ttDRWa
nPIT5NgiSuTtsQ57yR9rULDYm+VvSamgHYoCQl1/YpcM4uy+li9bmEJHUxmb
xmL+3lqkX6DHkIFnYObK2EeCo4Fdfxnf5N7TY42yQYwV38kW3B1cCpSCC+Bc
vstJw5Ahl8YElEBebm5VO2lw6U1EPBXr1tBtdob18wCT6kuct+GvfUfrGqBU
GE199FY+e0xzR/pSdf6B0dDAZ7UurIim23LUhn/iU7pSb5WZSv2SNkXoRIuy
+190eet0tEgF34/10cSDBJNqHxP+q5ZnZymv7dAtFLhm3jlqs2KHmcOArKEu
yp7b6le1NSNAzJoekBEQA0RlifotNr1/kJJiaNblEgYo76b6QY+A019cLQ0C
g0L5vB7RFm9sQiusAvqyCZcRWnGXO4l/3l1b+vO9Jjz24Lx+twtz0LCGCFdk
LUd8u7RxAUpPMmHo4KTs00/aAxSGNt/pk+EAqbM0FyKFWQufcwtpcccI6zyK
mvK2HUIfXeY05skAGqJEcZofFxkdk4qQJ20OiLJDmmxd2guZZhRRqvfaOQcX
TF7PYIfeIDlFUel4P8jrctKITEkPM6OePecYoWZ4YG26Zoa8UsrTlhPesH8D
ctqki7fmE4N21/k89iymcDhGRNlVYuOwYw2d3aYzlj/9poCj5h3oZHQQXLxT
5eyDujS+aKz/ZVc6EoLzlCLPnXcBuRLc9OGqVsIuJESAuM6ECaT7CqK9IU0S
bGgFKgIf80+iMC0FUi+Eq5UB27JsjPU2QffK1g+S2jY1Fx9ww4spe+8kMRbA
VHVB3u+0mLfTbxOeUFuEu0V65UVPq9ol22IsQh0WobU/vSQswHmNx1cciMKV
y98AHXa0IkbhFI0SY6XKMIS2zYu8Eb+NWUVtzJQRciBx4iIGM+tHmkRPbZIt
yoS3Rhl0qUjI3hGoE6av1BeDP1ln3MMvfQGyEeG5WmaBXJqBqz7OSBWqMSuR
NyBN4L0iQth7+5gpNv81oz97fOq/rp/e5PUYCjko3u5H3zIo6mk3M0eTEBYc
zgKuBeh3P74P1PnRvgNJPNL0Z5YCvSg43cB21U/DGxWTFjtBqPTN6DPt/Q//
LbTqavqsxn7pWjti59WKAx+hHIrsyx4RUlD6obetNlAuZFH/T5LhK+1wIN1H
g8+m+ZBUVcxHfhhxUgw3cBHWVkkc9uUaHyhZ4kGDT+B1gG56vgwBKQ9qDdJ7
Mmff4UB+N9FlRPJow8m9ANkIlWlQD+m6UgEBmvPLfmUJbXwZmwp9ctNkR8Ey
wv0P33oHmIdBiD6oQ9zgXDf538rBm5672OJ2elUVhntFEvpTmPvSvBaMY54c
IOTuDibossi0fHMnnGgo/G7sw1U8rSrQAh5zFMdjRQ+VgjeZte0zMA+1QGdx
2OlGoJVVyfcZBP19KCpK7qLW+sy+1p5zQzcocfDVl3PIeB/aDq5JFlGzIWUT
rjILD4Bh2NVa4x1Xp/VfNP882EmUBsFk2oGMbCNw13NZfMq9eVCfkEmRwBem
cd2RgMi2dbpUsrCjPENUgq0bxEAwZ41IeVWffURkLgPZFutvp3B5wYcdrrQd
tsPIEzXw1mTKltuZrdNIfje593ZOwh3OeHQPnmEpcCDu06VZKFD0vlVcrsC8
puGR3pWwoN7XUqtpwkXXol1T7cIjc1LvNGjo7L3ab1vvfUYgG19JNL5xN+ky
Z3wXug5VUxM+FnBEmQT5yw7csC2T+YAIIPZ1WVptYBhSJiygRHQPVFssuo6e
FHgrDBoVnuhQM6JSUKh0kR4tP3OdTz+Xq5zNxDnFXf7OjZOaGCWSx4jmCkpN
3dyfy5uZmP+V+5KsoPp2P9z1t5d6kpZ1pLs6Xdm1sSD+/7lMAaXIVIyBD60W
QR6tT1aQ92WgQTlt1MQDZQb9aSivxmPWqxhHp0Tu3MfkS6A1IafiBMDQl2nR
0MB8lfPbJJ3AaxEusWHqBQkvTQ5khrmxwlMSZfdONW5iuNhg62gDp2/JDjHb
i8IWCIDkI9wlev+Nfu7PpCfErX/MLiZ7aOcoKcJG+yNIPDfPO4fm0AQP4SFG
FXmq2+tvXp0VWa5Kjm2F0ovdLx7S/Qg+hNnYW8mg++KtDm64N6krvpaKE1c1
TvWlK/ZRJzGmI65XkXEXVT88Hgj1dhlVJk28KhkURN3PqvlMnumFPrrIFIGt
mMvl3ihHm04eXHRHME6dFQMvLSfHwHk4o+zgVHEU1ir0FZTDh0Y+ZH1mLGPj
umJC57VqX7/07G7rcvjzl4kcOJUgk4LnZhcqdBZqZVUuvhkvqNouXnz+mSs5
Kkg4AajJ8BtT0igwIyFI821l6ijrAzPuF5GfFN+uBMaj9WTw4ES03mz1q4v1
ODdndUkRl2RVzR0Yy6R5WUJgL8WeSPrwJ/tCbM1RbJshy2+AHhGqw47S7NqI
VlfbqUffLiSHKv6PH5yo7On+iQbgdn2B7/0umW+jPfWx5vKXd4RgKOg/rRRT
7EPMfUSAvU/FgJ2lsTiKYD9PvbgP7G1Br0C9zKBnSOPc9eLulvl3nlMGlPTD
UcdWkZpbAmKroqDkptzwZF9BRz3guI1otl12jbDH77prTSeusLNSwdMm586u
JwbiUrNajJTGcz5tR2EDfgqGHSW75nZ7vlnp4Tt2V5ldmznKN8C4ZQvBNiPo
H9emQgKNy1TTiBAi3CLWzjCZDhywLTJ2wh/aI5H5VOQfEG8zyJS5VVsifrUd
+wpMKNmUvJtldKjQWdEvHbiPl6EPMP0g8nGLNJgSx2fmue8JBPPxBCNird+p
Gy4I3ikBiMwwUx93imCwuFSSYxZytL81ARXEMIhCIpD7e1/Y6kbgfA2sgRFQ
fksd8/bm6Evpu8Wg8cm129UaN4uKJJhHEcgH8Vx1eXDZQxQC9MDcjLcAwA/N
izv+TUrGymGu/NSM91vZyaQo5wZGclEPNN0dBSGx2CDNVkNlvUS/jCebM/hh
tpymEMxIz5uNpXBrDqN4Vp7uxzGyY21uEVczc5/O7ATVI3CePC5L584n06pF
tkVJ3Bkz02525Ef3dCCECFPuyuSbmCYAhfQoI6Xp6Mzj5c1FzM1a7vRQtHKA
aOg/I7A1iG1I8Hh/lCw5aUjyIXwPlqH3/mKVdWMJPCSujHPyXK1z+j9B2UHM
/o2u+zLVXrfpIe10MGZwm1NOt88dQbhMJhQ3jiDegoWgPdRGSObyKk5gOTTi
gh5BVzy1e1+kf6mNDY67X3zjFbnA01JnfXrpQRoEEZpfF3N14SqYH1F9PtUE
38vkcfd0XmaGU5t4Q2P7XCjPyoEbO8ef9qPYmRIxdkAX8WPW0BGDTKkVdoA5
6vA/6FQJ8uHvnoYxcY3Fk2kzoqKcNJAa8DkZnuthpmqT6nMIaA/XxJAW3gkG
6upgDW3fax8MFLG+c3dK5Na40TJsLTOy2+KVX3emIvj0KVqFvASQ0btryx5P
RcBLx6xHl7eWRodx93S7MnB2vkNQZFQu3v/X6wKFsqW44BsUzlKPMl4LeIPB
B97298sNVT4avPFvBJc5HculCfECH2CBqFbRfaAxrVCZabmTgQGWChCdLOy6
w+YzZ4iYdPgc8RDGbDC89MxkD0Gx9d02fzFaHbBiI9Vy+9ZGdkfIH1Ejj0LU
fGsUYzp1Nnu9One7vQRB/E+boC/Noh9a53rIZwNpkXkLYPnUE3xlkRsV/LGa
s6IWd48JzO0oN04YF+IFIke9kig74uzobx8RXvsxeBnNdY9CpiB1YfuRgFko
LrQH/vSMIr/EDB2BUeEyQoQyj/w8eD6ZFI17UYYVfm8RFV6JW+FufaBfPYkX
xSG6H0oVMoqfiWjMISRQ4PfBqqOas41IQHWgzxF4tLkJN5XYJMeaX81a6gcr
SXzY+w6Ejrhb+7sHV1/q08UFRkiKsaqMH/u2+kNySqLAZbWKL0TOXKIVDvqH
efVMWeUKhzFRT0eQvEBs2OIVJU+VVPvHRJbXB8YBSYwXHyKpgVfOwk9sBwjX
FWKD5wReV+QGpmeiqbHoOp2UztF+c8/2g0aLReIw/WBqJ82y/HIVmgl8TmwE
3KFvS7y6zApGH3d9TIoRDgxrSbpvvO6Pa4mXWWRlzK+95s/H6gAWYEHeXSHw
BJtG720tQXd9AW8/wZP1HMjJci+frYA9hZ54NUxVY74WJOleQI8h3s1A/Yoq
JsUGGftSeXRDS6+0/RVp0T7fWevCkEYw4OO/ONZWXbpgcFTjSwgw0MX8IwHX
dv0PwZ1VDjGSiXpZRe5BCxckXwqh6M4rxcYmTcywbNIOJSRV3gR6kccssMNh
ikgdQQVMsi+mRr20y3j8S5BYbUK37KeT7Ab2xutprIZ8yWcqDIqB5v69SfGu
4S5GMJAAs3LPLGeDN1iyGVfh4N1vKIN+2zhvZrXjK3OBxH+xB9uQMLAzypVm
8dWeToA99BSTYLQVvlikyo9lqO0hh7cwXmvvUU+41GSHA2cfe4Hy3KNowhYc
VrhzrYmPn9qhiDg6abSi+ojCgBWBZHSU3pFm3cLjxvnYxv4r9dJN5M1FT/1g
DYEUuMV6S4b7MJX1zhNq0iwGWP9KzeR61TI44aSMVNpLND9urrR/4WOMPvFT
IU2O4Nz8lkY4x5w0ATA+WLm4IqEsl0MqI+ETVoU6hdyOuv0oMjfkY8p92FOa
Sdn92jFNtSEbsp8knJ5d0vJSc6byvJabNBcz+t7/0xt/+HCs8W5qdTiyT3/F
GRoahxfjltkh41SB0BIZfpC9GTL+yseFQUWvN4epnuSpY2+cUfr0DfVZCv9y
jBaD8JfDPmEgImfNYs626QWZGpIR6rL/7s/0tMUCXIcSSIx5A/tEQoPDmBJ6
MESOOwy6HAxkTWC0hgTqdfFV3HrCD4J6XzrWOm/jAjC8JiY0yVy7i4ycG7GG
GMsdYoZ/tThgGOkmo6cLBUJg9/Szcjn+oXe8H5AnRrSQXdSsvY0pZjFGgC0P
dkUHIQkLOX1Yua8vmW67PlPqQVTORxTX8evUEUswK+pqRfvA7frLkOnI2Bji
cOVsRaeziU8oDdvjOZeKU3wivElikRB9QDnOauewACQyanHldxMuIh8KnpKl
aqytMi7V/45bEmKSxbctevTeHhkybd/hMON1N5SdPelCcxDh1L19SsKqGej1
tn1h0hXADg2bP2g28aLD/Oh2W1P45njmiQdEJU/sRaKMWFa8yAAmsuZJcLo6
8Iok07oQUUQ+rps3H3TNTikuZASNKHuaqM6jwMYZ2L9Wm5LDM1ly+X2JoFs4
Hp2VZ7eH+Z4h8vtXBJLPt6hMg8AC7Z9rNYuKe9luoIcVaFy/Z2q2hbC1fCE7
F26gjaZqU2CpqbJuN7F4JYBNg7E+5MH7lWz309ZSANqEID//fczGsg1sqOxZ
tZeaPEUrKDgwadskTyJcy2czhS4Gy4YlKo6P6HnOyu3VqDqPlGjwHnv0tg0Y
RrUtAogUnOiuDVdSvnHZsPJnpvdMYuW6+uGTf5RjWo8wMXSK+fzxnAsru6fS
5Ib5W8JyRUTVHc6mT6G+nfqyVHFtSYH/0S25E1KXqeMA34mWG8F5qnhnpCDl
gs1h5wXq466lEyt3315Upb7dIkV3Qzhhu49CbVroGqCVRvJ5/a3zoovKjuL6
2rsgYK2EwITa8dNkUr9aOjCQH5XgHOj+bs/ehdho+dq5Z0uXCOKhaNOj1JsB
KvyQ5Uslc3LxyDx4hscfqBn1sRMvnTUeTICb7zAH7AxOF1dpxgxovYpVg7Dv
znP/7fDnejAXxspT+0WzUeKM0M1GOS8xU/feEZwp1/DxkjxslZopExKU/lPV
Vo/ofGAFtXKr+VAwvb+NnKdJTHKO8T05tszDWad7hc034JnGCLv3WaTf8U6V
BwoWw8JqZViOZHjoQwaGWbdwscMzrCiE3G57nWfCsOMNrI9bmhSNMBla5Ok7
BF7jHbzn8MlCG3JH/+8ht4bRnXty2rzOiSP/ex50GKtKnr4WbNFkgvD0n576
o2m1gjIMFzBpXGuhflbcL7Ep3fCWddLE4MsZBapaRwQ9/i7cJg3l9qP1BOI+
x1dU0zt0rzppaYUpjClvlBP3Hjn8lsHcqXoWvi6RwCZI6IF810zEGqe9a7kW
5fDeXeXHxnLQpvCsWNBjdlWbI6qV4VIRENsJjwMcwTaQj0m8vSDM/HKCMSNw
o6Di8lGN3IdqtVzIvBssNKX5j5AA676XLHjTp7hrrwuQkZPjt9s5c7T9Q/9z
S3Aj+003JOKjO4otZstJ7NLPrOIvB0qEw0PW8tStf8MkbKRGLaIEUVAgXnRL
/QbkbqJ2i2eJisKSQoSXYtwoy2iqPU9anRp+jn7UgFx54Twzld9baJr+6h4b
jN/d+WHAq5QpKVXZE3fDA7RUnOaJslOs706KGvLky1R/V7ZsYerUOB6CY/4T
7/71iKXtihdFoAPOnlE+5a/JsUidJW/h4dULZUSerOvLVoeOcq+U/UqaECiL
kJtkYPJFP1W4kfU55sEgGTcE1Dj3fyg1k4IY47FFMH9Hqct5IdJn3xBJAhA8
WT0BWWccxXUdK1iC5+NvFMkPNo/H4tPJo65uO9K1pX+2zBGvjxJ3MSWiXieI
mnyOAiSjOxJZE6h96Z9xXchB57kGvWIcfKN8x+T8QWWf0MHZyvjpt67ER8By
+kHEA6SMgvj8HIT86lR5r8IDkKtoX5gVR3ZskjhdyILqAeBT8KhcYvTIQlxS
rWW+Zmzq2vT3U6Kj0P1Pb+lKnkX1JPSMGg7y3sy7D+crMf/23si4N6RQ4DzN
JZ33DWyq67zM00/jMXtcX0tkyI15N6mqZRw4+urt3qzfTtcMTiHaXQ0FlL+5
s6ojWvH10H5ds3r84bvR7BO7GPmeQdargFpqJXmNPjV9WKBkAa4cbMuW/7Uj
ylWp/zbwez/+8Vi2CJDq/BlMjoSOA8XG0iMu6uQt8JKmOWuYddE17VcQ1vEd
HY5Owr2wdzQX1n+fgAtp74x4wfhHg9RD3lTtsofOgBYLfe/hIV1pc5gwydGE
FyAP1K7V7QZjvcMHdhpn4zJY3DX/wFKWOHy2NmaVxG2cHOfL9QHSJnDIHvkm
6AeD2TF9/8NGQuOqienS5WUZI/MvC28KNI+C8r7f4O6F5CWIn8Y8vCjjXX7h
4EhJWshO/kCOxzNmZ8ydr/EZLE4aVSALVtcdRyslTTcjfQID2fCmXYf9gghU
/NDWhmvfum6CqLuI/19lZ7+cCNRM5zxg28JEaDNj1ijKczUELLgFvkX1Nrei
TFpZ1hkCBXNYy0mGPom4yEk95pfKvflPtVoF06jN5zM0V/g47OTBWfjb3RsB
jhswuBfrP+HchOfppC/axKUwlp/EReb4Sv6oNNlfik9rN9yoSNkwnslB2t7o
qYvUK/8c4rDq4xhl/UCkClGasAXL3lBPIBvGQYDEn/IG6qPN15EmQx4nUR5d
nBnk624ZxMZ0bGvPjaw0Hz0uPL+28Ri7r7neGkipDBu67bzjev5aisz5ulQs
OcWiOfAubwhz+DrJH27QlXvoS2MTG660e/cb6qACWI2DOXn6FuK/HxUcJLnz
VBdxTA8JNSjASgtXa1ln6h5hO/zl7eo4f62kWgLb7sHPltdcVBJ19s6J6AN2
v/bh7cVOPkkjvt7+MFxZv118NNvccBxQ+HPaIsLv4G/qV6lObiFIsFpBcKBy
kPJH62wdbkiFhTf8a/hXHi6zjwqOeSfVxLo0wa5n9zWhhtJeDgrBcvNBlbqT
PrLiBolXZVPlt90xs7tHWD95ouHUdYTO2jOBlNqjfBB9HiGWVVrXsZs9J5yq
31qK0y7FkslKlDS1f1etK+2/cMTtT2rQHJo/Zw8NzCx+/HC7huVdhGi/yo24
JRGh+pz2Nj7i4X4Vp3SaqV/QMnrRcIeLXDMG1aKqXV6EAZ9GzKnLPGetZzOd
925nHOmD8tOCyxlzYbwPQRirjWHa5X2OESii+35cpCfjJ4azMqnk2T42im1e
LR8jO17J1OdnXaUfXNW5m6p+ZJEzOIjfzLoPA//k8HF0cc+V8kl6AK4Y6OpQ
qKvbc4qm5wtLRwyrl0vwdy66mKz+93O60e25bRDr1rgTGF1i9YbLZDb3ACQs
6uuRdPiSw9HDTChOfYJDCaXTRmz+mGbVTZJl3/1sN5zxDIHmAQ2ft678IKsn
g4Jy11f2VWd/AtwyXXfZTPfpoe6Kcgr1x747owTbJWVtJSIuw0zIRSZ/Aw7W
CrI446oJhdlPS7UMSZk9IC89/3RbxMc9QalDgy0IgTJyJ+e16B73UcWSIWX7
QdZzGm8ohOTkc9dZg1reMGO0M/9ErLOy2RAIDaNtxtWk4MSHiKaOdKnevppl
iBIxfxVGn7NVSubBpvgTbzOLL7s5xet+RqNrqRewsFaNFwF4mUetMl2kCH2a
yzpJLctmUY0XL5X+b1g7lBHPznh8cyrODqHq9KvIUT4fbl+C8nIAJckZ1wSi
OMzq0vRY1DkLE4a6Q2viqoOkZvLwribUn+mB+ncsC+QywRUA6hCmmDRS71As
i+Cylr+rsDyZk3vRMjEsQdlvNQXy+q69FULkab1SY9FdjsOTxLmPOqrfmo9S
fuJ0II07eE5FRON8AjgVFvTSPAtqOR87SDUHMHL4ZmU9mvAIEr7fsbG0egWq
1otWS7n3j3zlkjsiZVHIbviNVeCUH5NkF19Vrwun3fve4oKpxOvQ0iFfVIsP
whVtjlvIGJqUowgpsg3X4Z6rsdFrWW0MixWJQ2fmLTT5mV/3n/BbCWCj/bIR
IbDnUzLZUIPqKqOcTFP7vPLVvE0qqsKu1Nh648ot9mvkCEdm6GWnIiAbkZaC
uzjuI7dIuPb/gw0q+4GOW6VCAZ5yfaYuQmFBFnJlcrOUMe+5JSn0AmV9w9Cu
zaTS1YYTXMr2MwEnGrRSVSierN66pMlpdrvtIDGpSKB59k3U0YPlW9TOPAGH
UflSlwQlWyU4u3Lu6EmYtaZWqDG05D3eC4j4ymXVnFa+BJT/KRscII8FeMth
0CJcTi4G1mLeMey9hbdWM+FkECIf1Xnq5g49CzRScOFJaeAbS9JX0qnu4zMZ
ZVkD9pSkqFB1KittO1dnLKXQEP+20Jr6Nf6BSXbpvkOOZZPVlAtbU7AkCZ7/
M1ZZx3rPxLLlqIkcSwSics263Wa4Vge6jfAAA7FghXm36dhBDp9o9Wsu7+JO
LBhVNAcU3WB20f6V8SFbsf8KQWTFNVd6qu9yqriUHoQoU2L8yZpRKURzgAxV
1XfEsk/aSyfUWKdztpsXglgWsbZ7rh1gm7SxNGkkE4QIctn7Iez7OkhM1dO8
CkYPc+7Ov8AG0RBeywQNqc279lZbCi6idXGuoeBLmV/J7S5NheHJ1lJ827bh
Nzt/3WtIS2xNOr6VcbFl5osb/zuZUF4P8DwEGizYg5WDe6mfWPvOlYRUAkVp
NOqfkUMCxSUzhxeG7wEgCfGpLk/OeOnX2Krqxc/pHkB/44Mc29zb/m+1ybLM
VJup42SKCmFrL/+Skgi3Xt1pWuRyJT88CMI58SnUQdI0XhkuXnjWP9pKYr8k
AKs1F7efY/sWRxR54+jIzivvUUHAZJ6jAhepq9++F8CTWt+wNCa4d0GH8SA/
53rX40Nv0otDOXq3Dxgb8Y7bTtAMXkI6FPvcPEGW/c/KeXvHSCSgeYIG77Mz
KHLJiNaqhwctnQ0X+X6VxqwovT3cfbAfjdKNaI9FJlRzGBp3EutcDRwOipVK
km2Y8GH292fRJEhTf2bkhEL0O2KJZYXc/qMjvfUjVhVglKrxywq6Bhn0Ae4t
GhEJYpbE1TcYoDaloEemP1TBlnY7iasw5q/8bDW/LnCxGtg0QxE7X0QNNwaS
rDOpiUAyAF/7iFO1vflZxcXKj5Br/ZpJnmqnIuheUmhU08+j4b/Lt8xsVDLe
6J6VrQ9SnARfa24x4lCdKPZlTgV656CBjNajOGzMnMh/RuBJoFr8GKDjmR2E
y/zS1HZSWgeGxXjg9j/QiwO1fxNzft/1NiqqRqDbq1+gnePv5N5hKn20+LA9
BtBWCcYajRHjlbzXW4XJOsVj1gVYEpuxTrDa5Za/TYX/B/7nWf8s0/f49Uw+
rzmSI0H/0IjW0/kOwXrx+yuPKd1zK0ONS8VE8q9hNRmO34SVNXp2pC+w3EBv
Fi8fBHJ+FztvZrOkXsmv7Rm+90iRfGhZp2JzqTBPhKi2ui1XzoBc5fK1Zj4S
/v6ylH4Snz6EpH4uK4rsxYVRslORjkbpJTyUFk6ucwNyf/ffxIyLCdIBBfph
ZxwakUC/DZaFDUCHPfYcqevQ2YITEQ9SF2lkxLoAOox5it9U4whzhkRdktry
suYYvPZLr3OtazBv+23Vl6zA0Cuzcukh1HM8TPuYGpkaEnuPU4nRY+ZfeHnz
HMGSiSAHEByql6xt+pq6wtiCpQiBS6xs3qluwdouA/1w0/HM2+RIXeKrD6K4
t42WHUFKrCGCPM8dxghrWHcAaj49WUMl2ykJERR5hYCIMo++d6pnTAm6QwTE
ANovRgcddc3Bkhk4ghohBZPp+qaqV9kifoNzYKkxJAfbFnwAcTrEWtPizPhe
L/AskCNzewgLCPk/DxyiedbV2JYMCz9ZnYVXxaM41NYGYX0M9mMkVb3nQY7x
ixvspE043NzqRwkTHS2/WfgS//cl270TMOPGAnf2E7dg++QPcI48ehQddELl
6NeWvvFglPX3mPjkg4FyLm7GLwkMxNIB2pLDhIxr+ILUhbn9+7LpSINqGbIG
CFAzJ51z5aKOTMMRb/1aLIT8A6/EhyxA8CDapJBOhOS+3mkKCWdhDfBi3by2
gPnLg+4+UmrV3XzY7x84XXSLyylukyxgDMaBa8Zsy8lH0bcECxo4JC1360OZ
ufB76H4qxbVK483GChWe7uHBYiEu/ZqpFyRcr1hcA+SgJG2Tmphf0tx9Bxce
/DOyOS98nHxx0QgrKH7Io2cGzAgSubZeDZlwfpltszdQmA96n5ydV2DijPr3
jbADgLl6xhnL8MxtHXpTab2i9TPBXlEkqeQPX+rOEFM8HDbmpQ9GDCQSkput
6GteC1QOK1F2lDCG0ct669biKy1ThQ4crKG1D93OIQ96dkkHO4tIoCswtvdc
VGdH+kaBQwOSV6WKC4fFKQO+ezGW2w83SethRQMjuggDdgbNRSWgHVlUBFW/
60ZaKZW29uq3DKHwbZIORTjY6apLy5qGafTLRtMetT0jlmBdvun/iFx1w5Ut
ZQRLeei3TfDL2VEfViCsSIgkO8i1OMw+q00qFJVNbthL37bmXVyBU8c0dphW
DIpvVSPOBJfTTpXe8xAYqTlTOotcG5QcwHtKAD/nyQ7Xk+DFcyC4OMh9Xl/G
tTTyRJrWM2Ufb/RUfP4CfgV5Lz8K4UGnQgRl3ARHpSomBoea90H7wLe2jdVB
Oo3BsYO8HsqOnfX9iWrwUFNh6zkptscznS95xvbT2b44nN7TvDy9gUAwHBCa
XQvOpA1Vm0VuPal+00ZFqxAAweoxPUVMP2ZSuKbM3eQK4AN26VQhqsn7prmN
Ee/b5ydRO9ozHJ1U9kwbQxNs/P4z26QC0QKhpZh1psNFfBm3reEOUfF/sIuy
zDMGKyqqR4ct82yCoj54tPIlAAieY/2qoGF9puTtLfOQ3vI+ohJwvj2pv2qX
qerh4LvSxrk98ZH2RDQy0ZVxSxN4l+dLoE3RmJjNL1gfxPZeK6QRUlmE80mv
FTjEVN2oUN+ZBKGmQvYwHZgfKcTaZFGFhy4CT9Ihvqu6a8fwlozFtr9En6d4
BXzQMUHRLZ1cB8Z4m8bHnZWsDz89blf9Gr7iM06IVoZv4tepMytOLS9SOgwd
SJAjAboAx7digmXUaFfItOJw8WLiLIQiujT6pbX5cIfxZ/SOtP0peE4eq3fs
IgTilxvlWgneTIBGJjVfgc40i8UssPXxdvvcKVuIch8T3JsTWa/vDPN7S/Wy
ziTVxRlL3Zrz1k0zzsm2XpLpOJJWAMqYXlo8g1a6O8PFjRgNADWOv/7v2FUh
JudAmj5fEzzr9c7ShqD3HrBC6JlxB0HsNynL1y5tWM+cwYP7FU81EJ7dQKBS
6GultAxQZGweIFxR7pnWtEh0BHhq4GVPL1inTSe3a/FrzSemXCdNK2cxzBtf
zk2EUi5LZN83EYHhHnSb2DdnR/snVvIjvg43dYz/p9biRqAcxcGaQvVpPGqU
8O7E3TOg0yIz+4UtpZw4V98MHDOXJGRyCRwcCBoQMXZGpxS1g1C+/svuZJH5
UrsfY2V847/gq3QgW6xc4wun5olpLf5vOb78o34EWXA04iEyZeBG+gRu3BmC
/wJeTPjrajandYqWclVp3emW/MzvRx3c9kKfxnGWv7yYycZXj2IsPyJAztka
uMN44MP7rjNtVrINQfCv8Rq3DL6N+AMENzoG4cpG5LCNSrLn7SA0Hr6pYHp5
1fzmlI2dWP7Th13wMBLLknTJHajvdY2fBevtUw/Hzq5M86WKG6kRapxtcOSb
8GfkvjwvZhddDyvCIyYgKSjx4yz4oXlKUycx8eHRjVe+4FlH3GBoQ0VuvpyX
V1+sSxE9ulmX3U3sVDQhTYBpI1yNOlC0Wlu1MNjSABqycX9zZsUPWGbuVAZI
/EzYKbrQIu5m7Z5t60z1wRYZX00ZQMkj1WjhaMdp2z7SoUl8UghB0AWYH3L5
nbjwHHjvSQyHNPdtS753BTnfnhNnR79kcYq/M0BxZSCRxuLNb2CvLmi/nBe2
bA9ncAa1oGV6dd49eyyIl0iUobb2IipboMBkYXakTfNyCUAt2HIrR7dm+8zq
im/Es0MfKY3wI/+chvLYDv8RFogwqYG5UMSF/m1aV+Zgr/WwIL2oOGx57cyx
DRWb0ec27Og/EFGUv902c8+NvS20QYw+ikFEff03uFPFpvdUc3owiS5pLw2l
cpaky8VfT3t1ziIE1AFgRzo+7LwURPnGgoLuzLNFEm1xjAS2Vn0Jtcowfj4l
z+7fdXqS6Aro/+BtaqGDz98V+kQ30dz3Od84rThL2gVddnGmt9uR+uX7bC8f
raIJ/TwKs8eNHqJKB2s2JFuDMwMNVWjDzyGpsuPG1UCcK6grG+x8xDSd3b86
XIIQuGQfLqD0YY/wZlZo4nujoW3Rdx9pRdD2exkX6B8uId0995f86aq0bdoO
vsaC8AuMBpEH+vDrEbwV0/mlZ0IZaj3sg0JSvAwj/teU9Ux6W/VZKIpvNQge
5esbroWy8e/iHgGUIjEoDrGS2HTWHKceJirXWRg4t6fAAMlHwoysyDfn/5Cb
aCilfIuQZaA1nLrz9dQ4SbHE6E6J9fWo6wIIiWNcqsO/blfhvI4cXR9znyaM
7uEa+ox8cXPbZpHaUwsa4J7M2rKYXdIbCxCYHRuhFR5qSTKASRJTGD6YS1/P
F9PegbYcpXOBCcbSkpHLUi7mFSGvSl9tiBrb8tssflKQXX4iGe0mxd3cFsYM
c6YB7StUFsaNbJFEx1x6uphznXgvzSuMAmAqtkw+LcVhSo/R9Q98sbr+4SK5
ukEwt48aP+qAFTlUDQPJGCQELZFkWT2tgA9/YADZAAJ1PxUYgZgxw9XG9jG+
VV5Kzi+YTXeJk0do14RXMw3ratIXsZRf8JzGEA4suhwCzz7GNBA0F0+b4ciI
Uf9VlgHSPhcu6eTh7vVNJxwsrIpILgkB/f0ZED6WBRYt+L7VDV2ZjWxvt5Jl
7Vilf/0Vx5xDMAYuByiEq71sycLZVokgaP8xp9XJo4no6ngFuptbwn7X2Wl/
Vs2tynxlB2fTP1EZp6Fhj25P66OmT11vi8qoU3j+ZLB7CdVAw3jwJUePqOs9
eIlu3MJezELpWh2fe5fCNYxIFXdgqXjM5b0OTQPdgD9Lk64m6upyp1+ZDPaW
pHVb0wfYeaAhQSgIIEaSKGtsSiJ9r4SToYg7mxHZfBLPCOaeeMZnT3ntZrxw
cpX8CxC34NHbPIH44g5rquF6JOSaz3zxk5Tq05SWjv4s0ZXv/OrrXK/gzsXO
KTnfGD/lDC7KsrWwwSat4ldKqQoba01UXHmwkL3sRs6wHhCw0ctLt1uKUv77
p0E3hF0HURR4z969ZreqDn37IvsN1Ne9hHXeuuWs5uggPH8TbU7PJq9A1GIT
u8kRIFcUmJuxxcgrxEnte192z3uJKnpqdeJ6xIZIJCVjVw5uea5u94dj+odx
suhg/HI/rqAVmHGbIprEfk7HajGMZGs6rgGGngkgL0jBWThpVccW8FoYi8Ce
zuIgzVL9qqOqMeDE4G2skri0RI2jAKlmoNJpU7N+Gpztd366IogbLLsW1dkL
RWn5JnMsN2xCllk71ytjsEmrZSpvYbAJbEOKnrGsqbWCmrbmlJ8iu1GZrJVo
zAT/J097yx6TXXcuhMgxT9VWP2mJhWDznwQ2ITRFKL1LISFER3UvjyLwDJn7
40Ey0uAdLyrlw/7ZdiBzOU9hi7IDcs/oFKMrJUHnDSRohmVWcKQpmlhrYpmP
S42PHZXYJVuAH00hHFH/d6qtPPphvWddTemC5JXh3c69b6fKwZ9uBh7D+dsi
vze9sGCWa552SVkt7+3a0iT2rM+X7oZPOfKyzoLoS3ch9turo/GTR8SYOAiP
f3qAVUIOy+UCpayxvYHrcWlGdz0wdzLxzHl74JBoIkEdm0vyjbufESA8WRbG
sxG+JGxKpz5zuEr+5UAkcind0LyZbfLrs59CSa5/QnDVMSqeDl4W38sMEK5W
k8juQVjztALBOoSb7jSBHn3ML6tJsiMlxGMlWMY320scH02O1JYJQgNb1g/c
CH6EBtg0ydZWufK6qutHHu1H4hXERYs8e7HeO3fQIpYo6DIFNYSJpLzHStlo
HyaMEXnSfgccY5VtW8U4n/er5y5pviMTXBKMczJSzQxRLOqMHQQar5OGs/Pe
6x08lIvBhRKp6z+18a6M+Bc3jNIUtPPnW+j4uCXvm3FFYD0VQUjyVkkIhIqC
d6Hdh3aKSBKAZ70Wel7DlCcm5QwY7w5FQX/csRm4TNoO1cXI+dYLaYabn+xG
MLb1qFn6sTMhjAinV432UEcJvHGBzAwsd6D+05gK/qtXNczhcRJ0XTaPZwJ5
J1cFeoOjagTGG+oQ8WK8ibkaMFsPJpJlvnFgXeTCC7p0IgY6YWZaziXBea6s
T5KvlowW8lf0RzfNzmVgXOdmsxFgZIisntM34i2NkMq9FTBLdJOFFpSFeMHr
XRB3rNG016t1oJ+ZxhT+WdH4UB6ME0Fti8ZXVNMaMcTGfeKiV3PiP/dMPXnN
nz+DOd6Bi1Ge7Rls02RWpc67/NtwEFAPuJP6R+AZxSMEVZ11sgaXiYE6XDOS
hAhfd1xAPQKwvgxNURwrvva09ARGkY0cA8Fe14Bw/9w6DlcL7OouFLHVl0PR
OkdEkQiQ48q29z3Q8sEk0jxzqjG44JS9jsdIdSkl5pjOkfV2uf/oJW4hByUC
Y2Tc/NyHCGFHQDQUBvH+kGe2Sca5SAzk+215Fa2kWXvM3zuQPH8xV3YKMtSU
/lGVweJRNQJCBdkBWN+PXYWiqyEilVy9G0CGstnI0ROIQ9KVJHunO2/7vEWc
Gq3eoKgASpdTj4+bMsIABEgQ0Xa0M1KrW0B5mJXIxy0wlIommr/9i391Vpgt
24o+DjbkgBNY5FUA3gn41qxTUcdMt/6TXlATRA5o1dnUVgXtLf+fHJsovmIT
37nrwTZqPeFzvmV/5pGucSZymUE2cCT1cp7zRX1EikxGQj82iPrPO5B/X7+H
rFHQJSJdjB1Eli5sBff4bMKzmfphY8qje6IJ9udPmPu/hxrcQic3N5w4+57D
VOQWI02VClur20tp/LIenLrzF/ibwNSkNFVV7r/umVdPMt2CP0FgiiCzstsd
7H9i24YeUVbyOw5y9A1316emf6KKdnEbFzuYAnfQSUutfDOg6krzP/v577UU
i9JTnCVuJhmJenv523+aHFXDWWttFuEnYUpNeehuKxmtpA6XVfO1a+HDRblI
R39RhpNekOLGMQ/nO9mLFGM1MweZ1XWX0MJSpxlkVlmmcuPKox/C8O81RCbf
R0BfGqJRCc5vcyt1Pt7swQYGA+e+zS5UyXiBTLeH0JpBu0kBGz1AUBSNDrce
Qz7EtUjrgFaZb433vXEXav7RKhleV1ZImIbZmpcmzeRJZSMPuf+Ax5RbdiKq
f3awJBmEwlQdem/TAYhywXOyAAvqVwTdLIRy7GFdD9YNz5+3ZDzKN3GeSgLZ
VLg1dcW/RxNCHpS8jTH6g6EPflL30seqJOQVP0w5CvHrTwvYaKLC3b8Lprbw
p3NoAB3x4/nDZ+uyJbOxnQ9Xgq9Aqh8hATIO5nsAM9itfDQPzRuwmBtx4by8
YUA5Mhp6YxdOBCpPAji1EKzZ+A/5yzJSCDDDjY8Vdcpth9Zsh8Z8XnZ1c7h1
9LGxfDRONoIp6Ykg56Kgp8B5yiFIajZTSgI7EwOmHGClYb7NghNCA2iIMl3n
77NXrDhiCbPUkImBi2+lNZFldZV+Rjyy1AGNRrnf7YxlS6DKe4l5eWhbO1G0
P34Unv5C6TInxsbhuUyGJG2YvO+c8qeZ0XIielMbG5Ycln8dRRMN64H757Z1
CU93Xyk/jbDvYyuNfN5SkWy0hg0iEZUIXFTcbx9jmVY5oDyoFIkSCuI+zSqn
CNyicLzsZlzDxJXH92sM10Ah5wtCIK0Q9gq2e5ie7WioWnidNr/LoeBf0D8+
5Be0QijhU4wcjbH0cnWLjxdsMmA/5smon8UrYTD+qcgqoEdSzKx0rnu6rfBR
wVV0qypxr6luYCRFUaiqp2hBR4injBNXbQv9IvyBlqLoImClNPFT0CE2Gw7E
B9j+MzRKp/tS1VZjU9KtRIB9Mjeu15BmDonJK2FkY8tWoJOTlJes2Yij7mli
P/cXXvJ4ltZwcNz8RB0vXoXp5+NadzIIKRLUmSsh5L93L0JUX7mGkkhQE+Ze
ZDjKsA5ygZ9kn3wL9iP5q0+v0jnqBfuF8MZPLGOZ9lY1Wil3z2+0mOJxUguh
/No9MKQMZVSTVHySIA3FkMDM2CpnZ7VTodPR4ap9s5ifZG6+Dnrlr5bi1I4U
WVr22cpaunWcijbISzY7CazFCl1xYHxeOiLGhZsgCBHNNtnS/0gcMFij55ng
7sWC9YP3fFahbuO54cpDPkEDT+FdvghR2ME5BgnDztuJ8R3wh9pSK5HQv4fd
MFzAvFM9MfuBMZVZ4LCeREkZDIHSaI3q0bmVgkBPcLO4iCCugR9r+x6NpO/y
iLbhP44umiFQDpWCgOvSezK8MqtRXMMzpObCLbnh3j92hLHIdToAKUpgy7oJ
5rLeVggFoMn9OslxWKnSatqi6f0sCb0eRGHdACwKE85PcYI1HaxTkbIZx7oe
b8XPupKjMRtSJLBENqwEaVArFHzlMp7xf30oMTkau5hBqZolnVh5mPWr+7Y0
J+IRB/8pZefcJ1g9OpUutQpMkHxEsIcNNhL4IzzxPq2cY9YNDmFf+wNlzFuN
mnMxReD8JhVrjKF3vckzMrgt+/nwUF2Io1XFy/ERyXXumwWsgZ1mCibIv8G0
aBVATWwhu0sfCARG9dxG3yZfz+skMcESaX0uogeqCo/5hDHbV/1IStc12GW5
ZpRIBv0bt8fnLomeb2n5JNEQ/mgaYtD37opPQ1U+7ycjDHZxXn6XlFCC73/M
AWlyWM3wMFok8UztBnW7IMo6XUCG3DUYZ8ql7jB3Y4nEZkprdV6fbKmSF/UX
UBUN852RUteWE3pCiFlcc5B4OAAYMTtvE6t9k3SvlYHXHlWMiVPODzMpNG0S
fskGTrWBjJYgk+RFDT4d9C36+vdwPfsPl8nBK5WtoTRwkCNZU3qihGytfdXJ
hL4tiSwrvg0BDHF5BRo9cA3Mpz4vmUZbR+XJRRP+DuZLiclU1mDajJ8M3NuN
Xzg8J0HAe6AVgBcamq63+hUP5stYwoeR1Wfm8hII4U3nJLWmctxTHHzd+wjV
2qfrp9RIGOEp07SHTObh8TNBJ6TsDg5Y7ZRiXEMkL9uTaLyE+CgarhbXjQKm
HwCbghWyDUyHw/RlFfxhrCISJpOL+HgT5hNl+cH6efoomAWeO3laWu8X+l19
gWteWxBxv+hOP4YCIEf9/MCmUmblpTiyJGN/8NyYkO6UKDfT5cKr6g5ebKrw
V1ZKtRGfNbbl7r4A/2oypFb6/zGakDQjRNv6OOIJL+H0qbLfk4pSMmCiYIss
2E7uT2uuw5ZFjwvWIW0bLHpAKvsmF8/I2MI/iKg7EM80BdGFU0NvmGIsZzXU
J9OyMNvRu7RUhIoS5dRTXNYvparjUh4dZnH7rRDQWugd6ziOzxwOKzP2L0vM
roDnxiHEcOY6rF5G2MPQiefAzLMHPn4JIo2Sm6MulX7QKkkUHPzn1BYyVdMs
kgcIdfE57AfVPu5CaiwKAxcIQSr4BCBRfbaV8Rjb2RtJiclpTaRj1Z3PAWcO
lNW9J4+aVajnHtbuoMN0b5rFNKd1jFT65d3Dw2B4PUCNFFg2V5TYfwDlGJs5
biMdviH1OrbHpxKHBHGPtmasBK8O3xumy9O9/fKQBYvlXncwxf+uGoXAO3Nr
NbrfQ+3lC1CY4QfLnkbefgcG+uSSTtXagXMR+MoWcC29f48wPSylL1P6HECw
Q53dRypq2aKLU2sv21fBwL2R1rR3RbG9IHn8spXHL/5FbNlwInHYWxG88pXp
CCNDZJb2QSnMBINYcLz+QXE+3xMvi+HL7yaGqvwdkEg95zHQLAyqOckd12yL
kXQArVNcs4bLN17JuVJyTnmSgROBn6EROxXIaOayXJOrVmK+2bcP9G3fKPEB
WCcALGAECYhKOMeBcxICV5MCz3FFELxpMzaARDWm1RJ5aMuPQYu/TaIpA4a4
eyeuNtF06bHvoLGda6U6OyriYIsuKqoDcrsmqMex8RUzJ/PTPtylhKNzNM+Z
jA3u857JvRds/bv4595Y41cfnpYpRB2HYs+HnNWx0F/Q5YPEesy+mAFwmaqq
nH3YvydnUMvfo026sIsxbKfS6pUyyebR17rRsYwo1hTbBpBa24BhhTsoo7i/
ea+FrLBLRFzMP/YG0OiPJMmY66+6LWAJDWmxXEah9FYi6iOZGao/3cgsES5Y
rHdqAvZCFnmiphS7pdd6AjZQvEO5bOR78QiJiaoh+FrzLr6G0HGMNwUiVvje
bhD+dTZ6cr/KszrAokx+CzeZk3oX+N5niC4AQRyar1t/Hcy/JmCURS6vbrPO
zo39UmKO//o6Y+OkZJ+GqJPwa2UYZ11Gh/U3m2ayJg8YJJYarIP9xeqIeFgf
yJTticetL3Qa4NGpt6ab0gAx8L3ctIY45mKpV1AGH08Qvl0pUaQdTmIquvAL
JtVu3PnrXGpgMXolbXwV559cLY/rnI7fzE95S4F0IUsZmZ52F9sr/ycrStSD
skjAMyHg01VwCNiSK5sd9RDoJ4uhi174LIra+uaul2HfFvIGQ0ojQpB3L2AV
bOfldrQOs8pyS1/lQJf/DZdUHYM8x+TSwtMClSiyixzDPHvSQ9qqCNpOwMUo
9Qf9mV9NHzx0zMB2IW46aR+/eyZ23QrEY6NL5i5Z1s3kIlx7ZBLdy0t6Z2XE
JEBwjssCz9x8QleaAPtx2sRwySeymUgOIWWUK//7Z3P+iEj6kslDwUvzSctH
+7I92CnHik2TOvrT6BPDZMnDhGxaScEgL1l0suwtvouuy7of246GLp3/CrWK
VRjZAczNNzEXbxy9O/lYDjzo4c+b0OAMD8AFL/3epNBbYrp03vVSClKlZPGL
ZsxFqVjMYukb9tAXgLXkUcE18Z0hNgkMSxteU37Q8U/+SJAL0TQoi9tGMuVJ
DSBm1AarLRUOqb/2E5FjG4dd5QqOzhUq74A0DGvKS8b+EGwK+fq2cMk6mhNX
wTCJDRvxBgSDSuIjdTPPZ2GgDtg4luyNEdizmwFySbZFXxbDl+RC887PUSEF
ACYGpiKn/ixIIJzIV+aoWN+UMnFFn1bcyr+WfvwOpC4Y5+dULNL64zcFlu2g
D0+R84zzB5duhyxf6of6rCk6z2sab+PXchFmSllCRFfV/m/D95cYnfuYDoWs
Ttnl6tMdMA8dQB7tWBHJqMGzvaBqsDkdQPNeNExcUS0OA6ZGvGVi+DU76YGz
zC48NfnNXb+a7I1FB5nbcdJ2kq7Yg4Xrlb/nRNEK4z3TxXVTDIEN2N/y7ah1
WPP3eP/8Kr27vXFW0RUDYshclbj7L2aLUvd7J+RGCg76xtND6fPF54l9yWcc
ygBJ4JnlIuQWaBpygpgIpvFwMHIymmF2Itejc/qU7TOcCRfpmDYXvjTES9v3
goFptYb2K6NDw2zGI45AGdzCejtMeIPUqmLK5b2fuuIWC+KSXr95AgFmr5gm
4noWS1I+1xeT3qplu2+k7J5zcV4g4EsiAys69TBjHSP3uZFWxZQygiwnjbub
6abowt7CNAHBRxLnHrNfsjFuY71cTvstuCRo4fEen03eh0F1ND5h+i7cf/Zt
WG6Mt2A78ll2a6GaXXuuE4QmGpaDxMDu1glyN6Z+wKkInkGl/REZvRvxLn8/
1IlKMJZFoIxh39d6w53ZuN4hgNctf2l1CzJtlJYhrv1xpHOy/mr/eKUn5M9A
yKzGKEa8IpjFTeYEte1WmhTlgFCVM2nPPzF5yT9ImlOnZfORmENtSoLlxdnk
VBJgjLi7/0Abvu9p1YuwiTQfj22behnXQ2GmraimM/xjRUh/DjekAB3+apxj
FoSmhrBB+ZQc9nQJgEDzdKulYLMgI2UgEsec36nzJS3/Cro0aMeHR27fqqRT
Zmsoj1rpZoLFwB49wXn+F7+P0nwtdJ8oHjIqBBjg9FtQa/9OI+uoaX3vw4tB
T7NX/V95qeXbi4upRZZ6AgjPpUcvtevQGUk+NNKbfCuKFROwnmRmgM3btPG1
eZb+BkxQ5IU/tn2dbjfuMXEwkPXicwbtjQ/FFvJFME85ku7rubAHS4rt25dL
ikQpO2K6dPi8vFSsUOYvf0dAEpBnlSkgr3Rp+oLSxa16MCNAh7BkSdyXtNWf
YR2pKi4txTA3hzfifrbv37ACZ7YPZbaTV7jseiJpxY6TbVJ6UWpJ1vNK8tLW
L5gu0XUUuId4V5NVXSpL1HH7xw+8I9gXrPlCkW2SOSip2kAXGztq25lz6uUe
336NooW3kV4aKyExJMlAK4E+2i193ZPJbRuUxcttS3mer4p6Ya+3aZjF8vhj
Af3mqBPeT7lAK9dYva9YL/xnloXWm3RV9RPsnpuip13uqhHkhWQHCc09Mn7h
Q8tUGbWZABYggx1k4ZlZHcB7Ty8kxYKKN3vmuePrJlu2+eUY1uZL3OmK4zb0
bPkttYLDZYlgOBc/zI6ll0OKAIXHATJaNjn5owAXCyL8IHE4wwrIKc4V51pz
EyodGKTqx1EWOCZI51/emkFKjt1vN6QMRHOyxRSdM/kVqpV3AXMIpH2aRB5u
TddzyKAoox+v9gGpPZsMNHEMV8amHbykXrU1yD9ZoBRiPsQb02lg4/YGimg2
QWeYYZPnSczjgZHVHlEnj/IuWnN9nTCKWfxrTGXBmHe3B9VKEBkMeJgdrmbi
OCucyFkHUvC0+CjSHKy4BK+WlQv97XjlaMNx1LBIwJ5f967qodR2uDMhalOJ
fZopYPD7KSRae29IrMnIFMFppRW+078y/+UBkrZY02hoytbb+xFmIpTRy5aI
G6KFQDzekG+OLJG4nlgljEW89lYzQEt175MfTVmoB9czfAEiqmo9qpeIeKP8
xaJhEvYbbMAp2mNAnU78INUlQOg5jCCAH5RAuxNa1gpggpEw0aKMCFcPac9F
UwCYwcZcvNKGzxK3aS2U/k7ky06ye6GfNWjy12JjUADZeYMjZeiFBQ+AuEdE
rIUaOGu1BIaYa8M077qMisd2yterrWQOo9/LeQdGXSQ9dA6sUtnj60JAJBhh
lgzFXph4ZBW1lhCwtfuQDsrX/1x4lFLwHYjfE9iPgULOGIp/+l0QMhUmbKjV
YAV6sZJeqFDE6Y9uxc6kM3cxZEm07m05TUFaiShGO0ooG7a/l5lWpuZsbnZO
VQyJOCqnXKTAZMD8kg6pR4sF2J/GAES2UenPkn6woIhjwq4EPxSo97PR8V9g
9EdOygj6AZgvLhYa2JPzrumwRTJWT4yaVTKlunh6QedBUQXZAcVzNF4aogUJ
zGP2UVmTAMVEAg99lGqLy/0228cl7rXzMD/KKG0vrRvXBQXc+qLdyPj/fDkR
CotfaYkkviMPMIbmAf/dhPLHalsshbWOfnH8DOOpkDqZNSQKcp4hEtdWteqY
SbfQborzFtMkjcNh1lYZXiCG7UGzOzuiQqe5rUpr5elx4y550Q34kAcM+axf
z6h1wEp2e+nk6bvmFR5Q/tEnRPfmDnMyqPqf1tdq1rhDJhUOAHWdvLc49ydl
ZP+o/GGx1dxG9mxsnaRNQLnKr2bQsiXfku59SHeedTwugN/rxO376L5zhOCc
xX/Tu5owb5bb6ysdWD+K7amW5Oo5bnCDb40J172BpIqDxCO/pMFl3s075BBd
dhn9Np4PaF0IWe2KavThM/FgcFoU/ZjMs9QLaBF3Qj1dEXig+9al2TJ2AbvO
qn0eWRfQuXErmwVSN72VUo9H0dvq3uDcTmbBRkq0I7mloJ8MVJDNW6DzPWCT
lJ4ypKQ9AY4fAavqBsOgW6ng8hLgjrEiiK47ktKroTtCfHLMO7gKCA65RJOj
kS6KfMYhqqBq0XXli4lj2FTZuGwRyObXYtnr4lFvW6msoR24LMZu6fuJZGWa
h7BpxNG/WAjUuQfiK55YYh1xrBnBnG776C1YbHEOQ2kw6Huj6kV/HwPZK6jS
hGpVFWwnCcv7m20SBXM+C0PyqYcANrculI9L3AWSC5JZtDmswsrNQWCf6C+e
4FVKvYX3HIDsfVS6XOeDBgQ+SYSTny7Xz8MLb9i4CgxFgNLfLZaVeEyieUcb
S1NCxAEjzmnljxnWI03fq3e/QSSYvrUyH3az5wtoBfF0fRe6j9QgDruUXkdW
AiM/bslvQuFLS7nPkzkPFpKrODzMzke/OY6bu41Z6lUV/guD8neWC3l2xxq6
Gf/U3osUe2+cnVwP0Gg5qfwlIZVc9dQcsSbrYtdG3Mz3Oyfe3Arv8dS7HzAH
JxwACq/cy51tG4gTxDJa36T7xHDA9aN/jf2HY+thruXuu6vmRv94+h+v3iAs
ou+lQLbdpjan5BukpeQufdO84pmo2Uge1qS+L6qUNxsjnIXJg/3ZXor8MZIl
Mu8PCGoIQLxXgds+umsvHQ+JwZm6Kv4k+d5U++iD4yyYz6Ch2O3OCiF4zkDn
rGmL6V46WilPFacTrRsuKU0+7RFB9gYyV/gz48fjRSmSDGeBlZdK0xeV0Ult
CXlUilqEiA26nZ4F0L0yY9daJy4BfZW+775Uwxi9bB6t7vlpYujTiVWDX22E
fMTESIFzHx7gb2x1Bx/8rWoTJ4v9WWW71y9wVBvLPowQ1kx8x8O6N+X8CNvJ
xI5JuVcshXE520FJwSHY6D7ZsmAuZLuecCIGpLr13GOD0egoiHO66gGSpuBW
QhsYIJoBtSoZspbW9D2sjhD49tSp63H76wKbEFnS7FPF345VuHtpe6GIlPd/
dTRXRF8mJ3mRMpx7WE258titr+wcKcyBWFwuxMchDId8B7EVXpjGbZNb/lEF
+uAi18OWStOncZ7CDt98eKZHZO45dLKtBDoK+cwQIdUkycYguOFWsjywFdUL
YRHaswCFY9DY86GC/+jDPn8ejmEg8rIb6EXo0HIX+L/JP0SdFdP6JcqsklNb
JVrzp3MGgf7Vup/5T+KSFz/xppLPwM9hhK2VfVd5yNtLyhVzPKmcp8jTiP1i
ZMD41d4xpIoc2gCy1KjZr2gFllnFXgwzdmt2C+F3DpeyVubuK3NVELt5Hk4o
efuiVmpxXpDFhSSU+ivYSwA71tt4vhFkDVK2oAxRhbI7jySKy67/2r+lnVCV
19zqOf8AQFlQ5/WfgMxpJxhZZvgUC16uwYP2/P7iUFcTzQtg74DuOTow5gf3
Hs6Uf0IkhNMEhU5R1G27SN7MpWZZPD0xRJWUaU5+iMbpd7tMy0E6YxKbpnyT
oYvJg6ab84biD6aVq3gmXjY2E5yPyPjApCkDSMFjylyzmGhLNBOaQqaQNrN7
z1W7q/59yJ8atViKg7RuAUO9ex1TQu4GuC5mc73KMJakIyT86Xf7Fix+ffKk
g2L6asa/rdRdOe4yvimwRXxBZHWz9+40UIBVsy6yaM6iyN3tbj8iDpwUDzf3
MGRSHH3WMoULAHPssez+RS153vm3Qyunr2h4+MOZPzP+OXA80L/2UjJnd82C
inAKYY+iTrH2ez0cSEMFjAEOmCT9qUpl2ITMdtf19buxkADx8+YAZ1YiDDl/
4b3qPdUeCov0oM5J8ARhMBx1QA0kUr5opNf2UQ73QL55+ArqVXlofW8doCjj
Mm3oAr5nNpoJiWR/OeJwHxTL0GESD7hDCTS2hIIl8XJSbpb4VyxVe/Kd44Yf
IGxqPhMN5a+R8f6hK3dL52Zq4OLSWH3RUZIudl9YSp/q6Zi4plOzI5EGrHuI
IAix8mQbKEXai8Ok8CG8CbIO4ACVxohKfclZ2tCDi89U63+gEW/PuK6ac35p
l8ek10AJ615VVJljqrXreHI2rviJskGu1xnm48xPXHCkpJqu14m+QFfUeN7N
FN5NvQPQmF5FKL74ZFCNP/ALvzDLYOiQf5URtrVK16dXjx4Jh/zN0CG/yatI
C4KVnOvOmxZY6bsh6DDJ35I+y3rSGgIvppKL5vBghxIgB4V6xBMqaKZt5jCW
bMHmy1DK4KHVTpJzO+KKpXocXOnajWxN2klFoxsALgQGxH5mzOy7cY3Es+8P
LkIPQM0MnTVNwJFMQr9UW4vi1H9AX3t3DAn3Er0MjujO4GATlnxAQfMaxwck
rLzWeJ0XUnc6xPpKKNBcRpL2aIdEmxMh577nJ8AiWIAiqP6dA1Z9ssBzF/2S
xsthQpf182rPfsY4ls9NUESvzKmFxd/WkBZZrRFnjm7iLwqjt7tsVE7mcWM/
VMHy3zVslgfWpOoEHcEnN87BT434BhHzXO2Hif+LRYI2HOOSwGwmo95VmeEk
qev6GCu04cH8RqXi3T9sPG7lthAT/VQCASDtawUhTQKOpAH4CcvOSm99QcEA
ZO5Zqt64VBShiEVDoxEMxfNgRLScxLLcIwFbK2Z2MgemQsWTitw5Oo0DbB/T
1vmqvHawtnfKhK2C90u4QB/mzIkJQsNo6By0Y5v07SXgvKU/6+OPeUJ74aKN
9iS7Xr4CszI1A93ySpLorztPJRhnXV0T+xCX5UMwHWLsg3KtfnekIuyefbvf
ivNXPfLd7Ays74kPXy9lfEl5x4gwDtdNlynXpha8V3zewbxi+ow31HeSI87q
WL/n1yoN2B0TyZZOqTDvApDOczkPqa/Vh7GE6Jzt6Aq89rXN5TIwzQEKf2Wo
NFGXiSLHdjffMs19yKNUyhHDEcFjhPAnpswjdcMXX0uJuA12eGjv4Ks7F346
Smu9QXoTNMY/0B4VguIlfyrN/s/viY395eONOEC8k+N+qBzhncLseRz3F1V/
id1+VU79AC4BRWMc9HVUXtp7l/4rVVURzizhxUXrgIfyFUU54b6P2A0tdun1
W/df6vs1M5vRhCKX6+iKNLJd8OkXm2IEVqHg2AG8/GjDPEZBAwg02q9NZUNu
O48QWpBxn6ViVvpMKifatmu8FfVeaxwamFZVgk4/8EoSyhQcxQCvSTrlJ/wg
NS/TXWulFPKjG1MvoJF4sKxgsx0noDrLuRLNhivh74FwDetGubIoqaENZ7jh
qbclivDzYPA7yIYweIqyXTuZTj/1RxC/T7gGLT3NKPXgTwDilBo2+pKqncb1
PCsSBvxqShO+oh7615Y/fRsZl5btzeoO9YR9AuoCTYf+/iIWw0L3yKJgNnbC
BVYQBnDcTNsbb6N0YAJc87x93nmP9Y9vNLTrzSZ4bcdiHGHxFyBX/gRvIfiC
LcGH8r4aAU77ZVHXHUQETUlIzxMknJtJCVAQejmOMKlL6YOPdICl0j6wkoR8
i/iEXxuXSyHkwX7vo1Zj2PYlhAgxuMZebbT+PD/rCbl7I8ejqSFFt4jhNHGU
NziqvukQ4dVw/htLmjYWCpyZo491e6NXMPZVSFTIglBxFzhONz7UQXCnmri+
FvB2RF8znl7UxciNEakoyJQ2d15wjl0qD2EgVfhDo91Z2P9AZfYNagsU8W20
WjfCGJsegf2r7gxiL8F1wNcPQ9V4IyzAtT7Uef6rx2HP0K4nlmgUW6Yl8EyP
sLVOKrwE/dd2ZW6MmmVsc+hTJV9P4p+9NNUavobgMZJS9GbDkI45hyDP1OoJ
eHtuk8fetmzjOzfOHaNB/xHuMRSAnY3/4HSK6fHqcnJ0h16i45uY5rBqh3V9
t4sum6e/fkrDg8ZBn1XYXRKqWLTQmIO004/tvY028wGYc43En9ZbCoFHscgO
ERBB7qFIsR13OXSaoPwFSoJnd20CfOYrQAfvbRmCn3XFlx7kjRd8jJsgiddq
7dYLcyOdCN91a7FKUh2i1aRJ1mRt75/8VXNkG/pVc+1N3m6PNiPjk0sDXGXp
MXQO4Cdk65IbS3d/vsXp+TBz1nDPRtj6riE0an5pBjd+Ho2Goo6cn1GrIf1N
sS2KNmA0toBjzps52FlroPvWhkCB8/xtmjLHoBmh0f23TAla6Dp/xWBn1Qu6
OCazIWaA6JpBIByUiLANYBZ3fDHKrHwwiQLPnz2P9pifv+qO1mXmXRFaEuAA
evU3TSyF4J3pmi5uvINBm0FY3309XRfF9vLYiZZZpI6SmNB74hU+ADShQSnw
UBa9M1syV9TiNu2h7WeAcQ3KRo/jh4fsWeq6vIV6k516OqV0pDSbYoncMxx2
K/IaWxel7ftAX2FgD/T3GQy39jMx9m0MO83PqZet5jaMV0IoaWwDRRMDI/aJ
BY9RiiEUgPr7wBCqSfHnJLFBh40izgdlhad6qvp6IRgzC1hQ0wopj5j9+08U
TQfnL1dZ9IFYck+G26A2F6y+ObX/PMwW/hedzDaVX8VIt2MITqtwB17xO7Wh
lyFaHPQ131tD7hIy9V3m6xWeb6SJs8SYS52hJXnFgEjfM+jnlbZB+tHR2DYK
906cIxvXWveqinPaE80gyr9TZbdt3R2V8ZERzd08ezQnIpz/rplUoapjFQiY
EIMhQIiHj/ajsdg+sZ9uRsRZcbOnt+m15INDeGfPQgaCl+xK5SRzXu+Slxik
Sgqy4Kn7EDkUvvwMZsjXafHyzqG/vaXaUQD3X5vKNJEYhLqaf7+ms+mHdgll
9IAouNqy8+kVXu7euCEiOwf61k0DsEG/8k0ur8kxCKZgmJpzae7wjvzdNwOq
4el6iaBz0j5BU9Vx4xtBbHM6NI8+d5ne9rg7kzpDCX6N3df6bQe1BAwc952s
0e54QZ2OdPZjOTKxN/KT50HC8pNHfusYEz7P9uwYR6TT+bFUtJXMXk+bqUS2
Q0Jco1nRJqaYq8r83J8y33GXv3jp65b0X2t+nyQsNa7K1nrX5jGu7b017WIm
qqUz5ylnlKf1Wc72BoKAoxnVckzGuaKwzm/SSqzYe6H/FxoPYGW8knFk7g66
SiQAqLW9diznr6wPoSmWAjvlF1N/6WoimGdBNzJdVaAp+quUVoZ4BVS3JlpI
llLI8pqtgF9DUOCC0Br7q48fAImO6uI9jUELtpoOfuAwJfTsNL23Ya82/2I7
zmyBlEtoqdXuHxK/wlNCYVV9e7grYjOoIEIW0O2z07OF+TDWXxFjZyjQbzL7
QzXwKdFrmrpt/qVyO6QGy9VdkfCROEfYC2PSxhPztDjD7jhEXhpcQ7kmkTBS
gqlVBYmp7yrEkZAHKjlBahXCOje9gk7Sxu4eUU0tTKQSc5K3QE7l3gDPz36u
khIL5v4xgP/2o+kAdY0UwO55HOGx4scPdoPTQbZwg8tcc30YcZmT1x0lhp07
CcMIfO4lbwZqYbnORJ68+sP0gRiofba4Auiy0nS+3BLA827Dm4ohB31luGSp
Nj9j/5vXDjcMetkGp3QYHRc0AdutjvomG3ghBPMB0piqKZwuEK8a4O2He16h
4pjVkeERe0Klzujdw8bUC6AfQq2VDh0W2DoJeLZJpVrpwVMoleKBrcP88IvC
5IBwuTzyGo1+0dqkhvmFml/LjYZV3VvKEY1xOQ6qLBQG7rFFEFSO/BqWGbN3
GDOY7SlgnsSAr1ViP8wV+FjvuXs9Rwq1umb/1jJN9i65ie92ZVGXNcqcuEyb
Ajdr1HyPRW4E9CSXxAvY0/1FmmfS1+uChRsbeF8DBaFjvCeWOI6ykyjTg/ma
8y33SycreVWVDBWtatELXxqQnh4nHn59G5+TzeIN+7ezY08E8u6p1sZSQfRq
tNXeKWml+7rGB9xtwyZWEkFSyzmQ/+pRveCnH58/f9w/FNtiry9uD4367Bgf
JnV58qAe8E4LXdyEp5Ydh4cIVb6Tqxaf4ktKDvjuyRDeEReWa9CP77bLHnIX
dAO9HT9EvuPFUut30ghbD1cfaPXb42fK8Rqc7p/x/QgMp4ns61Nlbu36yj51
qm/SVzP7zC6B+yjHbqBghoANjBds751y3lfRJMtfPBp14soAgWra51T0Z7fC
WUBHPWT5HJHcTevakUyLIxuguGQqAZc1fY/RXBlc+exfg+bMUG3akNzco7k8
he+NDLQzzl+XfgaCh5aVuCi9Mjrt+G1z4DoZ6YQZtxx5L7gV3bzZkVDmcgfc
R7bxRNm100LSBrPljPruXD+QycTSyTx+KUJ84h+Iy1NQ1po8+uKZvCyc+8d7
PwzTJxkKObVVtrwO2+VSHYEguJujb/FsB5oVc4R2V+9BdDmF8c9Ch3rZT/rm
kRrHwmCkUi6bOJkpZdYxWFRw+2gPd3AGwoIXBdD3Qk1YerHCxoeCH+T4P2T+
+P/5e1gOmOvtJAiQiiyqpgDeWOSDYzeSpNylWFpRGhIL8dHzvvvPdbIflyFM
xg9KJhVyvRecVHf0Mpi40ov1/bem19oopfixwhnJURn2k5hHo6eEoubxsEp3
tXETzujkCuE/L6EISOY5KREfm/A8kxMzb1eM5Y2HDM6fJxKq7dcu2C2z9VMt
QZ7QOctekBIOae86SsmsAJMu0VE2f8p+EbxwBD9FU9eY+nbJ/OBpwMmFX45e
fHe6Zo+T2o+Q1akjomy1XrzvWjcya5e3Xadmw3ZC6kFqEIcJ4uij7PUYK3QY
zJfOrz3Y45Vjz35v4U6c6FTwNGm71BbyKhT4I3vB4chPzO8aeQCviqcdlJlr
yXk9n0cNcmpq1q4ts729g7Tzqfe5n6zYCaBOyKm703Q4Kxu9LdScai8yncn2
aF1CcKGx1sfKNvgMus/yfR1Jn7fTybcsLnJ1m0Ceap0XNsZCAlC4yRFCtvKo
cFQi2fU43UVcxMl/El84G4/anueYLRRQwndgLJjWg67BmNZuxh1L6JRLpPEO
v7713saxYLIFyiclEcHS5YTlo2+2qgRyxSuFhzWvmyCHEAsMiy9Im2oHyd8f
8XRNUtbysIV+zZ+zFyVJfhdSYHcB1OQBntQ2N9DFV8SQh88b5QM/dkHxWxql
xU71hA56X1niDdGwXM8zgL2VmFi7zoH2mGNrmANVxhz/Itgb7NsM/dP6Duox
3Y1AuxU3HzoVESJLCFdojD3WZYHDJS6Hsf/A4TDI/ajKKEd5we2C/nVHJNzC
X0l8+wKlptfMrUwwp6vQjRktO0WYwZXFujyTs7ikK4rG/vtIDoBoHsGW+Pg2
z8v2LKBD8/KdKH1AKAjjIgovOVl6zpKmy7EpIcxADZulDOKUo3qZBjLsShU9
T5pIgKXZ0/VQV14nyMZqvUGR1UwYFo4B+Lj0/sxDnLcUMhnUZQTpkvRmBESc
DPmukKVod7GLLvaSZHvHO9sPe03GZzOEQDY6Rx2KvoOCPLXJSgtq8uIPXNpL
e+EOfMoWJhgrgXG4wnOP5yuObeeW+i4yOcAEyJ6loyI0WJJbETsM9lT9Jvqp
d76QmAzUmAf5k7eFnQWsGXo+l9MT5I8a6+tmSNPp1dI8Ub4qYP/vYUXcHnls
GoLQWH3lxSTJfG/qzRQHpsVVtzf5sD4P8jGfLV/+9+DzZDR+nyafEQuOhkyL
ZcHPVgJgTtQtkqf9G47JcUQzyQ+bFPLmdQkrOXpzlKli9l7dmRb1J47NwXuw
9Kreyqf2FawDbdBBcNR/jOg7rJoOF9pQHz6XtCihx7KT5YU/QyfYGio6q2ER
QR2J9Ic1OzR9Tx92+1yo4PmaOW1ncGz5OSVBGE3xgRcx38IwaZCORdx0gSPr
UmIqAe0NuOl31UY7akYJrJT51GoIn9QsykjSdYEqtcsDVy/FrMyCGfDuG2L+
QwVjvSn75PY+4EX5MhOpesOgBKxghvg88q6CvbbMwz9bNy0qeihLsPmxRE0j
MToc6pjhB5PEKCwdfzyEnQU0dOWcYB5y8fC6hYtNSXUycOdPFJIJHyD0aUFj
wrXX5Kd7t33SP4CdjGUacMQHTs9oF/UxMXLtW4sJzJ2nJV9sBkAeO+AqFIiL
WkNYAnBx9qV8nzvzWbN/0ba55VVi9FK313D2XyR5gvTXqG8x3nwKMii/hXu6
HiFhtbaQPiRZRhOj4zE18kkYmDAcr2DsegnrAh2q9EqOtt2gFXfdXViIETse
U2YSGNhkdoGfBWVCZrw/oFWfSWUY9Z2ApMQ4AVNCBCUz20AbbW6BayTIxmuH
tCq5G57UAApAwAhvwIhwJfI8HkcUk4zEvaMt6hP3UkEzdX3r6igv4pQedmh5
tqCdy+y0N7GW3lzJs420ukVoPiNlr+ebowjTxtIYc5mGGvZ1Dl58USZlQoXz
YG4/mn5JpmGwX4jSfW5pEtzx6DJUTpz+Xv3Q0brmR2nbp+V908jow15TtH3j
Lr8jq4FrbZV24uyuPCSkVfk3+vi8dkH9JCP8yv0iwCszix0s1BCfcWB+npiX
i9IyR4TdCsKI4oxrkN+fYR7P0rRiHhdB9FsMKdGRaMnJB6u2KbJ9Ss4RMz+V
wh/YWBd4u0J3VZZmD5CCEWXmpz5bBMJz/r40nJ9s32KzCzQf55dKYfB82mqd
uTOnSmGUPk8jL8kwKxoG3VlXFipOsVX/GHvmHtVg++EmLvU32lP6NB3AYyWF
RuR1lYA1vV9uaGCHiFfF4p+vOw1YcPj/6eXUfmYXC3U4+A/Pd7GuSA9SUUND
uSQP5hwtHAAAx8+SZqSM3ANRlLAwGztyXrpc4xtKyGgLq3sl6xHlVLSfFmf6
L/lcAWBi/7k9z1yJPDagB+Ng/kQ/Y9KVaq41KZ9294PDnUEr5wRSsDfCg/U6
PSgyzQYBxleC2IZ74XSpH0InOUflF0qhjZ46NrynRgl28G4kjwRGMx7Ap9EA
RVBn9it28hKL2kw55ey3n6VrbH6QaHaZT4TyrLTpp9+XzF/CuMc3La/Dyy7S
VE51Rbmpg2ZorfcSpdyrqNxkjZauSLsvJdS2a8u1z9ZNCrFQXZ4dViVXlP3p
tE11GD/fMdf2zV7amVNNvsKtKcLBAfEe6YwZvnwcv4uagP5N2uVz7OV8UgYj
2VSI398r+ggm7yfkYsePlZsdwM5t+6Q96TGif0p+k7Jlonwr6ob9Km2fCKw/
It0MfPDUW6Q8nazSrmSkyOyWrer4QiQ0RZR7dA6ILRwP6yP0+2LmYPcmzqqD
Y3+kmYE8GFxixGOO40PfB+tQ2CLNQafyYdFFL1YP/rgyl22ng3r1bt3wOXGG
4LC52GwTf/pHX2EkomWiGxKqV6YWcC4wxR6uytMnRcpq8r2xJiiYG7DuuVNy
aOX8erHXqZWjg80e6hqBOKWfLg4EmbhrSOEHjIg/DqOG4KRBtOF55CBrJ2sI
e0Gjce5UAN70US/RLia50xMMqVZKEEVc8DjEtJvN2e9JeCn5ur0SVLxmOgq7
3KyIrSmnP4SVxieR6ezmIGYQZudp+TpjsaGlpNAkcqGKWyVl/BO5wOkvOc/q
5ddQF4t8XwAhJTrzZJmCzV+JmSRjEY/wVPij8WGPRuCubP8Wozn/dRb/PZ9r
WC1v0OSVr9qScWHSsR6xEzVFGfFPAza2GNxMtiD2HZpKMhsiPGMtWmD/45yT
WXG82CawHMfwD4I4j0qss5MOuIdSY371ETzjGjhinqIDi4OOxcuqLJSFSsFi
76Ba3G5ddvCz9ixOt9W9of5oTWxUOQGBmHzbTn5X4HoNjU9QpupArw5uPCg/
dqGqFOgoB+xA+TQhanUmHwd0xiruSS/zphNinxI+8l3N0bEEQ3qMCjdnPTb4
prYOW+tWmS4gVzpi/lRIV/gQ1XRrfHRptOrBQ9b2WXykvIJ9e6Uc9q+t+s/k
lCVX3wz4+767NLVuCfuzHnBAXpQm0abdM9nYtBcYt6LAWrD1ZYfnjcAuZ0PO
Jmu0pejO3sLPc/sxPc9fZMBcC5Sgw0ed36UV7BvYEpMZowNraF6XGe3tDck7
dIa4IbVhy9mAYw9Mf47aiIbc6+V9K3DlS6KToSRItd0lx6jz3TVW8lZNAB0F
2LLS9xqV2KniC2aWcITt+KdYympABKWpf8b4s4bW81WccqWAQajQsK14w2U8
XlduM1uXz0OGKjVrpEBt6kMGROiegYEnK1dE3A6E8i9UAVsJZd+iz/2HGSWG
RAyiU4QZkl6K5V1Wyq+Hq78DrEN7UFsZYTXtrkneRQl4TYXWwA+ixJIoPL+y
w2IbgpS6iDO9jZEmBcA22c+CetEooa1sSLNssZgPLEvMU1CU67nPzEM6/CwT
fPROToKIQ7QNrk0xq9hFsp/lwXRD6PEIjoO/kwUwZyLBVTGazKVLYMkfMZvx
wKC1W0Qrb7SIt7idpcHOx51JI/3b6CWifm0Vtna1kMpMA1v2ZAnj0hGGafcz
xwb3y1O5XWleIATPHUqCHlhMgDj671lEqzlrto2Ey+0sj32lZ0/j5swUrfkw
DW/wfFRkQh7uxShnRvovJHpmx1zt7DzcW/kXXkdv0haAjiQdkH2fENzeYami
RNr6SI65w6dbFgXgygDRGl+tgwCqUlRNxHot2QUQfBO96dc6mTU/RdAVIMf/
xDUK6WQv9creUbeVlDY0Du2T83qwue33nr1585FnU2N3cVpfFodk3BHP225r
YQL1Ffgna4E1YY9FmppzBUNeqUVHY7DIRlpbPOS55krnfDQAA05VKfPm8eQX
/geVdPokeZURHkWqct+5NIwRQWXePrHZxFCor85s6rg5DrdFWE1vDmpnJvTy
qigKkFyqGlrfZHyUew1Q98sN4B4+K/1BpSUOmkIQfbcAqUjN6VcdgC5Wj/cV
eIBxrtmGqJVNAvFeSvD7pX3v+jf3EyTQifye0hgFp3FjLP4Zzg2Y4SD1/9UM
11/wfqra0UEJVmfmjpkZ3wLoAwmKgqmDbnFImEusZCGTB7YEFMHsc1zKXkrB
POibm+w7LIY/vQbrbXctNzf5DNDnWLZ9g2x+znK1+nv5ESzE+DYDA6X/ZUAE
G0R9rBARbwuSVhYbUZm+Ay2GSNOQ3TEHDrKmL4WYPApg/4iVwERrnU/6ClHJ
q/EcPbysqzpdW3U6ipme0ChQ6MWKkLoEPEx5YtxfVr38r4EnWPUVI89sFI2r
rmbsiPFDWoGFe5DohVvraRz7FdfgQ2HEYvvZHF6XHIIeZe7ZxRoPT4dlrX4k
JdZS/gn2n6RoZY8BmhuTr5uJa9bdhZtYF65lQnlVqDWozmcmfVoBVnxI7qFD
qgjt585SvhXe2Sb+xXfSZhu3VDH6ax95BLYgRmC5gloAWeWRzlWS9JT+OvXB
5yHAvZabB9p5XJWemeeGA8k+TjI7Xyur6OUNFHdvjJKkvKAf8ukzmxGl0zVA
8h88FCHSvgeQrNdpwAPAnHAbRMv4ytUKGA6Hbu95G8/dZVA5FaJ565vByHtY
MkW6UPch1c0YViV9RbgGJ/s9cmI3npIpAZElp0jw/NOyPAwg3o+VCYxTOcMc
cAI8PwvOG4xRmGNddrtZ+QvuBiJ/APQ9/9GdX5cOpsI47gJZyAUaKwMgI2wo
pnCEfyATSZrMCzIj2/SvJwG26fQZDGcbNlLZW3OXv+e+faj8FjtGtJwANnnD
c8SrjnCbCgBs4H/UiD4I4Fq0lG7RKA8qNbWv3Rig6fl6C5WCjYJ3eRs9YErB
uEPeHw8wume99xTKmhmkVpXgQJf3TQQ6KyJZhxpP9wl0VYJyezP6vSd3IwE6
qwDi0+n23EwKxgCc/yP7cbJADctCP4oMTq9eUZDOHvQf24R9eyyrdkXGHBCE
iuNAQf0gN8B7uHQ7m1257wcxR71TKCmF2oCJ+1w7IDQM3D8jnZufusGHL8Ky
VCizY2WkNTTYcQfwKZFg5HVvRQRxn0d6BdeKV+1GAgpfLpdxFyIoWodvRjhj
XLVbiwp/Rwq7qzJxF8UP3mUEQXKdG0DNL1fn9vAaN6zFQriEjb0hUA/BS3VO
HMG+yYgIxAhNO42zVq0UU1fCiSHjhpn21k+cBqoBSmKmmFHUDgiS+Q86Sb1H
STVPDvawdl4mo2Ifr/E2d8S+CQtT2Fww7lk06+OlzOnR1HEzeWRFxKLFwPa9
fykAXPwfgu+XAdk2CHs6YdD9kZW5l6EBDaeg4sh41R8kj2VIDy4hRThygqXW
kIF7jeNMCISBjXLj0B56FBjzRXwHxeLlkSMtxJio90L9Q+XX5vl01arhWVvK
lXdyHcMHzBExUB+RuedaLyDxmOeAG1lABvBkri5ftn1Aeq4JfSDcsYjHIFZv
1PYKLe+ekw7DoByiqUnF+Mww9wLGTiBxrNN+HbWgxftRGxI8amd/wp9jmIVF
g1ppnupdroTa2csBhv/FZVgQ8spK+sYe/qWM9X4biEvbMd19hvJG8bvyw96P
EYcxCctI++mjbMZ4RtJUbraGjvi/knttBch7a097TVW75Ap9lYNKgopViAHo
0UdMPNQ69wG8rMbpOgWuiSix8PWwnVdOdqBS+iwMN9Z3aiNwLGv55GFdyqyo
pxYEK6TOIdTqkU7lEBSbjsVdVPnyWzuMA5dKSGrxE//z41w43xqbmRYrK4mi
V0D5Mv1g2jv6prqa23yzamnqtlRkgvHigeS2wWxOm0GiRVSkG8gqqBxo09j1
FgKH9LUO0gq9z6KjD3fNqufA2xuLkFOvH2YmHC1Xe9QHE5/0JE1ttW6B8Z6j
oDfhkslS4U7HnfGuzICXwnrkGBoFRDv3mNWcRZkLyPyQMYisWOXb19sYgqZl
FKh9JEEYHZjX+LupFJ2jY6u7p2KnFbfQH0aL9u1Zak0sUIDMHBJen0GaBr8f
iEesYpJNnRaum5IycY9EkGkT/+SwU1CDir93sSycCu/2LOvWuuoLICJ4B/oH
3fqlnsoVFMNwzYBLPnhl8l3Sk8NhMwWu/VL2CIUZ8ht2CWz0AZeCHM4HQGpi
3e2JNaJ4SBt3hjbjJtVUtwkANdTkUO3JYSX88QlHlmOYFTRxIRCAbH2q6nme
UqRrF5e2cSVGZ9/dtwM3dFUoLg/bNG7/sHxOyX1BBEmVBUrYBny7UrWZNkG5
i045+gZbtmG63TvenidkCHHlSJfUcoqDmL1jIcCXs8eGmzqVuLmR61YLURIA
si4G0dw2kAT42E+g/8G0zwTK7ObD1NQ9/POgPa5NCyUCyOeXr/PMclvnWkUu
hHUEaS1mJ6fdBhR4H+hny1wo8/zP8QQSDetJvkZ0+xTqTpmIjDbGO5MhLH44
usH2Z7XWp6OIYYwEvVksIPHEneDujoJPfESsTBuhhaeT476w/yamhJT2ToZl
YgevAarF0p6+XMolAyBoj+jVY2rtR+pVKaZwCfsJLN6GwfQbkFBLXcuw+RGa
303NumZXzYcwDydE0rzJ/qiAO8OOkAxkdy1EkQVnKpM5wM1wJJIIRl2gKqew
TQOef53bUBw3LIYpOqb60EbUDBqfYTTz8+49ccR5u7E1JXaX8YYwHXm9dCBm
0O4m52GegOkxVNT3DYds2VkTHCt7uKBJUKXQuRkI26zT/MHww2meel/YClhM
Mc5kBRtO/Iv14gzhH0JDUm0ImRrgbEVTXpYh9+tN480qy3EiU93Z8jJyWit1
Ijwp2/uIieYsAJoNCqzN3vK4YvlqqxwQkFWk298LaQYDWxAOpNL4CWgw7cMS
T9SdrnsT5Bg0CbPnuFwZ1a45tM9NFwmJ7QdK0AXSc2dVsBN9Lf24iZaexajQ
eMLzR+8H9Z/28vOE1pWXUwAGrRqVluEzUNatUzCJZAQ62IzxYnyy9YfktQ3T
Zdv2keNhBIqbo8bWwo92dZx8/OUVG9YeFU2k8JeuOwcvFcrsFMxBfDogMFrU
Z5HBuVEPT1jnobw7GWvp/sIpG+aGuyd+NLP3AtNLD1ErJhEohrrUiehaCVn+
HjjK8kK52tYKjwIOyGJ6XcBWnY7aR/Ub0Ip8pdQ022zL5DvtyVglcPU7OLCa
Y6nyIeeM62PwVwYlleLJJc0GI2P+BzK3gEeiTQyXF3OtIQ2oGh8sB/pI+f/I
JfGHtDj2LWOk7JNpd4RHJJUtsf1nkVBui13yB1PA6f+s3u4kEP2SO0/j0hu1
SnCWXjXtck7UdGaXlNqXD8BJNG5iIsVegKsvDayehbC1gzRl9Os9jhg9GTON
2npd729P4fs0uvmSfvS+5nAmZcpPE0YVuM2uaep7NZIbudsqmnNguOQyQIQm
ZnJtw0NklPPCVj5J3NUKDsElj7zmTlg7vk7pAr/lOCWvKJx29u95EWTGgGoj
xBeV61bO3fzx/BpNHrZ+fjUKIZnIuZ54725RWtV+aMqCa4z3fx9mvANvR5F4
FmK443YX5adGsHlBHdxnRCLTmYmyyKkGyiDoVjxtjMwnw54G2J6FkBfFaFCr
cie0aTIOidEW1q6uUPjAk70Qki/eFBpN01uXWGIK1deXRqyRJEt8EeDWE5KT
G6hnf/KjQErdc+AOUOJWA7GHmBo3nY3gREeFSrnlG9FL+BssCJ2iaMHQybjj
8EEE+4UPSHzZJxD+jDddNGuOlz5pkwDl6O91ib6RTBGGCjfRHXRItP2CHrMn
nS1cJKcdYSwvXKtEuUp3DHjTrYFLh55tuJOMGuT26EzsRIrDK6tvj33jd+o2
2UqikJg5wpiYIo2Od1iG1QTM2g0t/QkRsFdE2AYQZ36stF3CkOjN5Hewxims
3pWhQld1KorKOPeHEFwTdHNXBlSHHsVfruaLQH388ISdIdBnHQ58oIVkRzr9
L4haUUavCjCCV4z9BEihllb/vw8LHH4sbfZI32E5WvbvIqhesJs9Mb42Xe+v
Gi8bDjQefTNrNSi7rbZKqLBQdMoeS/KqoH7eR1YikLJ+bLxRZ64drdzcWYeI
DwMLFrVJXxKgj7OEkDOQIa/XaIPBAqAsDbtkyJdrovY051qI5RlbWf/eEhKY
Kkq+XgNV96qA+xd+WXA1wtcGEsHSSYsEgVVWzlqVJ8dh3rlR5gxh3QN6YSFg
rIxkYjYvdFRH/lXnUNfrkjdHUaqXPebyAE3ppE7jP4PBeNLXzSb4ntDSOyEn
b7s9piC8/0hssayFfpE9VqDVhO8mNrA1PwLQQ6h1oR0c9wcvCfyaKS4TwKRS
U6fjPQuicD+TYZ1vP5zDpbcRls8br/ACxhJyK63kIGh248aL8f5xGxIlVoZy
S32Ou1jjG5g51gYP7lYllZsejiUmWh9IqLLU6WzNiDZOPhbmwzh5o/VZPIJX
9J44RLV0/pAHiVZQ1Xg8jrwHF9O/A0s+waBIC737JxqN7xmd1xTgeQ9YCsy3
xUpdSjY1Nqh82cX9pj3/kteF4xqx5AI8aJOciZFeqIEzNdYozgWwxK5DrWEE
9FEAewfDTrNZeOTNdTeHD1frALBWixmVXmUG3sk9T+Rk4ApVfZYU992/r9xn
lSDb0o5nFSxA2RQzCNPkHOGuPAdeJxfmWzmJqr3GwdEExUsE6qulTFTASIGW
+37/OW6XYms+jsQ/FWelWys1N1nW6cPTEgYraFJiH75QNbGpAj8XR6VxOo8h
AntGuST6T6oXC+E9ldfXOAEdWD7kKjskn20m+6rQqhiiND+Ha/mXEa+rhd2z
/hdTUgmVqvBDMqWgqe3eSOUOUqAbq1afmOambYXuyG8h9qAbZxDc40iMC5m4
42/veDU6lrz79jX5YL1Ia28KBRwfxptCrGR1AvhcxV2/GEEkJ+YxsqRIyO5M
VdNebkvnchUxKHZDh4nJY8P/Q9gi1oz6VIyqWSNDTVnFgOSHPv42ss4B8V7H
Gt4/7bOQaWCDZHkzUcF+zqd1f8lNpoi94GHeQfFVkSA69j+bnW2yOWISPBsY
GciO2NRhlK5Gz8Imt8DTGvmjbgphkKxyCWDCCzIpZoUHoyhb2bdPGixoNAPE
13960i5WIhdNgM9p98NpmfLlIo88KuPmhtgG+sjXdEV/Bm4aitDsAMWdJdB7
AtHMrxu/XEg6tqxqnzTSHT+vuHg8STlhAXSLqAml49yGe6vzxXRinNyrGjj4
RuCiNinc0px0aAzpL9uHYiTW71lreajvhqJWscykUy95HdigUeDw9yZZjRKu
YU1hHZ4VjT7SV7DrDa/LRzGWNduiu29xVGfQMGdI+hmY3Hr5TmfDYLaiz9fN
1q60khIk4oo+0DRHjRHNAV481WZlznSRddRvigAnOk5yFYgPC0sVet4btl08
q6FdhqNfNrKIJBey/NB/TQb14JPEnnBFQL21oaR3okSPSobo8LUrsSXpA6lS
sVDU90YTYd2u+ghy/rxS7g1lGwdPkeFA7cxv6NuU/J+8N/VDcdaOxAxIYogu
VYV2ZPAHpnZwvuY/H0BQ1uBusQ9YPHN73e2QohQIpZIYNAnD88cHCvDZRiaS
xlYFbT9UW6IWWj9gJaOm/Jt3SPOyBRB2+tE1IsyiRo8k5e/ixsRZmr3vBqb0
E0RbgbcRAOIXUKjrd6STZ2tLG3Yd4LAgDeNYDigTSecHCycLb33aUDCrVSSr
Lm41D6V1aheRq2OT1gVEETHIkVdiEs3J5ZbzJ6mP8Otl/j8/XP9Ghe7l2x2L
beNdNNYWV/OpoSFhi28WOtuE2QQn3Wqso25eVa+sThUFS4OAP7fdLKVQbESB
vVdpY9pqL8xgGN3BU5eGX5NWIOJcq24jdU7cJ1pw5ixL4Ab/dqwITIAaTSi8
H6ifkAcG3uucqRBq/ZWFS8nL+I2a9dkVUoMwrBsy1zCjq5xhwTy/bA4uwjSL
ALAgfzlOGL/YlFIBCOqyLQDbdvae5dH8cQ2KPxwwHch5ongEKJySzP/BBvgc
bcM1Xx7hzM+GUCb9ZLQYqP7ru8H1EPH2OtiM8ZxyA/dlZ+bw8SkdsnJJFVBx
/r67qsyhG0BZXciefzOUenV9Rl9OQ2NbQyB/b927z92PH2ks+iQDDPx0yxj3
NSWxVm0pbaUYXJ3HIBfjN5/DZM6cAfIE5cVvb8vOOq+QH/ZvBqrIEyRbaong
xd4i9hOtXv/hBHmkZt5OaIN3hth7zjcq0k67E1RMNlxCDzbwkLLUBRlU/aS2
RVxUDMctCAc448Q0hWm31n30q3OAS6GlqdHhWLcvk++TQLaUGNupQfKyUEFy
CV/R85d0MBWzpNHLapTRAdeJ3QgDXkdmXv0OJm02dt/L01iKnAezz+w7CPo4
4ErcVBR+3sOR+er1OmK0r4G9eLvi2OLfm9i4NDbcIGYRD8f+oyK+UcJHtaRx
dbh6NvpJ+lnKQCdw7RhgEbd3FTg91CyuEGtYCuxaFITw4wmdRDi5AdoiRaM/
r2I45jbFKHajOcvmRCcrQ3ZsVTOPtZR6q2BFFjTy2xl7dtET9BcXgsL5CZut
iv6A9OENlPBGpANUgZ8L/2T/IQjkOXu9cdVlf+fDIy150JpXxrhJq8b76NZF
MTsdV+4tKUC0/ezfNhJrXDwiDwFUnslMSwZwFuO3UadffBBeZme3OkHkeZvT
XeaGRdAV/hcEjJYmCwt2JUv70p/JAo4OpWGkWxvPZFbNKQ578zKNV+BtKT4E
efQ2s2meowU6Jj06wP09/gyu3wC7itQT8F1orXa1jZfRhPGghsANYsjrGos3
6tnrU5qI0cKDsKeLCsalE0lxFEzjzoYKdVpcMFIpG+3KinOzEHCUZkXOdOf0
nWENQaluVBod1e+DlWiyEXyEB8Hbf0apEjRTYK7kQqWc6tuurDje3yVCztmV
DbvT9vWbS93uF8MSlxG92UR+C4JPcNlErxxcwaRNyiGXZakpRa3in8bfoEPx
tspsW+kPNOh3P0/Ti/sh6PJ6dvVHquq0FTYntELP42sMX1dFyi/SPtbmcE3f
umswSRWxgFviljtiYuRTwkZFVc05gw0wjoevoNvUMzxcNsqVZWKYtNg66OWV
SXcOzQw70fH813G+ixqWHA0YJY+ixCqEuJ3DZ02R6JhiBcy6K2sSoLl/gQU9
htK3R/fO87BmwK0Qcqb8HwWug711ptUmUz9gEYWpIEDf6kvvZFBBhSxMt4c6
lX10voPB5b2T5Bpefc0JfIENvifHzhx+7itG/r0uJV5tPRuMdRph9lLLqSaz
QfKxptNqaVNtB37lc+wmMYmtuqnbF8VBUy+jNjR3qcA2uxgJ6cpp/5bGU+JS
LrTOtXaNE/YgXg894ELlFFbzFGleQBvloC2k7doobVYDQPNyUc8ft246ZFRR
jwhpl8aNc5oOcg+kZpmcy7FR6TZOD7nI5UttqedqSE0x/Mr4lTNavOFL2NNM
qtKC5mBf74ylRnc/AW5j/eb2gfPtRY/ymG4NCTvONE4rC7/g6C3Z8JhAFHe3
RBf/gYt6xizDWdf2CLaK24gVDK6kq3ABij0I1b59MwMCXYDPTOWX5UbExocQ
3PbHhbjOP1CdWbGlEnmZs9L0mv1Wi+YRuIZMNrGBW9YkULNF3vV9a7SMz9HW
E9c36cTjPhqmMxoAvhw/CI5I1gJUTr9lPYwS08qqm6dL5nRpzXID/1SzpbWI
JslMs50vF9kRKMEs4LhF05ZO7ACcSDuqfT6xo3Zk4vCbvuKPOU8B2ayJsUrJ
ficFW759YqYcUysUkJT1WpXuoTNqg+Iq6CWzJ1Bm9ZS8zMLRcXAyt3woT9fS
xljAxCCNCIHjVZCeMxvQ8wFoyMGmPuspKpuQ6SK6hQhOPykMMJ23nnWtKl9y
kJsYZ9yqbEBZwhSxJT+QwXBCMK5QBJbNfaclKHDoeJPL+vJCOggUHeRmUCTY
EwsPuGGhEYGh8SkXapU5BwRMAdiM9q1EJ10ZB8I+nWdEeeTYANKKsnHp/2yZ
6UWscQkG/TqPNsnPnaFAWZWgqn3eJAuDQ5C+04HGgrZfg1O73kC5rnQ0eDb+
D4p8xUoOefRbannncaNB/Qkxv6wdQbvgltDJwEnHLj7/1Swnqz+UMLOBYBRE
dt3fyaUGBCaHHjVDwXeI76lNdf4m41A8jiiCDv4fVOJe5BVzysUZl2TiMOpa
o6U16lyOzIaAjuUyQ7q8rzyz9HO3+EQWG5fUgEEnNuIuPUAb1Ftd7HQwuKQJ
RqrKjDQOjYWRiKG0Ntwld7EvjoZ07cxMuXdsYbmgxwPfKYgD5+tvhILKDKgn
vMpRnZz9xDGSMjsiL3BeMjyGZzxtdrNMxQf3H4B/9uTQJr8xdG0FwaDFAWtp
bgbDJ0S7Faj8frOFa+PzIo0oWs/f7a4PnT1Qdlmh+Q3IGZMdpSKgcrZwcW0y
6qHIKrx+v+O4IXawMVJQmHB9viC0P7ylEtFVQ4J6AzxdzKPveePX/LawAdUi
F9yTAuPNcVMw5mMsM1ayAQQER1yZbU/n4cNzq2irVMb00R7CCBivrEP1RifD
QhDaItwHph9KnZ0ZVOSljzLIPBTreyY1ZlnZFxbEerj2np70UkUlgUVfkutd
kJJMP7EVCmXikQVn0/JWiK8Wtqq3hyWKdeLlpYVAQUA+hT+eOPk1AQKLTMsd
mdgs+XqIXnibW74n7/3CzZNCC9giIwCo43+UxWhWqL9r+KsMMhrKBDIDgiI+
O6hBOt5emO1MGlgP+VheHUN4As0M2vg6td7a2kjAM490Dj5+9NaiGZPQT3SY
MFKd6nnqel30zKghg/7R7I9uCe/oPWi3T6LZkzkPs0zjBxVuYoQOV353Y3XX
b16RoUWG0ibUTI1bu+WVrsY4xfidt0pj+0FJvxSZ19FGqyfLwfJEvgHElvkZ
Ck859/OGXgDT6W6gfNEpTcYr6x5ht+EaqGZZo5AFQph64j9ZysWb2UGamrdf
/SMIHHxHyq1xIrt4DGqsgR1yOE4MxuDdumOPWgm7upr89A022GGiABxl5T4/
jaLh8/0Pmrla9FgxH0J8mQE4ENUWRahSvwjjFPQ7R5XAZ/yB++DlmTQZjSvQ
CFx5CZCfnsKWGgiP9Z/Eun74SVKFb1l//uYIMsAF41O1s3hhgsGK/eGE877q
LJ4ZlIBxVJYpePZEslo/CN51JWPWPPQYn40R5Bjt/O84DS+zjY/3NR4G11OI
wLEymZHOlXus8D1oUIyWcbL8hR4B8w5J/9cH6FjDfwsNb4hN9Pm+KuxeSo+Q
1upPiBwq3VK+hT44GJ0ACtQ9NmvIRp68GqTWlCrEmGQ1TXu0FC/Y2L9HWFe7
jCzcMi4AU44pm4tF6i5YiruMleH+kDwLRCXsX8+VTbm5OpPWIrtN/uOMVuIy
6Y0jzf7UjOGxpnRKxHvC7tDVKv47jWPcRsUW1G33qscITVK+cGkLReSILLM1
ws/lkO0UFOly5d1eKNxtAUabYJEDSZK7rO9/LXNIMGWd752RzZyTzRHrDRCa
mz8bN3rh8y9vS3Ajj+e/gveyudBoa6rpygHPXWrsmE21NRnKXss+39OiERb7
zEyUc8p+ljIoo5lYDj5cle9CEDY17d61uhbiWg28L+LQv6rFRpcgn4rrQQtM
vqoxYSlX5RbQS3OYywWlriqm67t3BWOmFnjsPgRQP2+R31N9QjPJNdV5SBcH
J/J62AvH8bX1V31O92AXRNOnVFivB59aTelx+I4SxxEqlJMO7fVJrSdMq1yS
keZb3IRfUkLy7hkzyaYq1JaXNQPPVRJhkZ06rrmfx6E5Y9xnVxK6DDhH+bMN
QDaKqbmIZ8hatAYfCEYLO6mqgytj37JUQ87/ZA5t6ZvbB2tfLoWWSduxuznL
zjdwIxVLBqAqQW95ykf8UyfUnwaO6POCZYQLoqlcmvEZ5Q3v35WtPNNvLiLB
tn4UTcif9JPIIBa0ppjiKudD1BryJTjHOUSoDVAvjIFDYGKPdAZtGGdqyr27
083UczidWNjZzlyWP3zCh8gXivR27YtD5iOSVuXBCMfQgDpiSwvDI8de+4Ew
Ul0uxV9TOpOCx9ybozQLiMkE3mJ5lZ0xleJiK2Rng6p2fwaQeXckmzkx0t1H
l16MYwYfd9TngYlR4KdCKuYGyLiAOCukuAcV3dv+D6RGYNeMERVinhr4eWXp
rW5DwpYtIn3DdbtC7LbLzA9IyO5blqAAcmqu6QrSgeDEZKdIsK8I3Xb+A+VL
1lB0fVMrU3/4pjdd25/QV80H6yKjSAr2xytUwdcooOFtI4FejgTDRxA8xEoT
x8BXmiFihwcSZ9IKS17YXSVn9h7QcV2H8xntRxRRM5NDIropBW7L+xGmQU6r
m02/1PFSRZC3mJLrM4Rw1MGXH3+latRfUIXG89fnJbazbeyCVaDVLBmkIus7
NanOmiZ7qm6Fm3BBQXsGF5PvcpPLho+kmgmPLLHRL1ZpAFi3NwkfA6ktHge8
7/UR1tiP1dbxW9EvRL6OBGdgf2wm+Q/x/Aijorl/EANRKE7xJ3ZRVOEKU1a3
2/p77h9VWLPPVX3cznWMxyuRX/5RGU90UChRoM+0tsukhR4Gj5PPkhFjiVCf
v0LQnDG7z1YWhalV4nT4QNmy7JrjE3qlPHNtlXancLbrgmj3OWX3odwcgb4z
2TI3zKl7LGlXeS5qUZ/QlBEhc4gnI7cndqiHEJgkbyNDzQ4g0fAmmileGFmq
PSjPl3GMmkBs5Zxqf5B3FgAjIxAmnGtF0GDjO5ZB5MyeJzjjkwOw296hDqCk
zDnPUOwNpx9ffGQLHxBUCBsFL0Kon5CVmOZMCF5juLR0ids0wGUsY7dh7zgf
Ld8jpBKg4Tiq0NQuP+JuPLh+6W+iVPFJJA9jTEpLL/wzhd5sn8nJdgHIUrBC
jDujmj7Q5u2YlMGNnxEG1hbIn2nk4Y/S4P8AXMbF+FoGwgmJAoFtlf7NDk/G
EWv3IrK3CDPTDRsuj4Luf2zPFKgSCZM1AixyyQ/hTLU85t17AP1Nju/QLUVe
pT8+RVQTVp+HYteeZin/ZHychtw7gJ7dWnuF4vwn33D95k4UJTnBvXp08SEG
NAOdkiBRAH32ovqJGk0cafdxkBkcmngvf2SEGfhPKJsWA2Yel/T3r11kYj3+
Ya1NYom7SRggByLBok5ykSv1yhOq2cAYQIrTQSLAWA8jizcmSTAZ7sf9VPL6
N5KwrflzUtdrU8k8SZJ+3lziJk8X2InjvsoDrTuQKqK6Er9dzMOFEW+3Avbh
zXkwCE/pW1A/S5ptBfZhyg/OJLQBU3VI7cpmYYrFMBYo3u/m7Ys32WBHNgGJ
NuYUl3e/j64qw/ITut2PLH1R9ff34GeFaKgsVWHHbvirH7abh3uOVVpQ82fX
8endW5GSzzFw5iIDUS6y3ab3X7L48I72N8ebnhROWm1pjpgH/ebH0HsbN6JV
8vynPTHQ4ElCFEtlw6xvncX7jEqqTEEnXycCGOf7md9SbBngADwRhAi+uK/b
VTh4mmLbHvTlcID50y4i4wz0HxY/dQQD3V08yKi5bbsmPKXtjKPowbqBlHg6
Q0qr2PTy1aAmr1tj0/NB9z3Vrnmq0EwTUlXGGnoZl2+SSw+SWsnapTu21x3W
yVPayxyGZRssUPc/r+DVE5ezUExOFNR/xtucPLS4W0HR+z+wFWrURy3V9YMi
2CHjyJpqzJZVwOt8dBeJRD9guVPxGRioF36/VMEvHfTBLlyY1dCzNloJhe4u
AItILZBKl/bU8e6oN7XoDftQovEnakJHbNL07uHgnyUF6ToalQIqcqwfLOOM
HOu1QRCTGfJQoQYaFIs3r2uUBoPbeOvJOkhsTW4ChOc8x2mh5sYTHph4lP0Y
dVgMZRXHnokjvtOeqMTVmmQ5HdycLLpGsPa3MuRZzV1PwEbvLt1XGZC4RqLz
FpUQRNwtMJlJzndHmQrXHPKTXw81SLOUhGpFJbSDv7NDnxGMLYqk7RdH2wf9
s7aEAKU/gO/ofNvYPYej1Z6IslNk8YjaMjrbR2dTe+hTtDKVNvjSE/f2CBwp
aDoNgxW9ebAWG9qp28GAY8iQLk51bKVot8Ri4f6vXaNIpp/alc9Y2FIVV+FO
XMA/LSCniOS1YsSQNBVSxc5IBbY+c1MTr89ETPjBBeywY4wPac3tRWj9muzi
TE6vEv32GFQIMqe+d2yk/DSRdB5phQUZMmBjDGob1gehMEEvb6RX6JZH1maH
oTHmAR1G0rKKAdOOWqMvQ7FMN0xOT11dBCdY4jT+CMiJtT1J6jtZmrHn3I7k
m6gLYVv0wP6LKBasI5Llzq4/kFbf8+Fo6pYMYKfjiB+qnpOh2rb1wQUeeZ3j
A7Y8f/8aUsEMSO9Bn0J8GLiuwbBvh+r2HAN10cePeXWRsQjrKhgygUvtyrAS
xvKAIjC8yRY3JZsyWnktdoLxmh3yBQiNdtvTyU70hJYX1t7cq4VWLM2lu/P6
p1sXmeY03KhreZxnr3U6nvNe68iST3NyFPFgPB3hdM/Khdw4a0NBPExIPh5G
PtTFzn3Im5uWCf4GrDmieqajeroU9xprqvQDofkla5t9xx5S7I94P4Mm6Vw5
Xfrg/5rPjbzt8nFKVjGerBBj7Q5lnnhH4qxj4A1pjha5V4Jh9ZDITKDjtKGe
RVJNy2B3oVdYIZA9lsFwDLggI2PpaqkERzP2c+u64czNKb9K6zr5D9E41ZD/
xJS1de04hQf9preNWqbfto6TlRzoYUPPx2WqXhZlO1d5nxyrjcuEcskfXIhd
Z8HoPemJ9CRSh/aH+k3OswwgTrgGJ7ASjuSRRbZU2xD4oFAlFqn3ZyEDG6Wb
GA4YLama+gD3mTG4VI5xv1BC3BxYeuYHstwd+s5IDlEKvHcm5xl7V3TKn8g6
9Xg+Q5mieiVFb67QhdozGzX4ARsSMNCoIT0YtkMyBwoJXuX4lkyEljoqHrQd
bSrDAPdegjqJED6rRgmcyhNuAA0eDGwhmxj/JKZLu0rDfRziT5h3ygvlBPui
C/qXmIxZj+miRKs/3mIylCi8B4FBX63KA1IbK3vZFngG+Q0KNR0V92yBaSRO
txAwxB5YG+4MpQob5QMAhrW5/4En70S6H14aH42eMK11ihLiy2XGtJBnPRg0
b8JXI5KOMkZvHDnzlUcEn9u4qM9LuswaftdzurIueRczsyvHJRcPQNPyADSw
tHoaN6km6vU8yCuedpxN1x1A3WFvkaLuaXbSTIJH/6BGWYOJiHlbs86J5Vw9
zMdcx69o6dP+buc9rscaLJWfUzOaeniCtBi+hgwETAfbeInTVZsF/LUmMaZw
brYOnduypRzvC7kH1QNgTT3Vy39yfeo2GWzA0LoawS2iR6Cv4ETbg6L+tHA0
lFgLaTQbfnwZg6u1Po6WL8xSwHTAm9TyogmYHP/rZYEo/Z7pHI9N/Cy36foG
tZE5U/51QSMVlDOYsBR/h6pbWub9Q6eOZqH3o+O4X41uE+MgY3exWk4RVZ+p
d8EfW+dOHUW9nuWfgc89JCvExTLkS9SbZvs32Pd7YRsgh5oxEHYCMZnWQHnX
YLh+Ws99376/jbJkV1KYSssQwgQGEk44bvFLIO54lAeXrsjMJLffpy3ups1U
0Ye2DR3I8kh6u7ntTJRsUgcEpWfam5FWzEgc17FAR0t7D5bxBCpBCqmhFkDA
gKe8bZO0kGC4Vqp4goZSrfCNdLDsOuFdIUz1CSaQCQJboS5lx3WAuiFg+mFN
qIFOnbphYVnRLk0TmYEhtOrag9qzBcr0vtQPvuRMyZ3e26hg/1X9jhHlKQH7
3eq94m3x2fRgaixC7Ko4r/BrN9LVB8LEXdIqI7ox/ZfVnHefOZu3FpPPOJgu
nRxOmQZ0LdB2/QupKF+HGmxuY+sJO3c8BOtHlc+KxMdeKueeS7Tt4I9S8zSQ
e+yhLhZNqEgMvQTrQMQ0dOTbFVkBYE8Jm2yttKJ9YtFZoP+wwXEqJAGK6u72
u/CJLCDzwpWdWLewg64qwFnWo3xNOPsID2agqJUs6iiU99oet28R3kphtZXB
l3uW1sJv4Gg+OqCa5HE+OcrDrzdOsfk9BIJr5Gvef/E3sdGLHQCWPwR+Z2ay
IQvTJQu8/MICS6oSWwf3uoM0ETGW3z9O0Zi1/KgIJmRmq8y16USJkRDcxpa5
bewwEm7NpJFdDGxjScSjTy/LiTCXscZFjlqwHZjzybK0UQms4blno7CTPwyv
QHed2c52vQp6z4kiWvmAA5ET++JFdCUhYsdsyqU64giIe5VAjPaSPYKHCPVa
9NzsrvE5+8Z9BkHk5mw0u3uQfkJwFLKtXY1EcZ0uFBBkozEUY+h1qiaRhXyx
7R3Gggvjt9GWkAviIL+W+4NzQlHGwax1uPW2gKOP/Ms1jU7G7kRe3QbgCzS4
42s3rmStKV0J1tFj5sQ2RM+fowVE1Cgqky4+YQbY1IT4CCrxRwvxwikzB9Hn
CyQkfL5kZbE0XWFXoDmgeNzONHLwphqglmhwumKB2jnQvl/PRO5QORtZdYNs
5zQR6objjxXyi/mfv7OfgJY1CAAVMGcNrwMgPOBuOXYyoBxRjjRPTQ1qiAYG
ZtcF/gNtUEbzSAT4XKsdAyx5LT2ZUXKAbkmwTl7XCMdzmdE+H+VuaRTM69cY
aCCCrjtwrMl+cFq5W262or2JLIZky3kv4M3fEfGeAzKkTN7yCI8UyO9s8g3+
bJ2adBrzOQ44srfapDPcD9QOq/AU4y36EoNetGzNvQctt0cTAk8K6eufOu1e
GpuSej74+8yPZOxxog74pKjX+aDM6KuVsrtb0jQ22Ux6XZ5NRn4BU5suTFeL
vOFFcci2mxLKld1VSPdg5dciQjWKblZoBJ4wHa6grqm+7o7qyJRPR4if1uud
sgb3tZS8oIRbJ1/CgHGYZqvzQ37IjFwewrZThZiiEzcpgFWC7rTmvY2TLvgl
BuMOsEsVVMXqAfx/96Eh/SH3myC+U1FDCZTP2j7m0LQIzv7tAPIIxGRu3xfD
VtqQaCqkJF1ufwhkkvXRtpC/X4h4cp0euKKFkawt+W8CvgWpuYXp/z/bd2Sy
x9diuljuz8b4U6/xgJd36toOB0T6CrVDxpAohyJ79GZdWyb9hJgrn0TwHq5w
n35bKoGWK3vjI2wq3rxCI1Ltvm3ATiuxu6XH4u+HK9+zN1uFLRsHxfzOvmPO
MGtGDNRUgsjRAJAZ1SfF4APo+/YvIQU9b0GTkh0JlXu+6vjgfSX3QrYQSR0m
Rwz1BRTpWIIqqMiKS7DannGpFFa8SOZ+x0uabuU5KZUamDFDci9YQddVzxZN
g0kCWDgax6EevZJzdrAJpoZAjd1M2G0rfS0zNoFK/fuQvUhiDywzpIto5ips
LHOYR1O280y/eOsVx/9kYq9mNca36I1b3IUTpzH6imhRaqIgG0/IeCDGlIHk
D6tk0Z1rKm1blQnRCT2D+/4DHHnUaljz0P8PMerdhU4gnQ9McSMqyJrE342D
c2woAombrxJCGw3NGcwrV8zpKZ4IDasSvJQ0b+bNvT8pRH99TDw3medB3y/s
Go7ECtAPFO6K9mnWzxjmSr1zZyAS9EirQBtBXp5hTtrzmqxJu0gmcLrUvZtV
lo9R1BCgUs4y+yiE5COUu8i7VeyXEPukQNFAZ41ZyZ6gdVwQADWjVUbPfXRh
0a2H/dlnVejSY5Yty2e+f4IWiOoUC71arc25I3pEaFkwXcVjikNhWPsF0Q+y
WZ+XXGA/WhUJURLSTjC7Rh1AZizyAtDf65WUDcdOB3mOhT15bokilNQ/TbQX
FDrWsLWyl+mdgMv0pxirwASI3nIe2eiOvG+UlFg/hAoladNc1HcoepM/L8AT
um2J9+it4ysT0nAsx86XlrOHmi7n3cPjVn/aHccnZos/aU9lFIVedZ/sbkYS
EwUN7a9aOEADYxiE7f1LEioHhNhPFTC5Z1bvVpXczmdLu6KkFovP7+6aYdM4
zmpMhPY/A1QUEBtZfFCdI6XOCCvmGEcn07BU766/WaZvPlY/+Ny5ArdtZyJq
bGKV+8ouJs/DFhDOfFXEOns5E6AKcEJ/WOWTiImt2jTfObaf8nfm2AgZ5SFJ
eO83p8GFteGCcx5YZwPjYVZkDkkGcFhcMtRc+5a2EihjWhJOiARPXM2gHHVq
8rbAZM9W+HonrbGCFZVS7qgdACiKpAZIhaVZ+7hW/lPwqAv/hMWoq6l+B8cw
sO6+0fTcj/K3A7xRIY4QnPQAkcWvg5mlFyZd7bfIwRSfXLv7tUmrUdocZmor
sfS/NGeGoe+JHN6feCvAC7LfOSeyF7ahb9SQBfQOvxkDbIyhkxoEmrV/QIMl
XkXBn5vSnUNdZDL1LkjFOh3UUmVBHb4m8nRhBm/Vag+IaDJz599G4OjDXtNz
pEfVDvJuxHfADZ/bGxlLaxejQJqQzPp905d+PQrMwRlYw1AtkbzZhqtFY0FM
bQe4wqQJ+CSZJQ/J1FORYQ7EH3xJwEBvE0QLa7TPZgyJ4s3LA8cn5l/oBuhS
+0ipktObi9I50uLVBm6LnTPB1J+oZu2EO2rqbUVVKZrDRkIfaU8y9ujHibtC
pzJnz9gaSXMev9dxr1w858w8GDAbk4RWDiZ9IDdj5hpXWc5KOvN87pajHXsD
vNNuPlLeUhCjCNS5/46Hy7G0/XwIaf334BtgdxUkVBtn7ldlLATHaRu/a+tF
NBpWpjoo0q/0ZqsV6Fuyyi5a/JUO6By462vtrpxC4iDGArlWwzVtserM51tr
yyK/d5XtFfLIHSZm2L1qDWYjTNEOdar77JXw8Ec7bJbiMd3nnhRRpOmpZ7pw
69IO2vvqIMieNMfFq37RDgEH+3Uidr1FsRR04KiAWw0sPBHZFetMe37Y8oqE
g2UC6P8awFT982krk2CYkmEcyZxXzIjXd2Ke/PbxWLrhxn7cYi65F2TcGZWz
PWagKjQCVt1cQv1cqzvA7feyqjWsdDEXbtQBLSSmLSD4EXGKLjQu8hklvMp2
r5lqBooEWHgZensf052jjQX9SCWxdkxO/VxQoC+Io8B/KwbnvNOm5pHZ2pYF
eIRZtiOvIlQTCX3OmInzgC5urRT+5lblupHek9UieF0fT0csGu4pM1DqVc/I
l+BaCv+X2nTbRKfyWvFZNIlThNBlKkrf0TTNBjtVOsN3XM4Lfuf6PpGSshq/
fUY9DwA8XDuD2u2AAvD9hwuG3GmW4SDOmJK7awB0oLxE75AHYtORop5erXic
HQll1XcCQ6MZKbvhk6QnUetrwEHv0Nsy9JIONFSwA8zZ/iuGs1SLrWOidBBO
MajKFP1LH+inS+sYzHxYlG6lByclM0TImRWNBCEjxhH75KpbPh1Wi5AyoL9Q
4Iox14shQDQdwjetLrVY23SV69fjzsom8wgJSVduGuBHr/rkTeOvyNOb74TC
iCcbNMoXJ6rnUjvpdiirV9D9TCvjCCCr2d1BmzinFfcwxAXJkSV8OPjK0Guv
16nu4XPlCTE8GjhiERdtzrL/N3Gwcz8eb2Ha7Vfg1LOe4j7hhjYCNqktBQoq
lZ0QfGdWBpai2vk4XVtkUk1P1blWJHrueAU1T50RTGr+bz0SHij/l0buFXwR
wVhTgzuj+YxDXA4YZKWOxvidF+wqDh3K6KJXxO6TxsKEs9rt350W+CC76kP6
5MkWSXlUVqFjK9OcIajS0e6DucCU8TExFUel8F5k7l7e0CMr74U+OKm+4yLX
9wEkq8AhppqtEm+QO+HZbJZDJz6Wgc3xDSBLHOxYuyhH5EmjORtKNQPdBZ/D
CL572+1s6T6ijf7Nz8nmh5mLQUxgcQmUZ+N/k/Pt0PiOJBdbOlQNZqlNOk1Q
lOER5SAVvlEUqNF2x1j00gz2HZVLTjodcyIdCxmcCR8F8H4ut5wZ0q9uMDTH
4Pv28W6E39BA78DwTyMIX9+Ebvhw8g1al67VNX9SSydz+S1TlFfrlI4rthWk
JvVvHkXunwno9zahad4u6vzJkVJ7pEZ5v9B1019vicMx/vF9Dyb740ZfBoPI
BSJyW2EdozrntSDyyGZghvuBEkxEVqoPqu0Hd1TV6+tXK1wjfW7w8sGnvYVa
jnjGeFERkas9O8Fy+l/ryue9121+aRtSAjXQktUZHnZs623EPxOQIqQc5Syx
9xKGVSJgCl3JaKlPhugFiGd4iplCH1OgpHe5dBEDmlKgdDOaUYV+kz51SNKT
SziDANS2IKX5KTHAkUU6TxGow4AXAw/LItMxIs0ynheLUI9wH7ZkWzFz8Xyt
j/tTDuymrnD61thHCnSGECUJ6h9QEmPmL2DPVGpCZkFQDWajfHKO9rxGIPZC
B+PAWDUxVz1I2djRtx/2KgyhvBHZkTefu7TxLcaSv2vDC27il3/1W0EPHKsy
+ilOhhzcZRNrZbnmfta0L2yc2VuLvyFKduCVe9745jkyezFBj7Nh3wXthpqv
t7/eF10ndeSnXsyv3y/O+hdxtKM2VlVR/op44GY0F+iVmXhPHW7chsqbc/Bv
GP876BmVTBeAbAQ8d8kTRk3ChA6HQ6/aegF75VJCAanWhYP2XyDLXVPRZNhL
K76xkze//hYPhxPXbQtyeFvAQOHpNkewD+Lj6C2U61+eaZDEPJ0IvWOaxiGX
IryrrfUHg0lyYwi9E+jl34AcGXbOcoSmeDOOyW8D4RAtqdMfnfHK7vs3oxqZ
oGFiQZvp5fnT70CjH3JXfi+vsde11TrnvGDca4Gf1E3uX+Ks8nat6TCedH6s
ihweEPh3r+vHB/wuLhI8PI4wl++JUINItPBzOCrsZuR9fSlJWrbaghg6NCpf
jQZ4YlD7yWF5b04Y1UW56l+iC5dzHHt9GYKUN0qo50REkjCUMqRoYG9a6UZw
9/qupn4RyAObVfB+ZZq0GQhHmYqLmpNg9qdY00wHTQWtuU/F0KTAJVNJPu6B
SnteuqADJrbtOLT6ao5nXE89fmw/BZR0W/BLoK3IcxKR2rq8g9l30+q7AnJk
KjeNk/eEznoW6oIkueDphLC/6jXEMCINnWKozeoZyDGiDyhXfi5hvrdvbf/1
sTOss93XNwiidFDpXfSzOB9QEkvbBrzBYc6bmCK1XKGBG1DygDksoVSMoNL4
+zZOHVeRvuhTSIHeyTIPgPK8tF5bQVtOmsQcZXsAamzzY7EEwBdpI0AA6vru
jwa/U/4KqIbwuLZ6SVmlF28cDrdSSzJnvdt43LMM0T8d7By7KirSHr8+Wc7o
bSj1Eo66IGFU3Jhm7lgo0ezOQw2kQBnJVbYWmomPuaJsvem0Rqw5MyW5y4K1
YpUQWTZCtdkVUhnoDLj7HZBAUwz1um9IQqgMkGmEj0ND0DdEYyzw2/7C0doJ
FdXSHZ5puMirHzA+ISWISS9vwgvVnVADGHIrZ/wIEdCWYyFrw9dsi5edCsoQ
xjd+haeorto2eNDTpqNKPZ5sF1sxqBW27ixHWS6l8/lTH+m954dBjlyQqQp6
Z99OgOJtdNMu5V2Fw43iRfrsebLBbvQSaJd9cvItpl1l85CoCqYA5Nu2FVdK
IbsKTlba9Bo1uo9Imsr7MxSzZEjQ/5kwy5cjVJS50H/cCW+kLZBfEVi9c97c
yipSIO68GF4MOiSJHQ2CDZbWvzyjX9N1Cdt1tTKIg1QhzTI/goNEJQuZrRsO
zqzwhN8NLMULP9SGkrsJ/xBGh9M36oqA2LER20Ko4DDUEEoWlDmw9Pp2Mi4C
8sUkvjnA6Gg/g1kG7eel54sftNVZmsH5i7aXp1LTffsUjYCCDq5gIt3gsEDT
q+pjKhGovBAg7WgCB3FJox2hQYdg1qHSDbQJ7OA9UikMqlsiV+IjQOA7q6Dh
3TPsBMaOUdwkPsvwWScPqYif0SM12YAgwJFlQlMIKqSVpr9fDm9zymfku6TF
kGdcD3BQLlPLLIWpTdZp5M+79GXjOdXQNdPCE+TV0VOmNZSZhae90tCUBphc
Z0KKn/EHNOU7468V/9ySYkE+NJfXMEAK2cIapzPA23Qtb8D6Vj9J7B6YLi4A
suD7Df8How0/6L8G6t2ZsFS/egWAhtCOlqVitkKpcUIQ84hRxFPqaU79AnQ0
fa5/a37LfveAkfRuvHX2NozjjYbLmTgh+TFtFwNARMx32obUQhFGWOcFqtaE
48+KG5HygdMAyj4o3KYKt3mRZ6tki9dfe8bTBeag7smAxOef1i43KYLBQSme
AHf1lbejN/yYZfxURJ0NULjWLyNQGOWkXPVn3jC91QtpbCSTzK9uINwRXTpC
zOOsg5do6JfJ7fxSmglzg5GOTIsyKb5594b51BPDszoXj9NDjNCSodlyvkJz
CaTOE2+241TJQTqlpH1bNDeV4m9n7rDdIo6w8rXTR/gLhQFOJWpjA35aDIrb
QPcTp8Q1S9asbXlpZN6ir3gPFQ2QdvblUuturoa4wBF0Vu8pg1qvtBcIf6p5
bTeSCJxyJJRWl4Opcod+7txU9Z72fE/hFNOFSk46I4mVBUcmYQXyrojF2rMt
k4suD6hX5G91A5qPJlg+so1OaOarT4XAihPHVRD2CPkmnlvGHx2txsH2bwFG
mlor27YlD48JYQOUExCXkDc3cTj3MB6eFe0Z7cPEJRj7MBC/w9Lhtt3e6GeB
FiMFmHn9AiTGR5lhwV2r5dsEIYJfiktn56JQUuy/KBDZpylOSuFrooxJcf8s
EJkB1JQZB/fauaYpDsCfXqegU4rQ7phVvCdMHXG4bSdNs7BuntqgJpqvkrF7
BOkMCR+y0rjFwsfcZ3xaurQzKEmCbIjtm+pOGh+EsJZNDOwPISbinIGjs3t9
tfCubvxOUUfSQNy2DbkGPCJaIYdZAumd7/edDJlrzKwjw6N5B9EUoWDS+gkV
fpz2IpZZBjBPZQPNeRy72xGWUkKIpwAC3X68VMurTvatYb0ApAKSVkwDx4tV
VvmbuIQYzNBgziSCyUpjz50LkylgBINYmfR84BGLOEBKDAxLyWyjv1d8zFHk
m6Oa3ayLKY+fjaHra2JT2MeDkuWa9+TQIkRnVMSL1KWeZMHza5wbPo2u7/Cm
8wWscQFfu8LH2EuZTjOJmvsV+CIT6cGeLdW/QoL/v40m4K2nepKyJ7huDb6D
crCwJRvB3ZCXmvd1Cg4admmgKzr12yaXS7Sl2nLz6bUEqF2GbuUlMKhVurdz
1KwW8eTt1juaRhqhpgUu317l8bF5J8EBQb378td39ykoHT+kSZtNFNngdV2X
wUh9K8Kt4nO7uPNtlQg47z4RITWf0kLqak6JxIw2yQQK6K42FKRji9A7Pazh
GFbc6x10OpQZkNX51bOb14d4SasWk9/BaRgQDiF9mU+74H7KIPIr6ovHNNsw
vuVg+tkMLmaDhZ42edUrCgywUBuqCOdvfjqdFH20vkJ5hxJRkgqD4MF3yCsT
d1T951YN4Z5WJOep9kTQs61bB4LEDcOpGyt28P3KRURAFGhzC4B1klXqlz8n
iphosmDo/zACLlesPz3MmF5mV9jeqGmHZD3NtEjYKK+BzlwadB2DUhPbQXrN
IKEgaJSIPbo9rgpg/+uBMu2J6uaewwmGTP07jEGB6HGHIGDIoPACUpK1VcrG
E6gZzGj5eJ1ieeRhzR2Z9RBBQCs6TahwCHfWdSeJQzRDaQ+uFQD/ZTOpeB7b
rUAnD89Zg3U0xmgAaeK5q+x8DB8DFJwuSAWTD1beaM3P/ti4DmV5EjsvbfGn
m7IlN/OaHTKFEiSJZMpPG4wPjvun9nTyOUgRY1HMDuBfuISwlISWpGEYZtin
INz0iqQfKBajLhNAmwmYugpjQmSkvH7iJnWaCgV1GwirSdNAhBSW+askdiY+
4tNdfufsR8ZpCQsx1CYUVKRfljkBnMVrg3lCMa+AJC5jyukLstKkz/Mmsq0b
ogNXC4PlYXTZPckJv+akOGaScF87D8R3YYEWnpxf2i6AnK9QFwFyNV/mUto6
ieLSYjvxdWXbtYENyHk4tRORHMColaoPYkTX6whKET9MITkU5Iypz87rw2At
KyLU+Aug5jShsdmGBMP82TABSF+LlsGhS3Q8hOnkSkPCB+xfqOBN800VnxRd
oLC594zy3F1WjNhpHVLi7tSoYuvibWLgXlIxgjlGpwNBC3RdaJADQqq3d9aC
LSAxLVXQVAihHQUDzLiqMZn+QtNfEeDFAjSCKR2OjqXZzlox+5Fv8e6gxxxj
3jR3sdkdbalHM+CwTkBw9NcB8EAoD9LmvaA+TY81xHOTDgt3VlF+MD8HxxYn
RakvD92rP2RwetRXSpu0smzX5ZghMxjLBhrq8qZYJOWtK7MlBv+1Pk0yzyya
C8U1gM+2act1XihmNhEKEHXXJifP3uc4P8Rg9bl6PcYIWe/7sFe+8gQMoaBx
qUt8E8RvZX4IXHGP2sWreMJ2On3Bon1VSe9ShucJMdyyjfvRY2cowSRBoIMo
plYVPwFCtlpYOC9gMTi6/YebvWIcMwayZ9qpEWluInRsaV12/SqbuSlN140r
u1TGz+bOwh0Z9GQD7+IKfzgzoi4TfMiXiJi3r+kSHQOSnbLKjOgvf0dVu1JF
IGdh/YEl6nvb1zM8ek99oHyWidabyAx7r0NXKyFiyDzXjIg9zU514nnMef2m
uH0hfj5np74fHrXB9x+XMDk7n52Eh9ka5oE8jLVMOQ1dAIq1G+hptgethaYo
s9ycGg72rYSQmypfUOQlV6++z9b11nYQ5z6I3ZjH9fZTQlfNZdEL9PCLhLy4
K2YSXNlKNnnHAJ5+iA5yeTAO37+L9oXGlMgpnEgucRHsE6ZQFY++W5S+Zjqh
GeRwVjqUpfx/PAHWGqIbLP+ra32XzSwjyu+fQcKG3K0824Lq6mn0fr4RTyc3
3BbbLR3CuJ+p3sEEI9SxZeoukLrMXhko0GiooD1ZT5wz4NIPEME/PVchhRG9
XvnIqkYE7AZcJ2qdv//HMupOBm6BcaYduba0/B5qs4YnhiHF+HN3GxPrOkz7
GW4isJ3pVSW9otNvBTneyYjvJCDwy0oP8nLRN407Wna9h8zJWZ6V0mpSrj4s
JvrnSj2WHdJoc0jTEX3iorD6UoxkTkBu3zIJ567B96XjcVH9JemxKPk3RTsq
IKRM1z2RhNKMkbCjkIkVv8AjnJJzI5SXtkDz/MaM0ApnuQLSdZr3W0kUiFbF
o2/lJt8hbGU2ENsVXrxiCsRNNNRRoBZfxHBsts9UpGslvA04qjSXHWhZEAQ1
eK5pRZZcIoT3ToPR23za8mTrYbhGyiT1enBS706b/5JYhY1D0ttMqxDtp/Ay
54fDVPgeMGWsZLHGrSoaUo4BcB6nb3gAVnAWFxJpKHrcKqxlaZjBEYfUz1vc
IVuwGdkwfwX+UO86vW6TdJbkizMfS79Wf0e81A/VUgz7YA/n5PUtkBdB2R/w
dYBR5E3RBkjQy1aWnp1Zmc1B8nM9sHAEPn9fTbQwpUy4slGumQpG6HreFvkV
JuOboi4dDCoLVMc9eJdgMx9t/idN2U6VqWmjFHOSbVf4NLbwhz+XtX6QWdvH
V4R8TKNTaPW3ue5ZbVCU7htLxmQqhB6b7uWRht05ONPjY7g0bddplUTOS2lv
5c3P7XJpvXeZAydGb2gbE5KaprKUO6jQQ6ey0+QA5H+iHM3Qh8h4SddsEbGB
xGCeSeoQBNsESqQw14IrY+65sWUSOcK7oqFkM6ZXeqArtm3V0F3Dj0bZ3aJf
rlWpA8QVCNb/SAK+muyIJEHUVGPG4cdcvGa918MePM6A8LLm1MfTPNb9EPfk
ycXFbVppqmysxW9nto0gfDwU49eGGnl6j7RCVRLzvMLqJq1EZ0M4+iDtFFdT
IV/J6v22YsVGcNpA9rgYZewGHiILvFbrB3Ldu1wn+acci65Ou12q3WawqtZY
iklAFnxmKNWoaAXCaPiaupqNMp1Ak21Bjw0OzhTM7hclrIVicke0U2pH+Mt0
o8dfDhUN/VyFcr0puue7C6DY5OGqJBfhK7pcBkDgfDpDCmMPsDyN4aSLFgMI
drspuTXjPugQaYPlKGG42M/XqvfAay6xsrXW/XfwXONpwc+1IHl7OHrabaK7
Mi368ack8aYi4FT0WkJ+Kn1Q2Y71AHyYkINPyHjy7xuX/wv9fIvIaX+BNeup
HDum5sInzpewsbKgUfOf+BozRK+X9jh/vtKJ1IX4QWsPgp+gcnSkW/OJvh8U
9jN2/E/jih6XQkGJbCZWcUkAlnmTJ+JfkHk8bE1LMtKGfQbArjiZ5yv86c0p
zLYZJwNHy8vNDgSBdNVHi9i8poaCWaz4WBNc5/F/03zHyVVxD+cJPTHpSg4y
ccKPKNq1CrmqO37FIJZqreItSi7/PbO2TKRNn5UTR3xo/FMxiL6EMC735VpT
Is3VgYf5tmBZ+EUqYyoQeY9V8YbW2eBJtG+zyhvQseZh3D6i4DT3zF/1AMoZ
SNg+Jz2QLwPz+W/NuDnEy88gfipUD2KA0dri8dpnisy0BLNjqTuFJVOJCjJi
po404d1jd1bdx5TfXtywTr8H9ZcNZB/KJ7Hi8Pb+pusqbyXRZ8jo+JgwYyYh
sJV9iWvyqXntOdDcHETbwos8cq1CCj/+ObUEGamBFBPydGctVeN+aIHPCCdb
wuor2ZgaY2s0UfMEDgP1LJ0tulrPDqZqlhf0KzHdxX/VldedHg05tvIV9dYd
o7Lennl/LNgcwxGVMw8l1LF/e7gJRSF36rsjyse/8wJNSf8OpJk6K0yKKfJX
EfJ3iG7L9gQ12Z3JBAyNZujDPsGI8u32Oz4rU5kinOAYrIygRxo8x5+680Ol
wzGnlUAnCbQu9zJAb7g83EvYVlkouHMNs+XK56r75DnkB1KN6RDw51kAevYi
nwKwX5dm+oGwSHYDd9SJzhNwS6KnETisxG/CsRyyMO6rrekax7/qgDEBDeq6
MYcs94PnSeilochcgkzVzVHWo6U1nh5JBMkfLxD8UJdalP6Q09la9KIeKesL
M6bvONoKevGEnYNWV2zDmKwFDwXsnWxgkmSBzMRq3MwgKRqxgJpIAZNOSK5h
9+zFzfjLaqyU6EP2tqWUQe7HHsGsphPYSKPPUdUlQrxozRK7yKeWXksgNZ0e
OmQD4UfVMpcTblbyhUHBJc+Jow/KId/LlH9pygmqk1qvZIzE1t6S31S3XNUM
feQX0TZIO568tz8WXjNg8XK76iT5Qu/sOGyvNbtwiuruiim74IxrADWPSS/5
zpuvdth4SvEP0wwW0Ur6yVwe0sKrxBgqI+Z6JRx6/GZ3lqswbHlPSUlKv0e4
Txn+K8UUmaNLxH9XMIk9LnUlPocAsKhdk+cHNh4gsVKZEpm0wQm2SjwxOo85
6CbJ7sMa+/AHu1ePQN9KStjxi5tvzJSdRbI3OUs9+GXUFhe/358ilowX4sbc
+HQfVG1ZJaOxW26B/HO+7d/Pzf0l9X/tZB4CkpyOLDh5xGjrZuAXddzj5klV
sAZVTe7yLIj4ZgBSKvRY3so1fa08vOmv0LaiBH148hGRiN/VBdT798wfk3IW
AAiKM38kWsD2vWg6xH/8OXKqCO5CmjDwufqiRQnR42ythe0Gh+KJBNnirgLn
X/Zv5uCv7czNuIJVH3zr0l7xIPoORU2ovVAIk8paMN16DZOUcV1yJD4lK8Yo
sk0DylhfqqosQXLPpatciVDrYMcsFlc814np309I44XJlVv5cdKgo8k0B2v8
K8HO7oKfPsE8FLCwCWKYzC7PmNin33POxV99p5YoyCa5E5UmsiFmKvSGWk+x
EtYlV/EtU7M7IY/7I7bpD2XfZeuSptK2tum+mhdELHancjXaswgikni8cUtp
flDbZiqsnEAva+gLNg3k475/NGOZM0ZKvODfs2l7fEuakGAAfK8TyU3xQ8pR
63y9apMFNlGb07V+/NSbwxO/pinIbW8PjUjfTlMjrM/zHMFtHoTo6dkb8/Cm
b4252Q1XbbbJK4ctA88+QpZvSiharFp6+tI/fO4t18rLdX8Fp6mumN+HGFlG
IOOa66Kw2v0bsPFF50f65RMLzXHwG8ha5n/MswSMo+wWMAmqbs7MAXD6flgV
ZIAFDbTTrhs+gD9h1tQN4KP2y4mLRFg5p5s30dcZ9G5jx4oOUZS3Y7L1DnoE
Uqupy1DAm5Ud4R05INLMcgf9dO2qGrydFJI+jjOzwx88Sza0k8KbLPN0Owkb
YH73MERKXrfLZOdZ9IIr08YYNrytVJauEanCq9SnCMjdH4btbTgYut7VewA2
YTRoeOdeacmhq61Bwra9fwmF94auZqYaYZ7xD9EAtAhIs/ErpRgHOrFaWihc
7JPyQ0Zp66McVN2isCXk8BT9FT1HGMjHNTJqNqJzTR5WB82C90I1miVvt0kp
4mTV3rm+w7svkpkAKMd+QiwiBq2DvB5FchBtF7elJtSS5+/VVYbKl4BVe5mm
37ayVfvFi5TOWgEm0JjePB+YvnncaghPAp/OYUc7EM16b457+QxiKcf0eCx0
4ct16LOZE+0KgND7J1IpCuJxQg+aG2keXtKtmw8tTNTrvaqYB2USF+fDdctQ
0iLR2EyXBe/MvIe7Snu3qlK+bSUpjZOGnWpPUI+sNBOpxRZM1Z5UcF047WB3
GG2lwXc3lqoS3TcGuYOgaTN4NUTDFiTXXi3unxQqe2N0VX7y6+t2b6SDDmbK
BgYzLEUURfWYMB1OnbT4luUXCjla7niDyYxbBfzhjdTitmcAaISgACVhGlMq
LTnPeYbPOk8oYr6rQLo0uwoZCq/wPIea0b9UbHFdQldyHk3AA2wHLsUpsZpV
mPrivaSUGaeOG8ViAzMfnsehodsCHS2RLJJf7Edsyj+lh3lFFE8TgOGO5q45
F5XZLdSITUlyguTMhlJisvtRXMbNmJ14XMRPceo4TmL7HCtSaYqzpc3OGdC/
yZKe/uVF4nFNcOTL4RV+C4XaTSRpFiahixRQQFLVCl9AlJbe9sJt5+pVLicR
pSuSXGRHmuRxRpkRbA/jkNaRbR5NSXThEtGnASbdKcrTTOW68BAQwzjkhTDM
tDLnxz8Bt9rTlXmOIrfCfw6O+g+QEzHpUlevuUBuIM9eNRaiEgr1WlvQhTFF
YR8umTaEB0kuemfBz/Yx+vrOmxz3jolsdNyRARCRHLPVAnpyvwHAqdKCNqJh
TZGjMHO4exxZsZUDCbOp61zL1M3zhfXu21p1ZfolHFixV5UDxa6TzoOOqjwC
aB1cte/N5n5HOSEf7DjKp4kXgKtm3vNcMKRbGPdeHEGmU0xn7rr3vOxK5Eaj
5gHbplUYJ5cJoOF9AYN16gjYc0Xj0ojU85lPHgTyd1E6yhm7sMrYZy2gD/XN
OKendfKLxxSQNGgfH8vsKIgDyWMKL5wTOX1WMxrPQkDMeYUcDX53U/06i3tG
TnrGimr4guYvPd+l70ads826dL0hPKGOHHfiCzOI7IcJD/5y6QNRme0eooeP
/lyD5U/yN2hB2yPnG76cIkboqkQRXuRDjsNmeXjqtnRoSnzufF4KJTsOYLIN
ObQHwaMHewZ9SdDqQh8/IjhXGuZnQAl5qQPvj9PVwuPIgFZyjUGaj/dINj0x
8d57Ruz3QFqLFPKdi8/iO2XsOAPiHZWkwXCdK/Ik8O1fkHM2kTN/qkYo33Rt
UhKgkM0TfCBIxZQEHOXFI671KSiY6w4CPEGS3DCuZ6Rr8QGP8HRnuep9f7zp
YevI6IyGCMuQeyUyV9c4vBG09IZPZM1DnD6SwVJe1LzLy0vGTGAKDa1d7boF
zyqDh2mzUGR095ixlFFgnOYLYGyZVE5eREiyBbmCm8cOgJfbL8EzKdX9XeWK
K7RMLxfOslvXo9wORwLgUIQc2jH5d2KRQ3tTTJnSoUBQe1a1FdHunvO6GPhp
zieU0seS+iOSNUy0UFfR/AWxsRuXnIhU//FH6vKOu56VzqnUyUu6m59Z0W5l
ZBf1qEpBlYBwF3yxouC9xrH/uQRWrmwXvV1VpWQ9p3dCyNMoZDO7VPQdfB2D
A1s/KUnhHBbPR1k69KMJf+8JEiPyGXNLXGxMjhUm9sMLLX99agrLkLfoHKGE
UwXacHZs6ZD/7KH3/zDzv74nVY0IKb27rAjYNGV54cvc+tgYPcFC5c0GmoOY
eWOhBaLw3FVGw/bKI0q+7qkN5n4nD8bBza5VoONaUpeHWXughC9l5uBVCAai
IiKAgo4OuucKCjdeYCfFgYyGwPv//0alQP27dg4QLMqHluz38R4h/e9DeIoA
IvbB/sy+pC6qddFJrEJYpr2G0v9YRLbqpPw5uVwqQvWxN+mPWZzHDDP+rIFd
TfxTmMGgt0jX0DiTxWtF3FCDWUZZhi9T60LxJYTya15MlqU7EpylYX2i0TgP
W/J2rnsXxje43DSuZOYlS/2/b0/UACQQF5TEqq3X/4F7qwx9O0YVMH6C6ljS
U7hwuqmKtaNtsfhHubcHpauoQfhcXFad7E5lgnPblIb/YDF4EikmYeYC/Heo
29ZYbcpgPv3lnmRfqBU5HSfLYkYI8r2xkh5YPAmZax84tYMrSWeFpwhjYZyN
zk56g2Tohsqj+u3zjbVMekVYFHowArF9ZP0JyldmVrDyz0Uf46pvjR5//m2O
VGFOqBEJMwYAHe1cQA0NFO5yBj9zWZowN9WAfu8/FUIoBBp+tlW7nwJ269F6
TGCga5H4UuNG5WRMbZ+FAnTiEPG2R3W8QK8aeny5azMdCzYS4bmyKRy/vTC6
dMo0NTYXRGmZfJMMakbNzN4jTwK5cfX3TMiOAelNbXNF1wcHZa9GPTJvA9WK
VvN7RoTNCDx6ZPcab8aOINqK7ituZRcfS2VVe+OyxbxZxE5UfKQTKB8maa/3
X3iMkp9uLARNZ5OwrXbtxqRwg39k4713+bZyKAxZaag2lkBnQi4JmeRGVWFt
g2zhP2a+vsCVsg6ARmri5YW/1Logh/oZYeTglNARPj23J8oTuG62oilIocRq
xVE5oREqIdqjti44r7a91vrJ57j+QzK+okCtW5UNlRGubcSY+7a6DbYb+8Wu
gcw9Zc3ZqQeWROgFTcyUMigdxzrPPigE1vefH1JpuCWYlJ39kqmJtixM8v+Y
r/8mhqoCphnS/rPYNzGt1mqAOzMLszJ5QC3bO4R+JAmtF2i+/EpGJwd9r1eu
T0ez8LKHVPZzijWTTCnlApzXP7wjAlj5DUIplSmfzy1033Pebudd3YZ03pCs
g/GaEEE+KOEimOD9BJhQFMnA3Vp3W5XfSAEW3wxf6+W5iFv6/kWsFb2e5oug
Qh7kqp6YuVcYmKYXB48QR3FysIBIDUbpIqMbVsfmClkIev+Z1j2QT58hYVSI
LI87HmfUVsEu+Ic05lPKO/J/Uz/6dbmR/hjkV3vPeOVt4rrVN2mo9qLglAQn
PkCgCMr4Nq4KHl9WRhOp0OoOlykeC9aE2S68b4GbIrA51FyYETskDXngdFNM
KwKhvxGpkr6LWpyMJ4A+1RHS1YQURGH1J7tG94C8EvZuyXzM3WhtsvISZ+sI
lgY9NrCsUg9rKkNEsNHupyXJ2/44SUsrZzas10EcO1ErM6HLqk288nbEjoJO
alFPl9Hiz8HjEwtQ+XLA9pHWdcuvSVI2m9Kv4G2IWpYJdoetJ0FaI1ZohPCb
nj0UeAj/WopxvNU0Uhcr+XLzm8zwT5D6RFQIX7dOPw3HBQ6tWqnDVW9l8StO
zeckfSRwzF+MCTQNf9jDo9PzXPKiJd8rosyOilM0RR111V0vDvqY7GWEyexF
tfmu0Th8LYUqWQ0o5lMEWQ0bELhZwZryptjZSR5FuJPEUHIiq1LC6gbT3Pop
jiNhNIKuqaFUquE1yujX5CfaziK7CyKZexgwH6bwYb+CE/drxTXZGLrLrpug
d6qbfsUdY3pmO/7mUZnMzGDepxs9ImKIq+Pj2dXUAjouioAtp2DMN7BEcwK2
gk5ReHO8JF+zrjB861xieA4Rw0xjWBWtOtbec7fzhiepMWuEw3W6242Bnwki
aiQAS6dt02ALl21iB01fDk4MhU0HDFA0LIUG+MvPvgk1VizWFY3FYyIsro75
O5V+FDpN7hBkC/SdF9YTMiiSjQTe/WzA7vxYAChAT1oV97x8y/JgiAigCleW
KlE4E9gvMA2zkQTUJcjIKBsd5m2LRIIGgwALcMK5cOTFS5yPoWYG0gHmZ15e
otFFjw+8wIicxnymuEv4wfxFTG/Bid7f05kFC/qpJCKcA48pAaCdDDdHl/25
SlyMOPeiaRxyHAUl+RBtVURMQP+onY7tOUvYGqdwHqq4aVMe6AX1CE+UWPnH
F2EIym8UIDlWNjZnUvpPW/o1QgnyyLiUhLS/mbyGJUW5+TchOO9+QgYga1pK
nzm6a1+IAJ2JjB0m2m3qIMMHw6mz/Wc1w5aHlL5i/d9PBLwnGcU0jXW4ETPP
wX6YZ4QOqQGzDQLK3wRHpGKV/C0dclcZ0Ek2hrPmHveaJC242xdgkJAZZv8P
jqGiaQBLpnPnqsVYUlpFJKNpmA76Kh6kQtvKNWXqwQVTm3aQNz52MkdC0pM1
4KkpLI7EARiOH83tQHCGGveFrE9qaHpksJeGwXyzdwzvHiz3Y1xZvYljXQO5
+vZvhTL724OxXSsZ4zZseJfRYzrNuoHIhZ2ti1gsGJ4kjvJcMQPCiHz0igYs
zbJd4j/I0FPPEv0zxqWNFUbYREjahMMq26B1qopg0rdtDN4TiuSvgsfYlOQT
Q2ZgIPCJ2YtRVTlIdnwP1XgmENAe6QUT5c+aTwzYHkBKR6YoGC0zYWfu9E8h
I0WjNFGinF+IggN9aqC76pcE5fCWtswVVWVZnS8jPda0GsUn/da/O4fdBsRU
kLKKRJ9ud4VFDsmmIu0MeB7ZJXt0PE2bQz6J8IR81f36k3deCSiU495PeeMc
fJ7mguB8GojAVeJryBhc+dqFFugp0Q9z2zeInwIiCeD149ovZAgCTTal27eY
lQ6+o0rWfE/usFYrV98yHFRVnutl86GJQRN24rKm/NNKG7p/7PbyCQ/7qhKR
sdveIXzA2/ptfzZUNYj7hBOQjWdbbyj7T/DASjEc6YCcm7XPzKaFHwQ6QJkR
1iL3wP+y7lwZME5IOn3Gf1oQm+9yjOsax1Nn6Y3CSo/EbRqod7n5sxUppVLn
vTrI2PoXW5jZRA5/IAqv3sD7QyDoenHUDtDZH/R7Wa4no2ixkWCM8pgcrIMW
WCmVytaqFfK1Gn90VwWkOFepFkTytxp5MaN3mpay5R0m7YfowSExhU7EcLWl
O1O55vX2B0SaNQbZr7iE5puOhnwjNPCOQVTpMy7K+AWPJwj1GE7BahKb2Ttp
JswWwsW9xpUAVIAXXqbRfGCoNGjR5saqka7Y0zIS2IQi/0cnB5nVelSBrpfn
qkKv2K0fsRDBMw2mN89fAh8u0Deh5EV+1WjRTySUkX9gPbt6cGeJm2QLiPII
GoTDdqbn9m6AbWLv1Z/jj+oKjRJ5VxFEnv0nnJnuGCpEtk3XMpHzGg+SinYI
A/aBzeOTgjgz142C3GzVgOV0nqwn+iVU1BJWlHmejzKsMyEPaTYyDj4LPSMT
nzD07IB1eXjL6NLO9JRBnouqU5Hx70mH/jk0NYiJe4qFKH+jxxFy/9SJYuVX
zku7QYfM3kEFOehHy4DlUrwlsZ9OFQcYWHKVfDNm9LA+1O847AJygBkjkakl
LyUAYuTWbGLuCpQDrDI3qiMx5K76FPHh0bSqMy3d6syIk6UXEI6oCOKgC46X
jKRgEtzvjv92fze8wMJefZbuItVnhU0htb0VOJeFHBO5/prd3V14KDpztr9V
GvBch647RPhqZeBBNT3OxbVMOQQrQKO/aC1mX7vsDz05ATncg/+g8J4iZ49t
yyTLxsKRNFgl1bO9WRA7+6ZOTn1yXDKtJUxyHxqhCrkfYERD/A0u1GI1Xnpt
ghFnhTgeWkd0mlEU5a8tJy3WusYG431WLvvmNDySYZPsfTG/Nn6XXw7UugJs
emExd5RWcJvtTcUj6Ha7Tilqm826nADEphngmidYYuhoM6VopieKQhAWXgAo
FLasoaNPuPJFmuNh/sVpwDk5xNqW61eQ+yINCx7o/C73+X8z8VogNhLPGIw8
caaLCUBl5rTa4yhiOIW22DYkE7rFICQ8D6ENpBuF3w1vG9Loba3R+d6BY+yn
xATbS8mUHmjSSiAGkhaJljif3dnGHT5BKmmZHnhErY2G7xa3/sN8g71x1YHM
v7ZRT/lpK5aG1EMN/Nj2w4orUZubKGnrnLZcy6QKX9jhxyQTlu9qPkzDUEPC
C+FU1MoWXOEKFecMl2k77mnuL2/Qh6iF7Bai4ItBZ6Zer3xNHn79MfnTSPmp
NyvCsznGFArkaHi1R86ciHap3HwqrIsbrkR6s9/HS4Ank/UpQFnuUIVu6Oan
1Ljj71eEpwCG+DzW/Kk3j2cEH6grkG7TnFI7gZu9g/VXfz4XAWiXMLpDVl1O
LMt2p4vkKEsvkGYpzG6wDXHVAn9xcwmtiHK9bQJj1y3qnxbRGDgeGbrRY5To
PPR+WkAbCy9nLGsEaGwdlNlPlsXtIWIwM60g9Wl+BgYZjvTWR0Eq23G5qFvG
SmtCT2iy9JyEELxd6zXoGZj7OSOuMDGgHG0axm6QjOe+OmGWF+ARcQaMBVpw
BG0Rc6TLqkAH3nI59P48dXJiDkqvjSxZfGA5QGJUcO7ldG3qXKUzaRWdWRQS
pVJYiMgLJBAZSr6+cDYsgVoKDZDpvqGi5/AYhlxMPfmuRTuYV0T+lZujYjgT
ZBxTSQfHuLEaCqD21DfxC3BWzpOJ5sVhx68wd2VELYR4zbgoLvVgJkfaqhkn
JmAel2kN0pTcVWhrQ4SEU6APajnWKSNfOJuB1eb0Yy5CC1MrZOyRgJO1qRe1
jsqoUS9cSxVDXMcoIc1CYBnnQG0rhVb1acFq2IO8P1+YlWvs7Sav1QWV++M0
xYOpZ/TcOPuZOTcJCefVFaX6JtYa6a+IOecgMIteqqkCjfShJMBkFPYSG9Nk
GCa8LU+QpzPjuB1UiyqkZZhStggboW7VhnSwQnCJL8iklYUxB7q1LkNcEuhc
HrMdJCYShme62wbR1cr9FPCn3JILg+eqVOh3jEQ6z8hrCDS3kLN/iR8EbS4u
x28OPOqukVeQjyeMdjYJd+epM9d7C6ZN0taLGGNHpPRog5V3sC327uSJj7TC
1F9hNihlXp2PY89p2mNGs83+ZH8HqfO8rLKhAzeWwKmXZ9PBdlOpA1yJ2SNS
zT9kJQMS+l9EJ2DYsMtkR7fs5XB4BwgW78NWmaxkEtCC39wkED6BWK/BUSPY
5mvfyHUmlvG0giMBtmfvaC8qYXaKDwgYXdCjdqHcmgl4fmL8Qqcq+oc1op4l
yfb3yCxkVSTC+sZPUZ0EPKFW0igtIbhhNEgrljtOO6QW7tkiyfLlfqmY5Vja
X66hBh0kASoryAtBBcMTCH6RgTbXirYjCvlLGICxkdEhomSYo/jBkiOhv1Ss
tFcb+nk+W1CUswVMCUy6Zc/xgLo5NF//Is+JdQHA5cj4kzu5Yadrkla57xP0
8tsZev+qr43rLsh6H04z9LX9iQH1YhGKu2WpvlnX9p4EtwLgYetHZCDcQoNE
T//cDtnb6iGI0WfVThQ9qxbrAw3EfFE/H0RVh9qYSzao9mkB/vybXS08JUdz
D4t0qjkalLUJWE2ncIBZ7Zd5euBGv3gfUpf1uHbbZnYepWv0s5ufu3NvE0ri
1++XnX+M43wnaf0KHRvRsPXC6a1eFQB3ua9jMlBRpcCK/xt7CWVFFtVK1/8p
ba9AVkM6TniKoT44z2qA30+npxx6/SIhI9gT3JpFDPgTyh/vg6EjNVF4Cz+y
tOS8t5B+Q5aJ8E58O7KrRxrQhBiMkKdq+m+VELc4fYonIWPnVNdnY32MkeBr
foadeWn1iI3aVvNL1NO17gQdqu0Wjg1SPK7s0tulAI4KZj+JtgmJSi7iHrHd
Y1LYzEeaIbUFNJrsEaviaz9qsqpn233/tHNQxK/lDS60wtJ2nEuCllR+B/P3
fHRacIRX+ahiuWK6g1T54aDChppWuNpgGuEQbujaeDmspWgv0Y9C6Pu/sTIM
p3bb0Mb4FowfjhEg7b5Hhqlb/rRv9xbG/8wucrtvDJrC9li7txhw7XNsCc5z
vFIqYO6vMl3zJ4VKP5Pktu01SGm68m+KGDpuIvYWg4FmzXAcVm18Jt2YDX6p
LV4Vj/C+Grysd1wGI+OEXFvy5HSGSnkXfySk6d3vj1gL0Lm511/nzUN4OiAm
tiTiGZd538FRLiW52eh2o2m6ViX1FO759GEnmotUvK+Rwczh89L/exR7BhpC
43bnoxAZMEXqdg1FcPuBzIpR+x51tYucdc8ODGbm5mZgVDCjdesyeNHhI2TI
QQDKVVazc/3SsF3GHpG+UQ9M0nllWZ5c70pGgpXpzoWIcLrr0UcNn0dyTGkN
TC9obdUYyEFTDCYmn3Hw6rSE2IwjjwAliak7oJ11CYKj3P0MrA+0QB6l2T7d
w/85WWXytiDqZLFmnj0HU6pMrIDlMwg16TTioFX/KFBkT11fGmfnEZHul/hb
1R87+Kvtsu06FxH7+P7pn9lD48iz1X7ERM5Himkp2hyiZToD7nvphQCLUFxO
0OLm5Qt+ObF65WhMgqoSWwjB1bf0Xnu0a8qE9cpfR2SvtM3f24IZOHBfw4As
6cKE8vdkCF3+8EpwzBg99fKjHT1xLQAd8MCUn2es4OTMfO5pbdv/euYIE21h
8RRy19KT5RbEO4cVLuZYWmrENiXKdWvCNBMW4gtsfONVJ5bui2M5xL1z14Ga
gr+7uKNqEmFGACWIxoW4+LcKomZbhixJY2AceQFLVAxDpREcswYbjh7VqQLn
VZrq3axrnXWrOzYmcV8p/1TC3p8RVoO2WHHBxY+4k+BxTSgaURmeFD4q94Wh
QbiDhCMmpxI0HyklkjSqhvgNrEt8dJkCruACYIdEMvDqXQARqT+6CdkS71qJ
QoRnzbZNrmY4niO3/5uHr6e1mnZOBKwrC7wT2uVdMquPhRJeFxHe6uesQi1z
dhCBP12aFxWiR5h7MUWYEf8TKotYFFBn3f1fyUrVdpf+mqCTyEcvSfOl2h7/
ur7bjRnKu7AE6qCA/HiWQT5phHmqpgI2YyZbF6DfuZ4FwWHxq2gbhTyO3Max
8r7wXs53TGyFeiCHNkXZLwxcqbKapHEFFE+hcYlUCvhhnuBrj2eTOCrWWeaV
kjcobam6qoMmIcfxkhsNWsalX4/lvjTKMt99e0+Q56n0BkDJlLemV+R9tPiY
2VNObNmwU6+R7rMkXLqJ6rIHiEJovQM=

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "Fs0mzxxWW3u1nDrkJWuiWcJg9N05rPiXDvI8zzUYttUvzv35r3ZFtKKaqRTR5jmpAZ4wc2UrLeI0ck89858nCqHFdBx8aPbdR0+WnBNhuS/XrodV08Wt78V2otPkmbiS50ZwohSE7w+cseQqgJ8kgxhpG/kV9gq3NsSkdpuipbgRRMtED2IZ7HrTJIBK4TFc/TBNzO5oUucrAbXAKomkxGts0/Oq8TCR4KQZ/NWOPfQg6/D7/sKlE1jE6uU+pNOvApA+jaDAH059YlXwK2a9p7/IT7YhKlRta0L54gxfho6VwfBp1CiaCEbvY8zP4mqEYZ2+p2Y9cG3xMxlvdBu62+4kyVjRHeTxcNmVKz66WZ2VfquDEBYJ7vY9r6puItC2Ks7CzBfOkVkNwiba0leMAfSTDGLdjfqwF8nTnHP8A+7zq6LY9PdC5wDCO91ygbG3E76DA6Ua/0JgCL32t+ay1r7pqT96oqiLiVlQaEv5vmBjwi4ZbgITJMT63AdCTEL7bEgCrUrnYsrEu2IgbUwN+9md6iQVounHZhotXhGziJ6ursHDCF8KPRXj7npSuhK59Uovi4xcjn//wEiVijvrGhVoW+XD/OkP49pxR8lCVOwktDP+aU7Ec8wcw/pGd4HIOeq1dyZS/2CKqWYEf+EVsacU+jlBYbjGxKr3N6XB/qCmmb8MRjHtQ/Cpp2+7/lAbfwC/OMTJc32ooz2fhXLGgI0wOstODkiXF1YrRrEz/v8kbTKbd4znKYztGvGgSkfj2MSGKbpZnQHNqq+GCWDC3qn7G2uxyX4F+4VRr4x9VR7MxEsyWsOK7KuD7gyujm8xrTpHipLzPfzQBackHNBpwxSao5LwJI4eCuoR23MFIwQ226KLIZUVEGE+YLx5QYYOVaLS3UURlzido4vpdcTrnuHxeqQ7493V9II4+rnPYZDHVHJkArtGKibeJUpzeKDAp4RVamu7vsugeZJSfO1NOeAr25jLII41DpL5vrO68z/Ewuqcaze1/pSn2m5IsKme"
`endif