// system_intel_pcie_gts_0_one_lane_pcie_hal_phy_hal_2100_4cpcala.v

// Generated using ACDS version 23.4.1 205

`timescale 1 ps / 1 ps
module system_intel_pcie_gts_0_one_lane_pcie_hal_phy_hal_2100_4cpcala #(
		parameter       ch_xcvrif_l_loopback_mode_atom                     = "LOOPBACK_MODE_DISABLE",
		parameter       ch_flux_l_stmux_rx_demux_sel                       = "SEL_PCIE_PCS",
		parameter       ch_flux_l_stmux_rx_rxword_clk_demux_sel            = "SEL_PCIE_RXWORD_CLK",
		parameter       ch_flux_l_stmux_tx_txword_clk_demux_sel            = "SEL_PCIE_TXWORD_CLK",
		parameter       ch_flux_l_stmux_tx_mux_sel                         = "SEL_PCIE_PCS",
		parameter       ch_flux_l_stmux_tx_txword_clk_mux_sel              = "SEL_UX_OCK_PMA_CLK",
		parameter       ch_xcvrif_rx_ch_clk_static_mux                     = "SEL_UNUSED",
		parameter       ch_xcvrif_tx_ch_clk_static_mux                     = "SEL_UNUSED",
		parameter       ch_flux_l_tx_bond_size_atom                        = "TX_BOND_SIZE_X4",
		parameter       ch_l_xcvr_tx_bond_size_atom                        = "TX_BOND_SIZE_X4",
		parameter       ch_xcvrif_l_tx_bond_size_atom                      = "TX_BOND_SIZE_UNUSED",
		parameter       ch_xcvrif_l_rx_bond_size_atom                      = "RX_BOND_SIZE_UNUSED",
		parameter       ch_clkrx_refclk_cssm_fw_control_atom               = "CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch_clkrx_refclk_sector_specifies_refclk_ready_atom = "CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch_local_refclk_cssm_fw_control_atom               = "LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE",
		parameter       ch_local_refclk_sector_specifies_refclk_ready_atom = "LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE",
		parameter       ch_l_tx_pll_postdiv_sel_atom                       = "TX_PLL_POSTDIV_SEL_SYNTH2",
		parameter       ch_l_tx_pll_bw_sel_atom                            = "TX_PLL_BW_SEL_LOW",
		parameter[35:0] ch_l_tx_pll_f_out_hz_atom                          = 36'b000111011100110101100101000000000000,
		parameter[35:0] ch_l_tx_pll_f_vco_hz_atom                          = 36'b001001010100000010111110010000000000,
		parameter[35:0] ch_l_tx_pll_f_pfd_hz_atom                          = 36'b000000000101111101011110000100000000,
		parameter[35:0] ch_l_tx_pll_f_ref_hz_atom                          = 36'b000000000101111101011110000100000000,
		parameter[21:0] ch_l_tx_pll_k_counter_atom                         = 22'b0000000000000000000000,
		parameter[5:0]  ch_l_tx_pll_l_counter_atom                         = 6'b000001,
		parameter[8:0]  ch_l_tx_pll_m_counter_atom                         = 9'b001100100,
		parameter[5:0]  ch_l_tx_pll_n_counter_atom                         = 6'b000001,
		parameter[1:0]  ch_l_tx_pll_fb_counter_atom                        = 2'b01,
		parameter[35:0] ch_l_tx_postdiv_cdr_refclk_hz_atom                 = 36'b000000000000000000000000000000000000,
		parameter[7:0]  ch_l_tx_postdiv_cdr_refclk_divider_atom            = 8'b00001100,
		parameter[7:0]  ch_l_tx_synthdiv_out_divider_atom                  = 8'b00001100,
		parameter[35:0] ch_l_tx_synthdiv_out_hz_atom                       = 36'b000000000000000000000000000000000000,
		parameter[35:0] ch_l_xcvr_cdr_f_out_hz_atom                        = 36'b000111011100110101100101000000000000,
		parameter[35:0] ch_l_xcvr_cdr_f_vco_hz_atom                        = 36'b001001010100000010111110010000000000,
		parameter[35:0] ch_l_xcvr_cdr_f_pfd_hz_atom                        = 36'b000000000101111101011110000100000000,
		parameter[35:0] ch_l_xcvr_cdr_f_ref_hz_atom                        = 36'b000000000101111101011110000100000000,
		parameter[5:0]  ch_l_cdr_l_counter_atom                            = 6'b000001,
		parameter[8:0]  ch_l_cdr_m_counter_atom                            = 9'b000110010,
		parameter[5:0]  ch_l_cdr_n_counter_atom                            = 6'b000001,
		parameter       ch_l_xcvr_tx_preloaded_hardware_configs_atom       = "TX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch_l_xcvr_tx_protocol_hint_atom                    = "TX_PROTOCOL_HINT_DISABLED",
		parameter[36:0] ch_l_xcvr_tx_datarate_bps_atom                     = 37'b0001110111001101011001010000000000000,
		parameter       ch_l_xcvr_tx_prbs_gen_en_atom                      = "TX_PRBS_GEN_EN_DISABLE",
		parameter[3:0]  ch_l_xcvr_tx_prbs_pattern_atom                     = 4'b1001,
		parameter       ch_l_xcvr_tx_user_clk_only_mode_atom               = "TX_USER_CLK_ONLY_MODE_DISABLE",
		parameter       ch_l_xcvr_tx_width_atom                            = "TX_WIDTH_X16",
		parameter[35:0] ch_l_xcvr_tx_word_clk_hz_atom                      = 36'b000000111011100110101100101000000000,
		parameter       ch_l_xcvr_tx_dl_enable_atom                        = "TX_DL_ENABLE_DISABLE",
		parameter       ch_l_xcvr_rx_preloaded_hardware_configs_atom       = "RX_PRELOADED_HARDWARE_CONFIGS_PCIE",
		parameter       ch_l_xcvr_rx_protocol_hint_atom                    = "RX_PROTOCOL_HINT_DISABLED",
		parameter[36:0] ch_l_xcvr_rx_datarate_bps_atom                     = 37'b0001110111001101011001010000000000000,
		parameter       ch_l_xcvr_rx_prbs_monitor_en_atom                  = "RX_PRBS_MONITOR_EN_DISABLE",
		parameter[3:0]  ch_l_xcvr_rx_prbs_pattern_atom                     = 4'b0000,
		parameter       ch_l_xcvr_rx_width_atom                            = "RX_WIDTH_X16",
		parameter       ch_l_xcvr_rx_force_cdr_ltr_atom                    = "TRUE",
		parameter       ch_l_xcvr_rx_adaptation_mode_atom                  = "RX_ADAPTATION_MODE_UX_NATIVE_ADAPTATION",
		parameter[35:0] ch_l_xcvr_rx_word_clk_hz_atom                      = 36'b000000111011100110101100101000000000,
		parameter       ch_l_xcvr_rx_dl_enable_atom                        = "RX_DL_ENABLE_ENABLE",
		parameter       ch_l_rx_postdiv_clk_en_atom                        = "RX_POSTDIV_CLK_EN_ENABLE",
		parameter[7:0]  ch_l_rx_postdiv_clk_divider_atom                   = 8'b00001100,
		parameter[7:0]  ch_l_tx_postdiv_clk_divider_atom                   = 8'b10001001,
		parameter       ch_l_tx_pll_refclk_select_atom                     = "TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter       ch_l_loopback_mode_atom                            = "LOOPBACK_MODE_DISABLED",
		parameter       ch_flux_l_flux_mode_atom                           = "FLUX_MODE_FLUX_MODE_BYPASS",
		parameter       ch_flux_l_rx_protocol_hint_atom                    = "RX_PROTOCOL_HINT_DISABLED",
		parameter       ch_flux_l_tx_dl_enable_atom                        = "TX_DL_ENABLE_DISABLE",
		parameter       ch_flux_l_rx_dl_enable_atom                        = "RX_DL_ENABLE_DISABLE",
		parameter       ch_xcvrif_l_tx_dl_enable_atom                      = "TX_DL_ENABLE_DISABLE",
		parameter       ch_xcvrif_l_rx_dl_enable_atom                      = "RX_DL_ENABLE_DISABLE",
		parameter       ch_xcvrif_l_tx_fifo_mode_atom                      = "TX_FIFO_MODE_DISABLED",
		parameter       ch_xcvrif_l_rx_fifo_mode_atom                      = "RX_FIFO_MODE_DISABLED",
		parameter       ch_l_xcvr_tx_en_atom                               = "TRUE",
		parameter       ch_l_xcvr_rx_en_atom                               = "TRUE",
		parameter       ch_l_duplex_mode_atom                              = "DUPLEX_MODE_DUPLEX",
		parameter       ch_xcvrif_l_tx_en_atom                             = "FALSE",
		parameter       ch_xcvrif_l_rx_en_atom                             = "FALSE",
		parameter       ch_xcvrif_l_duplex_mode_atom                       = "DUPLEX_MODE_RX_ONLY_SIMPLEX",
		parameter       ch_flux_l_rx_fec_type_used_atom                    = "RX_FEC_TYPE_USED_NONE",
		parameter       ch_l_sim_mode_atom                                 = "SIM_MODE_DISABLE",
		parameter       ch_flux_l_rx_sim_mode_atom                         = "RX_SIM_MODE_DISABLE",
		parameter       ch_flux_l_tx_sim_mode_atom                         = "TX_SIM_MODE_DISABLE",
		parameter       ch_flux_l_dr_enabled_atom                          = "DR_ENABLED_DR_DISABLED",
		parameter       ch_xcvrif_l_sup_mode_atom                          = "SUP_MODE_USER_MODE",
		parameter       ch_xcvrif_l_sim_mode_atom                          = "SIM_MODE_ENABLE",
		parameter       ch_xcvrif_l_dr_enabled_atom                        = "DR_ENABLED_DR_DISABLED",
		parameter       ch_l_xcvr_tx_spread_spectrum_en_atom               = "TX_SPREAD_SPECTRUM_EN_ENABLE",
		parameter[35:0] ch_l_rx_postdiv_clk_hz_atom                        = 36'b000000000000000000000000000000000000,
		parameter       ch_l_rx_postdiv_clk_fractional_en_atom             = "RX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE",
		parameter       ch_l_cdr_refclk_select_atom                        = "CDR_REFCLK_SELECT_GLOBAL_REFCLK0",
		parameter[35:0] ch_l_tx_postdiv_clk_hz_atom                        = 36'b000000000000000000000000000000000000,
		parameter       ch_l_tx_postdiv_clk_fractional_en_atom             = "TX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE",
		parameter       ch_flux_l_lc_postdiv_sel_atom                      = "LC_POSTDIV_SEL_SYNTH2",
		parameter       ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom        = "TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom        = "TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK",
		parameter       ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom        = "RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom        = "RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD",
		parameter       ch_xcvrif_l_tx_gb_width_atom                       = "TX_GB_WIDTH_DISABLED",
		parameter       ch_xcvrif_l_rx_gb_width_atom                       = "RX_GB_WIDTH_DISABLED",
		parameter       ch_xcvrif_l_tx_dynamic_mux_atom                    = "TX_DYNAMIC_MUX_UNUSED",
		parameter       ch_xcvrif_l_tx_word_clk_dynamic_mux_atom           = "TX_WORD_CLK_DYNAMIC_MUX_X4",
		parameter       ch_xcvrif_l_rx_word_clk_dynamic_mux_atom           = "RX_WORD_CLK_DYNAMIC_MUX_UNUSED",
		parameter       ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom         = "TX_FIFO_RD_EN_DYNAMIC_MUX_X4",
		parameter       ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom         = "RX_FIFO_RD_EN_DYNAMIC_MUX_UNUSED",
		parameter       ch_xcvrif_l_tx_rst_dynamic_mux_atom                = "TX_RST_DYNAMIC_MUX_X4",
		parameter       ch_l_clk_debug_select_0_enable_atom                = "CLK_DEBUG_SELECT_0_ENABLE_DISABLE",
		parameter       ch_l_clk_debug_select_0_setting_atom               = "CLK_DEBUG_SELECT_0_SETTING_DISABLED",
		parameter       ch_l_clk_debug_select_1_enable_atom                = "CLK_DEBUG_SELECT_1_ENABLE_DISABLE",
		parameter       ch_l_clk_debug_select_1_setting_atom               = "CLK_DEBUG_SELECT_1_SETTING_DISABLED",
		parameter[5:0]  ch_l_xcvr_tx_eq_main_tap_atom                      = 6'b000000,
		parameter[4:0]  ch_l_xcvr_tx_eq_post_tap_1_atom                    = 5'b00000,
		parameter[4:0]  ch_l_xcvr_tx_eq_pre_tap_1_atom                     = 5'b00000,
		parameter[2:0]  ch_l_xcvr_tx_eq_pre_tap_2_atom                     = 3'b000,
		parameter[7:0]  ch_l_tx_pll_feed_forward_gain_atom                 = 8'b01000011,
		parameter       ch_l_xcvr_rx_termination_mode_atom                 = "RX_TERMINATION_MODE_GROUNDED",
		parameter       ch_l_xcvr_rx_onchip_termination_setting_atom       = "RX_ONCHIP_TERMINATION_SETTING_R_1",
		parameter[6:0]  ch_l_xcvr_rx_eq_vga_gain_atom                      = 7'b0100000,
		parameter[5:0]  ch_l_xcvr_x_eq_hf_boost_atom                       = 6'b100000,
		parameter[5:0]  ch_l_xcvr_rx_eq_dfe_tap_1_atom                     = 6'b000000,
		parameter       ch_l_xcvr_rx_external_couple_type_atom             = "RX_EXTERNAL_COUPLE_TYPE_AC",
		parameter       ch_l_xcvr_tx_bonding_category_atom                 = "TX_BONDING_CATEGORY_BONDING_FOLLOWER",
		parameter       ch_l_xcvr_tx_master_pll_mode_atom                  = "TX_MASTER_PLL_MODE_DISABLED",
		parameter       ch_l_xcvr_rx_cdrdivout_en_atom                     = "RX_CDRDIVOUT_EN_DISABLE",
		parameter       ch_xcvrif_l_tx_bonding_mode_atom                   = "TX_BONDING_MODE_UNUSED",
		parameter       ch_xcvrif_l_rx_bonding_mode_atom                   = "RX_BONDING_MODE_UNUSED",
		parameter       ch_flux_l_sequencer_reg_en_atom                    = "SEQUENCER_REG_EN_DISABLE",
		parameter       ch_l_speed_grade_atom                              = "SPEED_GRADE_DASH_1",
		parameter       ch_usb_mode_atom                                   = "USB_MODE_DISABLED",
		parameter       ch_pcie_mode_atom                                  = "PCIE_MODE_GEN4",
		parameter[35:0] ch_l_ick_tx_word_clk_hz_atom                       = 36'b100101011100000111110010100001110010,
		parameter[35:0] ch_l_pcs_ref_clk_hz_atom                           = 36'b101001111010110110010111101111110101,
		parameter[35:0] ch_l_lane_common_ref_clk_hz_atom                   = 36'b111110010011110101111111101000101001,
		parameter       ch_rx_invert_pin_atom                              = "RX_INVERT_PIN_DISABLE",
		parameter       ch_tx_invert_pin_atom                              = "TX_INVERT_PIN_DISABLE",
		parameter[17:0] ch_rx_dl_rx_lat_bit_for_async_atom                 = 18'b111110100110100101,
		parameter       ch_rx_dl_rxbit_cntr_pma_atom                       = "RX_DL_RXBIT_CNTR_PMA_DISABLE",
		parameter[17:0] ch_rx_dl_rxbit_rollover_atom                       = 18'b001001111001000101,
		parameter[35:0] ch_eth_rx_clk_hz_atom                              = 36'b000000000000000000000000000000000000,
		parameter[35:0] ch_eth_tx_clk_hz_atom                              = 36'b000000000000000000000000000000000000
	) (
		output wire         oflux_xoa_tx_n_l0_ux,              //              oflux_xoa_tx_n_l0_ux.data,          Stats Snapshot
		output wire         oflux_xoa_tx_p_l0_ux,              //              oflux_xoa_tx_p_l0_ux.data,          RX PFC
		input  wire         iflux_xia_rx_n_l0_ux,              //              iflux_xia_rx_n_l0_ux.data,          CSR access address
		input  wire         iflux_xia_rx_p_l0_ux,              //              iflux_xia_rx_p_l0_ux.data,          RX error bits asserted on the EOP cycle
		input  wire [79:0]  i_ss_async_pldif,                  //                       asyncdata_0.data,          Stats Snapshot
		output wire [49:0]  o_ss_async_pldif,                  //                       asyncdata_1.data,          RX PFC
		input  wire [79:0]  i_ss_async_pldif_pcie_mux,         //                       asyncdata_2.data,          CSR access address
		input  wire [19:0]  i_lavmm_addr,                      //                          reconfig.address,       RX error bits asserted on the EOP cycle
		input  wire [3:0]   i_lavmm_be,                        //                                  .byteenable,    Stats Snapshot
		input  wire         i_lavmm_read,                      //                                  .read,          CSR access address
		input  wire [31:0]  i_lavmm_wdata,                     //                                  .writedata,     RX error bits asserted on the EOP cycle
		input  wire         i_lavmm_write,                     //                                  .write,         Stats Snapshot
		output wire [31:0]  o_lavmm_rdata,                     //                                  .readdata,      RX PFC
		output wire         o_lavmm_rdata_valid,               //                                  .readdatavalid, CSR access address
		output wire         o_lavmm_waitreq,                   //                                  .waitrequest
		input  wire         i_lavmm_clk,                       //                      reconfig_clk.clk,           RX PFC
		input  wire         i_lavmm_rstn,                      //                      reconfig_rst.reset,         RX error bits asserted on the EOP cycle
		input  wire         i_ft_rx_sclk_sync_ch,              //              i_ft_rx_sclk_sync_ch.clk,           Stats Snapshot
		input  wire         i_ft_tx_sclk_sync_ch,              //              i_ft_tx_sclk_sync_ch.clk,           RX PFC
		output wire         o_ft_rx_async_pulse_ch,            //            o_ft_rx_async_pulse_ch.clk,           CSR access address
		output wire         o_ft_tx_async_pulse_ch,            //            o_ft_tx_async_pulse_ch.clk
		output wire         o_rxcdrlock2dataa,                 //                 o_rxcdrlock2dataa.lockdata,      Stats Snapshot
		input  wire         i_rst_ux_rx_sfrz,                  //                  i_rst_ux_rx_sfrz.data
		output wire         o_rst_flux0_cpi_cmn_busy,          //          o_rst_flux0_cpi_cmn_busy.busy,          CSR access address
		output wire         o_rst_oflux_rx_srds_rdy,           //           o_rst_oflux_rx_srds_rdy.ready
		output wire         o_rst_ux_all_synthlockstatus,      //      o_rst_ux_all_synthlockstatus.status
		output wire         o_rst_ux_rxcdrlockstatus,          //          o_rst_ux_rxcdrlockstatus.rxstatus
		output wire         o_ux_tx_ch_ptr_smpl,               //               o_ux_tx_ch_ptr_smpl.sample
		input  wire         i_ick_sclk_tx,                     //                     i_ick_sclk_tx.clk
		input  wire         i_ick_sclk_rx,                     //                     i_ick_sclk_rx.clk
		input  wire         i_rst_pld_ux_tx_pma_rst_n,         //         i_rst_pld_ux_tx_pma_rst_n.reset
		input  wire         i_rst_pld_ux_rx_pma_rst_n,         //         i_rst_pld_ux_rx_pma_rst_n.reset
		output wire [31:0]  o_ch_lavmm_xcvrif_rdata,           //                     reconfig_xcvr.readdata
		output wire         o_ch_lavmm_xcvrif_rdata_valid,     //                                  .readdatavalid
		output wire         o_ch_lavmm_xcvrif_waitreq,         //                                  .waitrequest
		input  wire [19:0]  i_ch_lavmm_xcvrif_addr,            //                                  .address
		input  wire [3:0]   i_ch_lavmm_xcvrif_be,              //                                  .byteenable
		input  wire         i_ch_lavmm_xcvrif_read,            //                                  .read
		input  wire [31:0]  i_ch_lavmm_xcvrif_wdata,           //                                  .writedata,     RX error bits asserted on the EOP cycle
		input  wire         i_ch_lavmm_xcvrif_write,           //                                  .write,         RX error bits asserted on the EOP cycle
		input  wire         i_ch_lavmm_xcvrif_clk,             //                 reconfig_clk_xcvr.clk
		input  wire         i_ch_lavmm_xcvrif_rstn,            //                 reconfig_rst_xcvr.reset,         RX error bits asserted on the EOP cycle
		output wire         o_rx_latency_pulse,                //                o_rx_latency_pulse.clk,           RX error bits asserted on the EOP cycle
		output wire         o_tx_latency_pulse,                //                o_tx_latency_pulse.clk,           RX error bits asserted on the EOP cycle
		input  wire [6:0]   i_ch_eth_xcvrif_tx_async,          //                       asyncdata_3.data,          RX error bits asserted on the EOP cycle
		input  wire         i_ch_eth_xcvrif_tx_direct,         //                       asyncdata_4.data
		output wire [13:0]  o_ch_eth_xcvrif_rx_async,          //                       asyncdata_5.data
		output wire         o_ch_eth_xcvrif_rx_direct,         //                       asyncdata_6.data
		input  wire         i_rstxcvrif_xcvrif_signal_ok,      //      i_rstxcvrif_xcvrif_signal_ok.data
		input  wire         i_rstxcvrif_rx_xcvrif_sfrz_n,      //      i_rstxcvrif_rx_xcvrif_sfrz_n.data
		input  wire         i_rstxcvrif_xcvrif_rx_rst_n,       //       i_rstxcvrif_xcvrif_rx_rst_n.data
		input  wire         i_rstxcvrif_tx_xcvrif_sfrz_n,      //      i_rstxcvrif_tx_xcvrif_sfrz_n.data
		input  wire         i_rstxcvrif_xcvrif_tx_rst_n,       //       i_rstxcvrif_xcvrif_tx_rst_n.data
		output wire         o_pma_rx_sf,                       //                       o_pma_rx_sf.data
		input  wire [42:0]  i_xcvrif_tx_mux_data,              //              i_xcvrif_tx_mux_data.data
		output wire [42:0]  o_rx_data,                         //                         o_rx_data.data
		output wire [1:0]   o_tx_source_sel,                   //                   o_tx_source_sel.data
		output wire [2:0]   o_rx_fifo_en_sel,                  //                  o_rx_fifo_en_sel.data
		output wire [2:0]   o_tx_rst_source_sel,               //               o_tx_rst_source_sel.data
		input  wire         i_ch_xcvrif_rx_fifo_rd_en,         //         i_ch_xcvrif_rx_fifo_rd_en.data
		output wire         o_ch_xcvrif_rx_fifo_rd_en,         //         o_ch_xcvrif_rx_fifo_rd_en.data
		input  wire         i_ch_xcvrif_tx_fifo_rd_en,         //         i_ch_xcvrif_tx_fifo_rd_en.data
		output wire         o_ch_xcvrif_tx_fifo_rd_en,         //         o_ch_xcvrif_tx_fifo_rd_en.data
		output wire [1:0]   o_ux_rxuser1_sel,                  //                  o_ux_rxuser1_sel.data
		output wire [1:0]   o_ux_rxuser2_sel,                  //                  o_ux_rxuser2_sel.data
		output wire [1:0]   o_ux_txuser1_sel,                  //                  o_ux_txuser1_sel.data
		output wire [1:0]   o_ux_txuser2_sel,                  //                  o_ux_txuser2_sel.data
		output wire         o_pcs_rxpostdiv,                   //                   o_pcs_rxpostdiv.data
		output wire         o_pcs_rxword,                      //                      o_pcs_rxword.data
		output wire         o_ux_txlc_clk,                     //                     o_ux_txlc_clk.clk
		output wire [2:0]   o_tx_xcvr_wordclk_sel,             //             o_tx_xcvr_wordclk_sel.data
		output wire [1:0]   o_rx_xcvr_wordclk_sel,             //             o_rx_xcvr_wordclk_sel.data
		input  wire         i_eth_rx_ch_clk,                   //                   i_eth_rx_ch_clk.clk
		input  wire [767:0] uxwrap_bus_in,                     //                     uxwrap_bus_in.data
		output wire [703:0] uxwrap_bus_out,                    //                    uxwrap_bus_out.data
		output wire [19:0]  o_lavmm_addr,                      //               reconfig_phy_shared.address
		output wire [3:0]   o_lavmm_be,                        //                                  .byteenable
		output wire         o_lavmm_read,                      //                                  .read
		output wire [31:0]  o_lavmm_wdata,                     //                                  .writedata
		output wire         o_lavmm_write,                     //                                  .write
		input  wire [31:0]  i_lavmm_rdata,                     //                                  .readdata
		input  wire         i_lavmm_rdata_valid,               //                                  .readdatavalid
		input  wire         i_lavmm_waitreq,                   //                                  .waitrequest
		output wire         o_lavmm_clk,                       //           reconfig_clk_phy_shared.clk
		output wire         o_lavmm_rstn,                      //           reconfig_rst_phy_shared.reset
		output wire         o_sclk_return_sel_rx,              //              o_sclk_return_sel_rx.data
		output wire         o_sclk_return_sel_tx,              //              o_sclk_return_sel_tx.data
		output wire         o_ick_sclk_rx,                     //                     o_ick_sclk_rx.clk
		input  wire [4:0]   i_sync_common_control,             //             i_sync_common_control.data
		output wire         o_ft_rx_sclk_sync_ch,              //              o_ft_rx_sclk_sync_ch.data
		output wire         o_ft_tx_sclk_sync_ch,              //              o_ft_tx_sclk_sync_ch.data
		output wire         o_rst_ux_rx_pma_rst_n,             //             o_rst_ux_rx_pma_rst_n.reset
		output wire         o_rst_ux_tx_pma_rst_n,             //             o_rst_ux_tx_pma_rst_n.reset
		output wire         o_ick_pcs_txword,                  //                  o_ick_pcs_txword.data
		output wire         o_tx_dl_ch_bit,                    //                    o_tx_dl_ch_bit.data
		input  wire         i_dat_pcs_measlatbit,              //              i_dat_pcs_measlatbit.data
		input  wire         i_ft_rx_async_pulse_ch,            //            i_ft_rx_async_pulse_ch.data
		input  wire         i_ft_tx_async_pulse_ch,            //            i_ft_tx_async_pulse_ch.data
		input  wire         i_rx_dl_ch_bit,                    //                    i_rx_dl_ch_bit.data
		input  wire [1:0]   i_ux_rxuser1_sel,                  //                  i_ux_rxuser1_sel.data
		input  wire [1:0]   i_ux_rxuser2_sel,                  //                  i_ux_rxuser2_sel.data
		input  wire [1:0]   i_ux_txuser1_sel,                  //                  i_ux_txuser1_sel.data
		input  wire [1:0]   i_ux_txuser2_sel,                  //                  i_ux_txuser2_sel.data
		output wire         o_octl_pcs_txstatus_a,             //             o_octl_pcs_txstatus_a.data
		input  wire         i_ictl_pcs_txenable_a,             //             i_ictl_pcs_txenable_a.data
		input  wire [124:0] i_sync_cfg_data,                   //                   i_sync_cfg_data.data
		input  wire [249:0] i_sync_interface_control,          //          i_sync_interface_control.data
		output wire [79:0]  o_tx_data,                         //                         o_tx_data.data
		input  wire [79:0]  i_rx_data,                         //                         i_rx_data.data
		output wire [319:0] o_sm_flux_ingress,                 //                 o_sm_flux_ingress.data
		input  wire [256:0] i_sm_flux_egress,                  //                  i_sm_flux_egress.data
		input  wire         i_flux_cpi_int,                    //                    i_flux_cpi_int.data
		input  wire         i_flux_int,                        //                        i_flux_int.data
		input  wire         i_oflux_octl_pcs_txptr_smpl_lane,  //  i_oflux_octl_pcs_txptr_smpl_lane.data
		output wire         o_ick_sclk_tx,                     //                     o_ick_sclk_tx.clk
		input  wire         i_flux_srds_rdy,                   //                   i_flux_srds_rdy.data
		input  wire         i_pcs_rxword,                      //                      i_pcs_rxword.data
		input  wire         i_pcs_rxpostdiv,                   //                   i_pcs_rxpostdiv.data
		input  wire         i_ock_pcs_txword,                  //                  i_ock_pcs_txword.data
		output wire         o_dat_pcs_measlatrndtripbit,       //       o_dat_pcs_measlatrndtripbit.data
		output wire         o_ock_pcs_cdrfbclk,                //                o_ock_pcs_cdrfbclk.data
		output wire         o_ock_pcs_ref,                     //                     o_ock_pcs_ref.data
		output wire [39:0]  o_pcie_pcs,                        //                        o_pcie_pcs.data
		input  wire [39:0]  i_pcie_pcs,                        //                        i_pcie_pcs.data
		input  wire         i_sel_rxword_clk,                  //                  i_sel_rxword_clk.clk
		input  wire         i_xcvr_txword_clk,                 //                 i_xcvr_txword_clk.clk
		output wire         o_pcie_rxword_clk,                 //                 o_pcie_rxword_clk.clk
		output wire         o_eth_rxword_clk,                  //                  o_eth_rxword_clk.clk
		output wire         o_pcie_txword_clk,                 //                 o_pcie_txword_clk.clk
		output wire         o_eth_txword_clk,                  //                  o_eth_txword_clk.clk
		output wire         o_ock_pcs_txword,                  //                  o_ock_pcs_txword.clk
		output wire         o_eth_rx_ch_clk,                   //                   o_eth_rx_ch_clk.clk
		output wire         o_eth_tx_ch_clk,                   //                   o_eth_tx_ch_clk.clk
		input  wire [5:0]   ioack_ref_left_p_ux_bidir_in,      //      ioack_ref_left_p_ux_bidir_in.data
		input  wire         ioack_hsref_left_p_ux_bidir_in,    //    ioack_hsref_left_p_ux_bidir_in.clk
		input  wire         ioack_cdrdiv_left_ux_bidir_in,     //     ioack_cdrdiv_left_ux_bidir_in.clk
		input  wire         ioack_synthdiv1_left_ux_bidir_in,  //  ioack_synthdiv1_left_ux_bidir_in.clk
		input  wire         ioack_synthdiv2_left_ux_bidir_in,  //  ioack_synthdiv2_left_ux_bidir_in.clk
		output wire         ioack_cdrdiv_left_ux_bidir_out,    //    ioack_cdrdiv_left_ux_bidir_out.clk
		output wire         ioack_synthdiv1_left_ux_bidir_out, // ioack_synthdiv1_left_ux_bidir_out.clk
		output wire         ioack_synthdiv2_left_ux_bidir_out, // ioack_synthdiv2_left_ux_bidir_out.clk
		output wire [13:0]  o_rxeq_best_eye_vala,              //              o_rxeq_best_eye_vala.data
		output wire         o_rxeq_donea,                      //                      o_rxeq_donea.data
		output wire         o_rxmargin_nacka,                  //                  o_rxmargin_nacka.data
		output wire         o_rxmargin_statusa,                //                o_rxmargin_statusa.data
		output wire         o_rxsignaldetect_lfpsa,            //            o_rxsignaldetect_lfpsa.data
		output wire         o_rxsignaldetecta,                 //                 o_rxsignaldetecta.data
		output wire [1:0]   o_rxmargin_status_gray,            //            o_rxmargin_status_gray.data
		output wire         o_rxstatusa,                       //                       o_rxstatusa.data
		output wire         o_synthlcfast_postdiv,             //             o_synthlcfast_postdiv.data
		output wire         o_synthlcmed_postdiv,              //              o_synthlcmed_postdiv.data
		output wire         o_synthlcslow_postdiv,             //             o_synthlcslow_postdiv.data
		output wire         o_txdetectrx_acka,                 //                 o_txdetectrx_acka.data
		output wire         o_txdetectrx_statct,               //               o_txdetectrx_statct.data
		output wire         o_txstatusa,                       //                       o_txstatusa.data
		input  wire         i_quartus_flux_s_to_ingress,       //       i_quartus_flux_s_to_ingress.data
		input  wire         i_pcs_pipe_rstn,                   //                   i_pcs_pipe_rstn.data
		input  wire         i_ux_ock_pma_clk,                  //                  i_ux_ock_pma_clk.data
		input  wire         i_lfps_ennt,                       //                       i_lfps_ennt.data
		input  wire [1:0]   i_pcie_l1ctrla,                    //                    i_pcie_l1ctrla.data
		input  wire         i_pma_cmn_ctrl,                    //                    i_pma_cmn_ctrl.data
		input  wire         i_pma_ctrl,                        //                        i_pma_ctrl.data
		input  wire         i_pcie_pcs_rx_rst,                 //                 i_pcie_pcs_rx_rst.data
		input  wire         i_pcie_pcs_tx_rst,                 //                 i_pcie_pcs_tx_rst.data
		input  wire         i_rxeiosdetectstata,               //               i_rxeiosdetectstata.data
		input  wire [2:0]   i_rxeq_precal_code_selnt,          //          i_rxeq_precal_code_selnt.data
		input  wire         i_rxeq_starta,                     //                     i_rxeq_starta.data
		input  wire         i_rxeq_static_ena,                 //                 i_rxeq_static_ena.data
		input  wire         i_rxmargin_direction_nt,           //           i_rxmargin_direction_nt.data
		input  wire         i_rxmargin_mode_nt,                //                i_rxmargin_mode_nt.data
		input  wire         i_rxmargin_offset_change_a,        //        i_rxmargin_offset_change_a.data
		input  wire [6:0]   i_rxmargin_offset_nt,              //              i_rxmargin_offset_nt.data
		input  wire         i_rxmargin_start_a,                //                i_rxmargin_start_a.data
		input  wire [2:0]   i_rxpstate,                        //                        i_rxpstate.data
		input  wire [3:0]   i_rxrate,                          //                          i_rxrate.data
		input  wire         i_rxterm_hiz_ena,                  //                  i_rxterm_hiz_ena.data
		input  wire [2:0]   i_rxwidth,                         //                         i_rxwidth.data
		input  wire         i_tstbus_lane,                     //                     i_tstbus_lane.data
		input  wire         i_txbeacona,                       //                       i_txbeacona.data
		input  wire [2:0]   i_txclkdivrate,                    //                    i_txclkdivrate.data
		input  wire         i_txdetectrx_reqa,                 //                 i_txdetectrx_reqa.data
		input  wire [5:0]   i_txdrv_levn,                      //                      i_txdrv_levn.data
		input  wire [4:0]   i_txdrv_levnm1,                    //                    i_txdrv_levnm1.data
		input  wire [2:0]   i_txdrv_levnm2,                    //                    i_txdrv_levnm2.data
		input  wire [4:0]   i_txdrv_levnp1,                    //                    i_txdrv_levnp1.data
		input  wire [3:0]   i_txdrv_slew,                      //                      i_txdrv_slew.data
		input  wire [3:0]   i_txelecidle,                      //                      i_txelecidle.data
		input  wire [2:0]   i_txpstate,                        //                        i_txpstate.data
		input  wire [3:0]   i_txrate,                          //                          i_txrate.data
		input  wire [2:0]   i_txwidth,                         //                         i_txwidth.data
		input  wire         i_rstxcvrif_xcvrif_tx_rd_rst_n,    //    i_rstxcvrif_xcvrif_tx_rd_rst_n.data
		input  wire         i_rstxcvrif_xcvrif_tx_wr_rst_n,    //    i_rstxcvrif_xcvrif_tx_wr_rst_n.data
		output wire         o_tx_rst_rd_sync_rst_n,            //            o_tx_rst_rd_sync_rst_n.data
		output wire         o_tx_rst_wr_sync_rst_n             //            o_tx_rst_wr_sync_rst_n.data
	);

	generate
		// If any of the display statements (or deliberately broken
		// instantiations) within this generate block triggers then this module
		// has been instantiated this module with a set of parameters different
		// from those it was generated for.  This will usually result in a
		// non-functioning system.
		if (ch_xcvrif_l_loopback_mode_atom != "LOOPBACK_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_stmux_rx_demux_sel != "SEL_PCIE_PCS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_stmux_rx_demux_sel_check ( .error(1'b1) );
		end
		if (ch_flux_l_stmux_rx_rxword_clk_demux_sel != "SEL_PCIE_RXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_stmux_rx_rxword_clk_demux_sel_check ( .error(1'b1) );
		end
		if (ch_flux_l_stmux_tx_txword_clk_demux_sel != "SEL_PCIE_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_stmux_tx_txword_clk_demux_sel_check ( .error(1'b1) );
		end
		if (ch_flux_l_stmux_tx_mux_sel != "SEL_PCIE_PCS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_stmux_tx_mux_sel_check ( .error(1'b1) );
		end
		if (ch_flux_l_stmux_tx_txword_clk_mux_sel != "SEL_UX_OCK_PMA_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_stmux_tx_txword_clk_mux_sel_check ( .error(1'b1) );
		end
		if (ch_xcvrif_rx_ch_clk_static_mux != "SEL_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_rx_ch_clk_static_mux_check ( .error(1'b1) );
		end
		if (ch_xcvrif_tx_ch_clk_static_mux != "SEL_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_tx_ch_clk_static_mux_check ( .error(1'b1) );
		end
		if (ch_flux_l_tx_bond_size_atom != "TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_bond_size_atom != "TX_BOND_SIZE_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_bond_size_atom != "TX_BOND_SIZE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_bond_size_atom != "RX_BOND_SIZE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_bond_size_atom_check ( .error(1'b1) );
		end
		if (ch_clkrx_refclk_cssm_fw_control_atom != "CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_clkrx_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch_clkrx_refclk_sector_specifies_refclk_ready_atom != "CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_clkrx_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch_local_refclk_cssm_fw_control_atom != "LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_local_refclk_cssm_fw_control_atom_check ( .error(1'b1) );
		end
		if (ch_local_refclk_sector_specifies_refclk_ready_atom != "LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_local_refclk_sector_specifies_refclk_ready_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_postdiv_sel_atom != "TX_PLL_POSTDIV_SEL_SYNTH2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_postdiv_sel_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_bw_sel_atom != "TX_PLL_BW_SEL_LOW")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_bw_sel_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_f_out_hz_atom != 36'b000111011100110101100101000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_f_out_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_f_vco_hz_atom != 36'b001001010100000010111110010000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_f_vco_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_f_pfd_hz_atom != 36'b000000000101111101011110000100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_f_pfd_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_f_ref_hz_atom != 36'b000000000101111101011110000100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_f_ref_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_k_counter_atom != 22'b0000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_k_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_m_counter_atom != 9'b001100100)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_m_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_n_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_n_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_fb_counter_atom != 2'b01)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_fb_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_postdiv_cdr_refclk_hz_atom != 36'b000000000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_postdiv_cdr_refclk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_postdiv_cdr_refclk_divider_atom != 8'b00001100)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_postdiv_cdr_refclk_divider_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_synthdiv_out_divider_atom != 8'b00001100)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_synthdiv_out_divider_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_synthdiv_out_hz_atom != 36'b000000000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_synthdiv_out_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_cdr_f_out_hz_atom != 36'b000111011100110101100101000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_cdr_f_out_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_cdr_f_vco_hz_atom != 36'b001001010100000010111110010000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_cdr_f_vco_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_cdr_f_pfd_hz_atom != 36'b000000000101111101011110000100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_cdr_f_pfd_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_cdr_f_ref_hz_atom != 36'b000000000101111101011110000100000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_cdr_f_ref_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_cdr_l_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_cdr_l_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_cdr_m_counter_atom != 9'b000110010)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_cdr_m_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_cdr_n_counter_atom != 6'b000001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_cdr_n_counter_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_preloaded_hardware_configs_atom != "TX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_protocol_hint_atom != "TX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_datarate_bps_atom != 37'b0001110111001101011001010000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_datarate_bps_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_prbs_gen_en_atom != "TX_PRBS_GEN_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_prbs_gen_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_prbs_pattern_atom != 4'b1001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_user_clk_only_mode_atom != "TX_USER_CLK_ONLY_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_user_clk_only_mode_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_width_atom != "TX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_width_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_word_clk_hz_atom != 36'b000000111011100110101100101000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_word_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_dl_enable_atom != "TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_preloaded_hardware_configs_atom != "RX_PRELOADED_HARDWARE_CONFIGS_PCIE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_preloaded_hardware_configs_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_protocol_hint_atom != "RX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_datarate_bps_atom != 37'b0001110111001101011001010000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_datarate_bps_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_prbs_monitor_en_atom != "RX_PRBS_MONITOR_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_prbs_monitor_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_prbs_pattern_atom != 4'b0000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_prbs_pattern_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_width_atom != "RX_WIDTH_X16")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_width_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_force_cdr_ltr_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_force_cdr_ltr_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_adaptation_mode_atom != "RX_ADAPTATION_MODE_UX_NATIVE_ADAPTATION")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_adaptation_mode_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_word_clk_hz_atom != 36'b000000111011100110101100101000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_word_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_dl_enable_atom != "RX_DL_ENABLE_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch_l_rx_postdiv_clk_en_atom != "RX_POSTDIV_CLK_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_rx_postdiv_clk_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_rx_postdiv_clk_divider_atom != 8'b00001100)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_rx_postdiv_clk_divider_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_postdiv_clk_divider_atom != 8'b10001001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_postdiv_clk_divider_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_refclk_select_atom != "TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch_l_loopback_mode_atom != "LOOPBACK_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_loopback_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_flux_mode_atom != "FLUX_MODE_FLUX_MODE_BYPASS")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_flux_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_rx_protocol_hint_atom != "RX_PROTOCOL_HINT_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_rx_protocol_hint_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_tx_dl_enable_atom != "TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_rx_dl_enable_atom != "RX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_dl_enable_atom != "TX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_dl_enable_atom != "RX_DL_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_dl_enable_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_fifo_mode_atom != "TX_FIFO_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_fifo_mode_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_fifo_mode_atom != "RX_FIFO_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_fifo_mode_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_en_atom != "TRUE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_duplex_mode_atom != "DUPLEX_MODE_DUPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_en_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_en_atom != "FALSE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_en_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_duplex_mode_atom != "DUPLEX_MODE_RX_ONLY_SIMPLEX")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_duplex_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_rx_fec_type_used_atom != "RX_FEC_TYPE_USED_NONE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_rx_fec_type_used_atom_check ( .error(1'b1) );
		end
		if (ch_l_sim_mode_atom != "SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_rx_sim_mode_atom != "RX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_rx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_tx_sim_mode_atom != "TX_SIM_MODE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_tx_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_dr_enabled_atom != "DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_sup_mode_atom != "SUP_MODE_USER_MODE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_sup_mode_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_sim_mode_atom != "SIM_MODE_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_sim_mode_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_dr_enabled_atom != "DR_ENABLED_DR_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_dr_enabled_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_spread_spectrum_en_atom != "TX_SPREAD_SPECTRUM_EN_ENABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_spread_spectrum_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_rx_postdiv_clk_hz_atom != 36'b000000000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_rx_postdiv_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_rx_postdiv_clk_fractional_en_atom != "RX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_rx_postdiv_clk_fractional_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_cdr_refclk_select_atom != "CDR_REFCLK_SELECT_GLOBAL_REFCLK0")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_cdr_refclk_select_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_postdiv_clk_hz_atom != 36'b000000000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_postdiv_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_postdiv_clk_fractional_en_atom != "TX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_postdiv_clk_fractional_en_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_lc_postdiv_sel_atom != "LC_POSTDIV_SEL_SYNTH2")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_lc_postdiv_sel_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom != "TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom != "TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom != "RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom != "RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_gb_width_atom != "TX_GB_WIDTH_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_gb_width_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_gb_width_atom != "RX_GB_WIDTH_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_gb_width_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_dynamic_mux_atom != "TX_DYNAMIC_MUX_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_word_clk_dynamic_mux_atom != "TX_WORD_CLK_DYNAMIC_MUX_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_word_clk_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_word_clk_dynamic_mux_atom != "RX_WORD_CLK_DYNAMIC_MUX_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_word_clk_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom != "TX_FIFO_RD_EN_DYNAMIC_MUX_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom != "RX_FIFO_RD_EN_DYNAMIC_MUX_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_rst_dynamic_mux_atom != "TX_RST_DYNAMIC_MUX_X4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_rst_dynamic_mux_atom_check ( .error(1'b1) );
		end
		if (ch_l_clk_debug_select_0_enable_atom != "CLK_DEBUG_SELECT_0_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_clk_debug_select_0_enable_atom_check ( .error(1'b1) );
		end
		if (ch_l_clk_debug_select_0_setting_atom != "CLK_DEBUG_SELECT_0_SETTING_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_clk_debug_select_0_setting_atom_check ( .error(1'b1) );
		end
		if (ch_l_clk_debug_select_1_enable_atom != "CLK_DEBUG_SELECT_1_ENABLE_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_clk_debug_select_1_enable_atom_check ( .error(1'b1) );
		end
		if (ch_l_clk_debug_select_1_setting_atom != "CLK_DEBUG_SELECT_1_SETTING_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_clk_debug_select_1_setting_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_eq_main_tap_atom != 6'b000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_eq_main_tap_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_eq_post_tap_1_atom != 5'b00000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_eq_post_tap_1_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_eq_pre_tap_1_atom != 5'b00000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_eq_pre_tap_1_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_eq_pre_tap_2_atom != 3'b000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_eq_pre_tap_2_atom_check ( .error(1'b1) );
		end
		if (ch_l_tx_pll_feed_forward_gain_atom != 8'b01000011)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_tx_pll_feed_forward_gain_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_termination_mode_atom != "RX_TERMINATION_MODE_GROUNDED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_termination_mode_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_onchip_termination_setting_atom != "RX_ONCHIP_TERMINATION_SETTING_R_1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_onchip_termination_setting_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_eq_vga_gain_atom != 7'b0100000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_eq_vga_gain_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_x_eq_hf_boost_atom != 6'b100000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_x_eq_hf_boost_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_eq_dfe_tap_1_atom != 6'b000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_eq_dfe_tap_1_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_external_couple_type_atom != "RX_EXTERNAL_COUPLE_TYPE_AC")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_external_couple_type_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_bonding_category_atom != "TX_BONDING_CATEGORY_BONDING_FOLLOWER")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_bonding_category_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_tx_master_pll_mode_atom != "TX_MASTER_PLL_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_tx_master_pll_mode_atom_check ( .error(1'b1) );
		end
		if (ch_l_xcvr_rx_cdrdivout_en_atom != "RX_CDRDIVOUT_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_xcvr_rx_cdrdivout_en_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_tx_bonding_mode_atom != "TX_BONDING_MODE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_tx_bonding_mode_atom_check ( .error(1'b1) );
		end
		if (ch_xcvrif_l_rx_bonding_mode_atom != "RX_BONDING_MODE_UNUSED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_xcvrif_l_rx_bonding_mode_atom_check ( .error(1'b1) );
		end
		if (ch_flux_l_sequencer_reg_en_atom != "SEQUENCER_REG_EN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_flux_l_sequencer_reg_en_atom_check ( .error(1'b1) );
		end
		if (ch_l_speed_grade_atom != "SPEED_GRADE_DASH_1")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_speed_grade_atom_check ( .error(1'b1) );
		end
		if (ch_usb_mode_atom != "USB_MODE_DISABLED")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_usb_mode_atom_check ( .error(1'b1) );
		end
		if (ch_pcie_mode_atom != "PCIE_MODE_GEN4")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_pcie_mode_atom_check ( .error(1'b1) );
		end
		if (ch_l_ick_tx_word_clk_hz_atom != 36'b100101011100000111110010100001110010)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_ick_tx_word_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_pcs_ref_clk_hz_atom != 36'b101001111010110110010111101111110101)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_pcs_ref_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_l_lane_common_ref_clk_hz_atom != 36'b111110010011110101111111101000101001)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_l_lane_common_ref_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_rx_invert_pin_atom != "RX_INVERT_PIN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_rx_invert_pin_atom_check ( .error(1'b1) );
		end
		if (ch_tx_invert_pin_atom != "TX_INVERT_PIN_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_tx_invert_pin_atom_check ( .error(1'b1) );
		end
		if (ch_rx_dl_rx_lat_bit_for_async_atom != 18'b111110100110100101)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_rx_dl_rx_lat_bit_for_async_atom_check ( .error(1'b1) );
		end
		if (ch_rx_dl_rxbit_cntr_pma_atom != "RX_DL_RXBIT_CNTR_PMA_DISABLE")
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_rx_dl_rxbit_cntr_pma_atom_check ( .error(1'b1) );
		end
		if (ch_rx_dl_rxbit_rollover_atom != 18'b001001111001000101)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_rx_dl_rxbit_rollover_atom_check ( .error(1'b1) );
		end
		if (ch_eth_rx_clk_hz_atom != 36'b000000000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_eth_rx_clk_hz_atom_check ( .error(1'b1) );
		end
		if (ch_eth_tx_clk_hz_atom != 36'b000000000000000000000000000000000000)
		begin
		// synthesis translate_off
			initial begin
				$display("Generated module instantiated with wrong parameters");
				$stop;
			end
		// synthesis translate_on
			instantiated_with_wrong_parameters_error_see_comment_above
					ch_eth_tx_clk_hz_atom_check ( .error(1'b1) );
		end
	endgenerate

	system_intel_pcie_gts_0_phy_hal_2100_xvyrmby #(
		.ch_xcvrif_l_loopback_mode_atom                     ("LOOPBACK_MODE_DISABLE"),
		.ch_flux_l_stmux_rx_demux_sel                       ("SEL_PCIE_PCS"),
		.ch_flux_l_stmux_rx_rxword_clk_demux_sel            ("SEL_PCIE_RXWORD_CLK"),
		.ch_flux_l_stmux_tx_txword_clk_demux_sel            ("SEL_PCIE_TXWORD_CLK"),
		.ch_flux_l_stmux_tx_mux_sel                         ("SEL_PCIE_PCS"),
		.ch_flux_l_stmux_tx_txword_clk_mux_sel              ("SEL_UX_OCK_PMA_CLK"),
		.ch_xcvrif_rx_ch_clk_static_mux                     ("SEL_UNUSED"),
		.ch_xcvrif_tx_ch_clk_static_mux                     ("SEL_UNUSED"),
		.ch_flux_l_tx_bond_size_atom                        ("TX_BOND_SIZE_X4"),
		.ch_l_xcvr_tx_bond_size_atom                        ("TX_BOND_SIZE_X4"),
		.ch_xcvrif_l_tx_bond_size_atom                      ("TX_BOND_SIZE_UNUSED"),
		.ch_xcvrif_l_rx_bond_size_atom                      ("RX_BOND_SIZE_UNUSED"),
		.ch_clkrx_refclk_cssm_fw_control_atom               ("CLKRX_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch_clkrx_refclk_sector_specifies_refclk_ready_atom ("CLKRX_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch_local_refclk_cssm_fw_control_atom               ("LOCAL_REFCLK_CSSM_FW_CONTROL_DISABLE"),
		.ch_local_refclk_sector_specifies_refclk_ready_atom ("LOCAL_REFCLK_SECTOR_SPECIFIES_REFCLK_READY_DISABLE"),
		.ch_l_tx_pll_postdiv_sel_atom                       ("TX_PLL_POSTDIV_SEL_SYNTH2"),
		.ch_l_tx_pll_bw_sel_atom                            ("TX_PLL_BW_SEL_LOW"),
		.ch_l_tx_pll_f_out_hz_atom                          (36'b000111011100110101100101000000000000),
		.ch_l_tx_pll_f_vco_hz_atom                          (36'b001001010100000010111110010000000000),
		.ch_l_tx_pll_f_pfd_hz_atom                          (36'b000000000101111101011110000100000000),
		.ch_l_tx_pll_f_ref_hz_atom                          (36'b000000000101111101011110000100000000),
		.ch_l_tx_pll_k_counter_atom                         (22'b0000000000000000000000),
		.ch_l_tx_pll_l_counter_atom                         (6'b000001),
		.ch_l_tx_pll_m_counter_atom                         (9'b001100100),
		.ch_l_tx_pll_n_counter_atom                         (6'b000001),
		.ch_l_tx_pll_fb_counter_atom                        (2'b01),
		.ch_l_tx_postdiv_cdr_refclk_hz_atom                 (36'b000000000000000000000000000000000000),
		.ch_l_tx_postdiv_cdr_refclk_divider_atom            (8'b00001100),
		.ch_l_tx_synthdiv_out_divider_atom                  (8'b00001100),
		.ch_l_tx_synthdiv_out_hz_atom                       (36'b000000000000000000000000000000000000),
		.ch_l_xcvr_cdr_f_out_hz_atom                        (36'b000111011100110101100101000000000000),
		.ch_l_xcvr_cdr_f_vco_hz_atom                        (36'b001001010100000010111110010000000000),
		.ch_l_xcvr_cdr_f_pfd_hz_atom                        (36'b000000000101111101011110000100000000),
		.ch_l_xcvr_cdr_f_ref_hz_atom                        (36'b000000000101111101011110000100000000),
		.ch_l_cdr_l_counter_atom                            (6'b000001),
		.ch_l_cdr_m_counter_atom                            (9'b000110010),
		.ch_l_cdr_n_counter_atom                            (6'b000001),
		.ch_l_xcvr_tx_preloaded_hardware_configs_atom       ("TX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch_l_xcvr_tx_protocol_hint_atom                    ("TX_PROTOCOL_HINT_DISABLED"),
		.ch_l_xcvr_tx_datarate_bps_atom                     (37'b0001110111001101011001010000000000000),
		.ch_l_xcvr_tx_prbs_gen_en_atom                      ("TX_PRBS_GEN_EN_DISABLE"),
		.ch_l_xcvr_tx_prbs_pattern_atom                     (4'b1001),
		.ch_l_xcvr_tx_user_clk_only_mode_atom               ("TX_USER_CLK_ONLY_MODE_DISABLE"),
		.ch_l_xcvr_tx_width_atom                            ("TX_WIDTH_X16"),
		.ch_l_xcvr_tx_word_clk_hz_atom                      (36'b000000111011100110101100101000000000),
		.ch_l_xcvr_tx_dl_enable_atom                        ("TX_DL_ENABLE_DISABLE"),
		.ch_l_xcvr_rx_preloaded_hardware_configs_atom       ("RX_PRELOADED_HARDWARE_CONFIGS_PCIE"),
		.ch_l_xcvr_rx_protocol_hint_atom                    ("RX_PROTOCOL_HINT_DISABLED"),
		.ch_l_xcvr_rx_datarate_bps_atom                     (37'b0001110111001101011001010000000000000),
		.ch_l_xcvr_rx_prbs_monitor_en_atom                  ("RX_PRBS_MONITOR_EN_DISABLE"),
		.ch_l_xcvr_rx_prbs_pattern_atom                     (4'b0000),
		.ch_l_xcvr_rx_width_atom                            ("RX_WIDTH_X16"),
		.ch_l_xcvr_rx_force_cdr_ltr_atom                    ("TRUE"),
		.ch_l_xcvr_rx_adaptation_mode_atom                  ("RX_ADAPTATION_MODE_UX_NATIVE_ADAPTATION"),
		.ch_l_xcvr_rx_word_clk_hz_atom                      (36'b000000111011100110101100101000000000),
		.ch_l_xcvr_rx_dl_enable_atom                        ("RX_DL_ENABLE_ENABLE"),
		.ch_l_rx_postdiv_clk_en_atom                        ("RX_POSTDIV_CLK_EN_ENABLE"),
		.ch_l_rx_postdiv_clk_divider_atom                   (8'b00001100),
		.ch_l_tx_postdiv_clk_divider_atom                   (8'b10001001),
		.ch_l_tx_pll_refclk_select_atom                     ("TX_PLL_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch_l_loopback_mode_atom                            ("LOOPBACK_MODE_DISABLED"),
		.ch_flux_l_flux_mode_atom                           ("FLUX_MODE_FLUX_MODE_BYPASS"),
		.ch_flux_l_rx_protocol_hint_atom                    ("RX_PROTOCOL_HINT_DISABLED"),
		.ch_flux_l_tx_dl_enable_atom                        ("TX_DL_ENABLE_DISABLE"),
		.ch_flux_l_rx_dl_enable_atom                        ("RX_DL_ENABLE_DISABLE"),
		.ch_xcvrif_l_tx_dl_enable_atom                      ("TX_DL_ENABLE_DISABLE"),
		.ch_xcvrif_l_rx_dl_enable_atom                      ("RX_DL_ENABLE_DISABLE"),
		.ch_xcvrif_l_tx_fifo_mode_atom                      ("TX_FIFO_MODE_DISABLED"),
		.ch_xcvrif_l_rx_fifo_mode_atom                      ("RX_FIFO_MODE_DISABLED"),
		.ch_l_xcvr_tx_en_atom                               ("TRUE"),
		.ch_l_xcvr_rx_en_atom                               ("TRUE"),
		.ch_l_duplex_mode_atom                              ("DUPLEX_MODE_DUPLEX"),
		.ch_xcvrif_l_tx_en_atom                             ("FALSE"),
		.ch_xcvrif_l_rx_en_atom                             ("FALSE"),
		.ch_xcvrif_l_duplex_mode_atom                       ("DUPLEX_MODE_RX_ONLY_SIMPLEX"),
		.ch_flux_l_rx_fec_type_used_atom                    ("RX_FEC_TYPE_USED_NONE"),
		.ch_l_sim_mode_atom                                 ("SIM_MODE_DISABLE"),
		.ch_flux_l_rx_sim_mode_atom                         ("RX_SIM_MODE_DISABLE"),
		.ch_flux_l_tx_sim_mode_atom                         ("TX_SIM_MODE_DISABLE"),
		.ch_flux_l_dr_enabled_atom                          ("DR_ENABLED_DR_DISABLED"),
		.ch_xcvrif_l_sup_mode_atom                          ("SUP_MODE_USER_MODE"),
		.ch_xcvrif_l_sim_mode_atom                          ("SIM_MODE_ENABLE"),
		.ch_xcvrif_l_dr_enabled_atom                        ("DR_ENABLED_DR_DISABLED"),
		.ch_l_xcvr_tx_spread_spectrum_en_atom               ("TX_SPREAD_SPECTRUM_EN_ENABLE"),
		.ch_l_rx_postdiv_clk_hz_atom                        (36'b000000000000000000000000000000000000),
		.ch_l_rx_postdiv_clk_fractional_en_atom             ("RX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE"),
		.ch_l_cdr_refclk_select_atom                        ("CDR_REFCLK_SELECT_GLOBAL_REFCLK0"),
		.ch_l_tx_postdiv_clk_hz_atom                        (36'b000000000000000000000000000000000000),
		.ch_l_tx_postdiv_clk_fractional_en_atom             ("TX_POSTDIV_CLK_FRACTIONAL_EN_DISABLE"),
		.ch_flux_l_lc_postdiv_sel_atom                      ("LC_POSTDIV_SEL_SYNTH2"),
		.ch_flux_l_tx_user1_clk_mux_dynamic_sel_atom        ("TX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch_flux_l_tx_user2_clk_mux_dynamic_sel_atom        ("TX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_TXWORD_CLK"),
		.ch_flux_l_rx_user1_clk_mux_dynamic_sel_atom        ("RX_USER1_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch_flux_l_rx_user2_clk_mux_dynamic_sel_atom        ("RX_USER2_CLK_MUX_DYNAMIC_SEL_OCK_PCS_RXWORD"),
		.ch_xcvrif_l_tx_gb_width_atom                       ("TX_GB_WIDTH_DISABLED"),
		.ch_xcvrif_l_rx_gb_width_atom                       ("RX_GB_WIDTH_DISABLED"),
		.ch_xcvrif_l_tx_dynamic_mux_atom                    ("TX_DYNAMIC_MUX_UNUSED"),
		.ch_xcvrif_l_tx_word_clk_dynamic_mux_atom           ("TX_WORD_CLK_DYNAMIC_MUX_X4"),
		.ch_xcvrif_l_rx_word_clk_dynamic_mux_atom           ("RX_WORD_CLK_DYNAMIC_MUX_UNUSED"),
		.ch_xcvrif_l_tx_fifo_rd_en_dynamic_mux_atom         ("TX_FIFO_RD_EN_DYNAMIC_MUX_X4"),
		.ch_xcvrif_l_rx_fifo_rd_en_dynamic_mux_atom         ("RX_FIFO_RD_EN_DYNAMIC_MUX_UNUSED"),
		.ch_xcvrif_l_tx_rst_dynamic_mux_atom                ("TX_RST_DYNAMIC_MUX_X4"),
		.ch_l_clk_debug_select_0_enable_atom                ("CLK_DEBUG_SELECT_0_ENABLE_DISABLE"),
		.ch_l_clk_debug_select_0_setting_atom               ("CLK_DEBUG_SELECT_0_SETTING_DISABLED"),
		.ch_l_clk_debug_select_1_enable_atom                ("CLK_DEBUG_SELECT_1_ENABLE_DISABLE"),
		.ch_l_clk_debug_select_1_setting_atom               ("CLK_DEBUG_SELECT_1_SETTING_DISABLED"),
		.ch_l_xcvr_tx_eq_main_tap_atom                      (6'b000000),
		.ch_l_xcvr_tx_eq_post_tap_1_atom                    (5'b00000),
		.ch_l_xcvr_tx_eq_pre_tap_1_atom                     (5'b00000),
		.ch_l_xcvr_tx_eq_pre_tap_2_atom                     (3'b000),
		.ch_l_tx_pll_feed_forward_gain_atom                 (8'b01000011),
		.ch_l_xcvr_rx_termination_mode_atom                 ("RX_TERMINATION_MODE_GROUNDED"),
		.ch_l_xcvr_rx_onchip_termination_setting_atom       ("RX_ONCHIP_TERMINATION_SETTING_R_1"),
		.ch_l_xcvr_rx_eq_vga_gain_atom                      (7'b0100000),
		.ch_l_xcvr_x_eq_hf_boost_atom                       (6'b100000),
		.ch_l_xcvr_rx_eq_dfe_tap_1_atom                     (6'b000000),
		.ch_l_xcvr_rx_external_couple_type_atom             ("RX_EXTERNAL_COUPLE_TYPE_AC"),
		.ch_l_xcvr_tx_bonding_category_atom                 ("TX_BONDING_CATEGORY_BONDING_FOLLOWER"),
		.ch_l_xcvr_tx_master_pll_mode_atom                  ("TX_MASTER_PLL_MODE_DISABLED"),
		.ch_l_xcvr_rx_cdrdivout_en_atom                     ("RX_CDRDIVOUT_EN_DISABLE"),
		.ch_xcvrif_l_tx_bonding_mode_atom                   ("TX_BONDING_MODE_UNUSED"),
		.ch_xcvrif_l_rx_bonding_mode_atom                   ("RX_BONDING_MODE_UNUSED"),
		.ch_flux_l_sequencer_reg_en_atom                    ("SEQUENCER_REG_EN_DISABLE"),
		.ch_l_speed_grade_atom                              ("SPEED_GRADE_DASH_1"),
		.ch_usb_mode_atom                                   ("USB_MODE_DISABLED"),
		.ch_pcie_mode_atom                                  ("PCIE_MODE_GEN4"),
		.ch_l_ick_tx_word_clk_hz_atom                       (36'b100101011100000111110010100001110010),
		.ch_l_pcs_ref_clk_hz_atom                           (36'b101001111010110110010111101111110101),
		.ch_l_lane_common_ref_clk_hz_atom                   (36'b111110010011110101111111101000101001),
		.ch_rx_invert_pin_atom                              ("RX_INVERT_PIN_DISABLE"),
		.ch_tx_invert_pin_atom                              ("TX_INVERT_PIN_DISABLE"),
		.ch_rx_dl_rx_lat_bit_for_async_atom                 (18'b111110100110100101),
		.ch_rx_dl_rxbit_cntr_pma_atom                       ("RX_DL_RXBIT_CNTR_PMA_DISABLE"),
		.ch_rx_dl_rxbit_rollover_atom                       (18'b001001111001000101),
		.ch_eth_rx_clk_hz_atom                              (36'b000000000000000000000000000000000000),
		.ch_eth_tx_clk_hz_atom                              (36'b000000000000000000000000000000000000)
	) phy_hal_top (
		.oflux_xoa_tx_n_l0_ux              (oflux_xoa_tx_n_l0_ux),              //  output,    width = 1,              oflux_xoa_tx_n_l0_ux.data
		.oflux_xoa_tx_p_l0_ux              (oflux_xoa_tx_p_l0_ux),              //  output,    width = 1,              oflux_xoa_tx_p_l0_ux.data
		.iflux_xia_rx_n_l0_ux              (iflux_xia_rx_n_l0_ux),              //   input,    width = 1,              iflux_xia_rx_n_l0_ux.data
		.iflux_xia_rx_p_l0_ux              (iflux_xia_rx_p_l0_ux),              //   input,    width = 1,              iflux_xia_rx_p_l0_ux.data
		.i_ss_async_pldif                  (i_ss_async_pldif),                  //   input,   width = 80,                       asyncdata_0.data
		.o_ss_async_pldif                  (o_ss_async_pldif),                  //  output,   width = 50,                       asyncdata_1.data
		.i_ss_async_pldif_pcie_mux         (i_ss_async_pldif_pcie_mux),         //   input,   width = 80,                       asyncdata_2.data
		.i_lavmm_addr                      (i_lavmm_addr),                      //   input,   width = 20,                          reconfig.address
		.i_lavmm_be                        (i_lavmm_be),                        //   input,    width = 4,                                  .byteenable
		.i_lavmm_read                      (i_lavmm_read),                      //   input,    width = 1,                                  .read
		.i_lavmm_wdata                     (i_lavmm_wdata),                     //   input,   width = 32,                                  .writedata
		.i_lavmm_write                     (i_lavmm_write),                     //   input,    width = 1,                                  .write
		.o_lavmm_rdata                     (o_lavmm_rdata),                     //  output,   width = 32,                                  .readdata
		.o_lavmm_rdata_valid               (o_lavmm_rdata_valid),               //  output,    width = 1,                                  .readdatavalid
		.o_lavmm_waitreq                   (o_lavmm_waitreq),                   //  output,    width = 1,                                  .waitrequest
		.i_lavmm_clk                       (i_lavmm_clk),                       //   input,    width = 1,                      reconfig_clk.clk
		.i_lavmm_rstn                      (i_lavmm_rstn),                      //   input,    width = 1,                      reconfig_rst.reset
		.i_ft_rx_sclk_sync_ch              (i_ft_rx_sclk_sync_ch),              //   input,    width = 1,              i_ft_rx_sclk_sync_ch.clk
		.i_ft_tx_sclk_sync_ch              (i_ft_tx_sclk_sync_ch),              //   input,    width = 1,              i_ft_tx_sclk_sync_ch.clk
		.o_ft_rx_async_pulse_ch            (o_ft_rx_async_pulse_ch),            //  output,    width = 1,            o_ft_rx_async_pulse_ch.clk
		.o_ft_tx_async_pulse_ch            (o_ft_tx_async_pulse_ch),            //  output,    width = 1,            o_ft_tx_async_pulse_ch.clk
		.o_rxcdrlock2dataa                 (o_rxcdrlock2dataa),                 //  output,    width = 1,                 o_rxcdrlock2dataa.lockdata
		.i_rst_ux_rx_sfrz                  (i_rst_ux_rx_sfrz),                  //   input,    width = 1,                  i_rst_ux_rx_sfrz.data
		.o_rst_flux0_cpi_cmn_busy          (o_rst_flux0_cpi_cmn_busy),          //  output,    width = 1,          o_rst_flux0_cpi_cmn_busy.busy
		.o_rst_oflux_rx_srds_rdy           (o_rst_oflux_rx_srds_rdy),           //  output,    width = 1,           o_rst_oflux_rx_srds_rdy.ready
		.o_rst_ux_all_synthlockstatus      (o_rst_ux_all_synthlockstatus),      //  output,    width = 1,      o_rst_ux_all_synthlockstatus.status
		.o_rst_ux_rxcdrlockstatus          (o_rst_ux_rxcdrlockstatus),          //  output,    width = 1,          o_rst_ux_rxcdrlockstatus.rxstatus
		.o_ux_tx_ch_ptr_smpl               (o_ux_tx_ch_ptr_smpl),               //  output,    width = 1,               o_ux_tx_ch_ptr_smpl.sample
		.i_ick_sclk_tx                     (i_ick_sclk_tx),                     //   input,    width = 1,                     i_ick_sclk_tx.clk
		.i_ick_sclk_rx                     (i_ick_sclk_rx),                     //   input,    width = 1,                     i_ick_sclk_rx.clk
		.i_rst_pld_ux_tx_pma_rst_n         (i_rst_pld_ux_tx_pma_rst_n),         //   input,    width = 1,         i_rst_pld_ux_tx_pma_rst_n.reset
		.i_rst_pld_ux_rx_pma_rst_n         (i_rst_pld_ux_rx_pma_rst_n),         //   input,    width = 1,         i_rst_pld_ux_rx_pma_rst_n.reset
		.o_ch_lavmm_xcvrif_rdata           (o_ch_lavmm_xcvrif_rdata),           //  output,   width = 32,                     reconfig_xcvr.readdata
		.o_ch_lavmm_xcvrif_rdata_valid     (o_ch_lavmm_xcvrif_rdata_valid),     //  output,    width = 1,                                  .readdatavalid
		.o_ch_lavmm_xcvrif_waitreq         (o_ch_lavmm_xcvrif_waitreq),         //  output,    width = 1,                                  .waitrequest
		.i_ch_lavmm_xcvrif_addr            (i_ch_lavmm_xcvrif_addr),            //   input,   width = 20,                                  .address
		.i_ch_lavmm_xcvrif_be              (i_ch_lavmm_xcvrif_be),              //   input,    width = 4,                                  .byteenable
		.i_ch_lavmm_xcvrif_read            (i_ch_lavmm_xcvrif_read),            //   input,    width = 1,                                  .read
		.i_ch_lavmm_xcvrif_wdata           (i_ch_lavmm_xcvrif_wdata),           //   input,   width = 32,                                  .writedata
		.i_ch_lavmm_xcvrif_write           (i_ch_lavmm_xcvrif_write),           //   input,    width = 1,                                  .write
		.i_ch_lavmm_xcvrif_clk             (i_ch_lavmm_xcvrif_clk),             //   input,    width = 1,                 reconfig_clk_xcvr.clk
		.i_ch_lavmm_xcvrif_rstn            (i_ch_lavmm_xcvrif_rstn),            //   input,    width = 1,                 reconfig_rst_xcvr.reset
		.o_rx_latency_pulse                (o_rx_latency_pulse),                //  output,    width = 1,                o_rx_latency_pulse.clk
		.o_tx_latency_pulse                (o_tx_latency_pulse),                //  output,    width = 1,                o_tx_latency_pulse.clk
		.i_ch_eth_xcvrif_tx_async          (i_ch_eth_xcvrif_tx_async),          //   input,    width = 7,                       asyncdata_3.data
		.i_ch_eth_xcvrif_tx_direct         (i_ch_eth_xcvrif_tx_direct),         //   input,    width = 1,                       asyncdata_4.data
		.o_ch_eth_xcvrif_rx_async          (o_ch_eth_xcvrif_rx_async),          //  output,   width = 14,                       asyncdata_5.data
		.o_ch_eth_xcvrif_rx_direct         (o_ch_eth_xcvrif_rx_direct),         //  output,    width = 1,                       asyncdata_6.data
		.i_rstxcvrif_xcvrif_signal_ok      (i_rstxcvrif_xcvrif_signal_ok),      //   input,    width = 1,      i_rstxcvrif_xcvrif_signal_ok.data
		.i_rstxcvrif_rx_xcvrif_sfrz_n      (i_rstxcvrif_rx_xcvrif_sfrz_n),      //   input,    width = 1,      i_rstxcvrif_rx_xcvrif_sfrz_n.data
		.i_rstxcvrif_xcvrif_rx_rst_n       (i_rstxcvrif_xcvrif_rx_rst_n),       //   input,    width = 1,       i_rstxcvrif_xcvrif_rx_rst_n.data
		.i_rstxcvrif_tx_xcvrif_sfrz_n      (i_rstxcvrif_tx_xcvrif_sfrz_n),      //   input,    width = 1,      i_rstxcvrif_tx_xcvrif_sfrz_n.data
		.i_rstxcvrif_xcvrif_tx_rst_n       (i_rstxcvrif_xcvrif_tx_rst_n),       //   input,    width = 1,       i_rstxcvrif_xcvrif_tx_rst_n.data
		.o_pma_rx_sf                       (o_pma_rx_sf),                       //  output,    width = 1,                       o_pma_rx_sf.data
		.i_xcvrif_tx_mux_data              (i_xcvrif_tx_mux_data),              //   input,   width = 43,              i_xcvrif_tx_mux_data.data
		.o_rx_data                         (o_rx_data),                         //  output,   width = 43,                         o_rx_data.data
		.o_tx_source_sel                   (o_tx_source_sel),                   //  output,    width = 2,                   o_tx_source_sel.data
		.o_rx_fifo_en_sel                  (o_rx_fifo_en_sel),                  //  output,    width = 3,                  o_rx_fifo_en_sel.data
		.o_tx_rst_source_sel               (o_tx_rst_source_sel),               //  output,    width = 3,               o_tx_rst_source_sel.data
		.i_ch_xcvrif_rx_fifo_rd_en         (i_ch_xcvrif_rx_fifo_rd_en),         //   input,    width = 1,         i_ch_xcvrif_rx_fifo_rd_en.data
		.o_ch_xcvrif_rx_fifo_rd_en         (o_ch_xcvrif_rx_fifo_rd_en),         //  output,    width = 1,         o_ch_xcvrif_rx_fifo_rd_en.data
		.i_ch_xcvrif_tx_fifo_rd_en         (i_ch_xcvrif_tx_fifo_rd_en),         //   input,    width = 1,         i_ch_xcvrif_tx_fifo_rd_en.data
		.o_ch_xcvrif_tx_fifo_rd_en         (o_ch_xcvrif_tx_fifo_rd_en),         //  output,    width = 1,         o_ch_xcvrif_tx_fifo_rd_en.data
		.o_ux_rxuser1_sel                  (o_ux_rxuser1_sel),                  //  output,    width = 2,                  o_ux_rxuser1_sel.data
		.o_ux_rxuser2_sel                  (o_ux_rxuser2_sel),                  //  output,    width = 2,                  o_ux_rxuser2_sel.data
		.o_ux_txuser1_sel                  (o_ux_txuser1_sel),                  //  output,    width = 2,                  o_ux_txuser1_sel.data
		.o_ux_txuser2_sel                  (o_ux_txuser2_sel),                  //  output,    width = 2,                  o_ux_txuser2_sel.data
		.o_pcs_rxpostdiv                   (o_pcs_rxpostdiv),                   //  output,    width = 1,                   o_pcs_rxpostdiv.data
		.o_pcs_rxword                      (o_pcs_rxword),                      //  output,    width = 1,                      o_pcs_rxword.data
		.o_ux_txlc_clk                     (o_ux_txlc_clk),                     //  output,    width = 1,                     o_ux_txlc_clk.clk
		.o_tx_xcvr_wordclk_sel             (o_tx_xcvr_wordclk_sel),             //  output,    width = 3,             o_tx_xcvr_wordclk_sel.data
		.o_rx_xcvr_wordclk_sel             (o_rx_xcvr_wordclk_sel),             //  output,    width = 2,             o_rx_xcvr_wordclk_sel.data
		.i_eth_rx_ch_clk                   (i_eth_rx_ch_clk),                   //   input,    width = 1,                   i_eth_rx_ch_clk.clk
		.uxwrap_bus_in                     (uxwrap_bus_in),                     //   input,  width = 768,                     uxwrap_bus_in.data
		.uxwrap_bus_out                    (uxwrap_bus_out),                    //  output,  width = 704,                    uxwrap_bus_out.data
		.o_lavmm_addr                      (o_lavmm_addr),                      //  output,   width = 20,               reconfig_phy_shared.address
		.o_lavmm_be                        (o_lavmm_be),                        //  output,    width = 4,                                  .byteenable
		.o_lavmm_read                      (o_lavmm_read),                      //  output,    width = 1,                                  .read
		.o_lavmm_wdata                     (o_lavmm_wdata),                     //  output,   width = 32,                                  .writedata
		.o_lavmm_write                     (o_lavmm_write),                     //  output,    width = 1,                                  .write
		.i_lavmm_rdata                     (i_lavmm_rdata),                     //   input,   width = 32,                                  .readdata
		.i_lavmm_rdata_valid               (i_lavmm_rdata_valid),               //   input,    width = 1,                                  .readdatavalid
		.i_lavmm_waitreq                   (i_lavmm_waitreq),                   //   input,    width = 1,                                  .waitrequest
		.o_lavmm_clk                       (o_lavmm_clk),                       //  output,    width = 1,           reconfig_clk_phy_shared.clk
		.o_lavmm_rstn                      (o_lavmm_rstn),                      //  output,    width = 1,           reconfig_rst_phy_shared.reset
		.o_sclk_return_sel_rx              (o_sclk_return_sel_rx),              //  output,    width = 1,              o_sclk_return_sel_rx.data
		.o_sclk_return_sel_tx              (o_sclk_return_sel_tx),              //  output,    width = 1,              o_sclk_return_sel_tx.data
		.o_ick_sclk_rx                     (o_ick_sclk_rx),                     //  output,    width = 1,                     o_ick_sclk_rx.clk
		.i_sync_common_control             (i_sync_common_control),             //   input,    width = 5,             i_sync_common_control.data
		.o_ft_rx_sclk_sync_ch              (o_ft_rx_sclk_sync_ch),              //  output,    width = 1,              o_ft_rx_sclk_sync_ch.data
		.o_ft_tx_sclk_sync_ch              (o_ft_tx_sclk_sync_ch),              //  output,    width = 1,              o_ft_tx_sclk_sync_ch.data
		.o_rst_ux_rx_pma_rst_n             (o_rst_ux_rx_pma_rst_n),             //  output,    width = 1,             o_rst_ux_rx_pma_rst_n.reset
		.o_rst_ux_tx_pma_rst_n             (o_rst_ux_tx_pma_rst_n),             //  output,    width = 1,             o_rst_ux_tx_pma_rst_n.reset
		.o_ick_pcs_txword                  (o_ick_pcs_txword),                  //  output,    width = 1,                  o_ick_pcs_txword.data
		.o_tx_dl_ch_bit                    (o_tx_dl_ch_bit),                    //  output,    width = 1,                    o_tx_dl_ch_bit.data
		.i_dat_pcs_measlatbit              (i_dat_pcs_measlatbit),              //   input,    width = 1,              i_dat_pcs_measlatbit.data
		.i_ft_rx_async_pulse_ch            (i_ft_rx_async_pulse_ch),            //   input,    width = 1,            i_ft_rx_async_pulse_ch.data
		.i_ft_tx_async_pulse_ch            (i_ft_tx_async_pulse_ch),            //   input,    width = 1,            i_ft_tx_async_pulse_ch.data
		.i_rx_dl_ch_bit                    (i_rx_dl_ch_bit),                    //   input,    width = 1,                    i_rx_dl_ch_bit.data
		.i_ux_rxuser1_sel                  (i_ux_rxuser1_sel),                  //   input,    width = 2,                  i_ux_rxuser1_sel.data
		.i_ux_rxuser2_sel                  (i_ux_rxuser2_sel),                  //   input,    width = 2,                  i_ux_rxuser2_sel.data
		.i_ux_txuser1_sel                  (i_ux_txuser1_sel),                  //   input,    width = 2,                  i_ux_txuser1_sel.data
		.i_ux_txuser2_sel                  (i_ux_txuser2_sel),                  //   input,    width = 2,                  i_ux_txuser2_sel.data
		.o_octl_pcs_txstatus_a             (o_octl_pcs_txstatus_a),             //  output,    width = 1,             o_octl_pcs_txstatus_a.data
		.i_ictl_pcs_txenable_a             (i_ictl_pcs_txenable_a),             //   input,    width = 1,             i_ictl_pcs_txenable_a.data
		.i_sync_cfg_data                   (i_sync_cfg_data),                   //   input,  width = 125,                   i_sync_cfg_data.data
		.i_sync_interface_control          (i_sync_interface_control),          //   input,  width = 250,          i_sync_interface_control.data
		.o_tx_data                         (o_tx_data),                         //  output,   width = 80,                         o_tx_data.data
		.i_rx_data                         (i_rx_data),                         //   input,   width = 80,                         i_rx_data.data
		.o_sm_flux_ingress                 (o_sm_flux_ingress),                 //  output,  width = 320,                 o_sm_flux_ingress.data
		.i_sm_flux_egress                  (i_sm_flux_egress),                  //   input,  width = 257,                  i_sm_flux_egress.data
		.i_flux_cpi_int                    (i_flux_cpi_int),                    //   input,    width = 1,                    i_flux_cpi_int.data
		.i_flux_int                        (i_flux_int),                        //   input,    width = 1,                        i_flux_int.data
		.i_oflux_octl_pcs_txptr_smpl_lane  (i_oflux_octl_pcs_txptr_smpl_lane),  //   input,    width = 1,  i_oflux_octl_pcs_txptr_smpl_lane.data
		.o_ick_sclk_tx                     (o_ick_sclk_tx),                     //  output,    width = 1,                     o_ick_sclk_tx.clk
		.i_flux_srds_rdy                   (i_flux_srds_rdy),                   //   input,    width = 1,                   i_flux_srds_rdy.data
		.i_pcs_rxword                      (i_pcs_rxword),                      //   input,    width = 1,                      i_pcs_rxword.data
		.i_pcs_rxpostdiv                   (i_pcs_rxpostdiv),                   //   input,    width = 1,                   i_pcs_rxpostdiv.data
		.i_ock_pcs_txword                  (i_ock_pcs_txword),                  //   input,    width = 1,                  i_ock_pcs_txword.data
		.o_dat_pcs_measlatrndtripbit       (o_dat_pcs_measlatrndtripbit),       //  output,    width = 1,       o_dat_pcs_measlatrndtripbit.data
		.o_ock_pcs_cdrfbclk                (o_ock_pcs_cdrfbclk),                //  output,    width = 1,                o_ock_pcs_cdrfbclk.data
		.o_ock_pcs_ref                     (o_ock_pcs_ref),                     //  output,    width = 1,                     o_ock_pcs_ref.data
		.o_pcie_pcs                        (o_pcie_pcs),                        //  output,   width = 40,                        o_pcie_pcs.data
		.i_pcie_pcs                        (i_pcie_pcs),                        //   input,   width = 40,                        i_pcie_pcs.data
		.i_sel_rxword_clk                  (i_sel_rxword_clk),                  //   input,    width = 1,                  i_sel_rxword_clk.clk
		.i_xcvr_txword_clk                 (i_xcvr_txword_clk),                 //   input,    width = 1,                 i_xcvr_txword_clk.clk
		.o_pcie_rxword_clk                 (o_pcie_rxword_clk),                 //  output,    width = 1,                 o_pcie_rxword_clk.clk
		.o_eth_rxword_clk                  (o_eth_rxword_clk),                  //  output,    width = 1,                  o_eth_rxword_clk.clk
		.o_pcie_txword_clk                 (o_pcie_txword_clk),                 //  output,    width = 1,                 o_pcie_txword_clk.clk
		.o_eth_txword_clk                  (o_eth_txword_clk),                  //  output,    width = 1,                  o_eth_txword_clk.clk
		.o_ock_pcs_txword                  (o_ock_pcs_txword),                  //  output,    width = 1,                  o_ock_pcs_txword.clk
		.o_eth_rx_ch_clk                   (o_eth_rx_ch_clk),                   //  output,    width = 1,                   o_eth_rx_ch_clk.clk
		.o_eth_tx_ch_clk                   (o_eth_tx_ch_clk),                   //  output,    width = 1,                   o_eth_tx_ch_clk.clk
		.ioack_ref_left_p_ux_bidir_in      (ioack_ref_left_p_ux_bidir_in),      //   input,    width = 6,      ioack_ref_left_p_ux_bidir_in.data
		.ioack_hsref_left_p_ux_bidir_in    (ioack_hsref_left_p_ux_bidir_in),    //   input,    width = 1,    ioack_hsref_left_p_ux_bidir_in.clk
		.ioack_cdrdiv_left_ux_bidir_in     (ioack_cdrdiv_left_ux_bidir_in),     //   input,    width = 1,     ioack_cdrdiv_left_ux_bidir_in.clk
		.ioack_synthdiv1_left_ux_bidir_in  (ioack_synthdiv1_left_ux_bidir_in),  //   input,    width = 1,  ioack_synthdiv1_left_ux_bidir_in.clk
		.ioack_synthdiv2_left_ux_bidir_in  (ioack_synthdiv2_left_ux_bidir_in),  //   input,    width = 1,  ioack_synthdiv2_left_ux_bidir_in.clk
		.ioack_cdrdiv_left_ux_bidir_out    (ioack_cdrdiv_left_ux_bidir_out),    //  output,    width = 1,    ioack_cdrdiv_left_ux_bidir_out.clk
		.ioack_synthdiv1_left_ux_bidir_out (ioack_synthdiv1_left_ux_bidir_out), //  output,    width = 1, ioack_synthdiv1_left_ux_bidir_out.clk
		.ioack_synthdiv2_left_ux_bidir_out (ioack_synthdiv2_left_ux_bidir_out), //  output,    width = 1, ioack_synthdiv2_left_ux_bidir_out.clk
		.o_rxeq_best_eye_vala              (o_rxeq_best_eye_vala),              //  output,   width = 14,              o_rxeq_best_eye_vala.data
		.o_rxeq_donea                      (o_rxeq_donea),                      //  output,    width = 1,                      o_rxeq_donea.data
		.o_rxmargin_nacka                  (o_rxmargin_nacka),                  //  output,    width = 1,                  o_rxmargin_nacka.data
		.o_rxmargin_statusa                (o_rxmargin_statusa),                //  output,    width = 1,                o_rxmargin_statusa.data
		.o_rxsignaldetect_lfpsa            (o_rxsignaldetect_lfpsa),            //  output,    width = 1,            o_rxsignaldetect_lfpsa.data
		.o_rxsignaldetecta                 (o_rxsignaldetecta),                 //  output,    width = 1,                 o_rxsignaldetecta.data
		.o_rxmargin_status_gray            (o_rxmargin_status_gray),            //  output,    width = 2,            o_rxmargin_status_gray.data
		.o_rxstatusa                       (o_rxstatusa),                       //  output,    width = 1,                       o_rxstatusa.data
		.o_synthlcfast_postdiv             (o_synthlcfast_postdiv),             //  output,    width = 1,             o_synthlcfast_postdiv.data
		.o_synthlcmed_postdiv              (o_synthlcmed_postdiv),              //  output,    width = 1,              o_synthlcmed_postdiv.data
		.o_synthlcslow_postdiv             (o_synthlcslow_postdiv),             //  output,    width = 1,             o_synthlcslow_postdiv.data
		.o_txdetectrx_acka                 (o_txdetectrx_acka),                 //  output,    width = 1,                 o_txdetectrx_acka.data
		.o_txdetectrx_statct               (o_txdetectrx_statct),               //  output,    width = 1,               o_txdetectrx_statct.data
		.o_txstatusa                       (o_txstatusa),                       //  output,    width = 1,                       o_txstatusa.data
		.i_quartus_flux_s_to_ingress       (i_quartus_flux_s_to_ingress),       //   input,    width = 1,       i_quartus_flux_s_to_ingress.data
		.i_pcs_pipe_rstn                   (i_pcs_pipe_rstn),                   //   input,    width = 1,                   i_pcs_pipe_rstn.data
		.i_ux_ock_pma_clk                  (i_ux_ock_pma_clk),                  //   input,    width = 1,                  i_ux_ock_pma_clk.data
		.i_lfps_ennt                       (i_lfps_ennt),                       //   input,    width = 1,                       i_lfps_ennt.data
		.i_pcie_l1ctrla                    (i_pcie_l1ctrla),                    //   input,    width = 2,                    i_pcie_l1ctrla.data
		.i_pma_cmn_ctrl                    (i_pma_cmn_ctrl),                    //   input,    width = 1,                    i_pma_cmn_ctrl.data
		.i_pma_ctrl                        (i_pma_ctrl),                        //   input,    width = 1,                        i_pma_ctrl.data
		.i_pcie_pcs_rx_rst                 (i_pcie_pcs_rx_rst),                 //   input,    width = 1,                 i_pcie_pcs_rx_rst.data
		.i_pcie_pcs_tx_rst                 (i_pcie_pcs_tx_rst),                 //   input,    width = 1,                 i_pcie_pcs_tx_rst.data
		.i_rxeiosdetectstata               (i_rxeiosdetectstata),               //   input,    width = 1,               i_rxeiosdetectstata.data
		.i_rxeq_precal_code_selnt          (i_rxeq_precal_code_selnt),          //   input,    width = 3,          i_rxeq_precal_code_selnt.data
		.i_rxeq_starta                     (i_rxeq_starta),                     //   input,    width = 1,                     i_rxeq_starta.data
		.i_rxeq_static_ena                 (i_rxeq_static_ena),                 //   input,    width = 1,                 i_rxeq_static_ena.data
		.i_rxmargin_direction_nt           (i_rxmargin_direction_nt),           //   input,    width = 1,           i_rxmargin_direction_nt.data
		.i_rxmargin_mode_nt                (i_rxmargin_mode_nt),                //   input,    width = 1,                i_rxmargin_mode_nt.data
		.i_rxmargin_offset_change_a        (i_rxmargin_offset_change_a),        //   input,    width = 1,        i_rxmargin_offset_change_a.data
		.i_rxmargin_offset_nt              (i_rxmargin_offset_nt),              //   input,    width = 7,              i_rxmargin_offset_nt.data
		.i_rxmargin_start_a                (i_rxmargin_start_a),                //   input,    width = 1,                i_rxmargin_start_a.data
		.i_rxpstate                        (i_rxpstate),                        //   input,    width = 3,                        i_rxpstate.data
		.i_rxrate                          (i_rxrate),                          //   input,    width = 4,                          i_rxrate.data
		.i_rxterm_hiz_ena                  (i_rxterm_hiz_ena),                  //   input,    width = 1,                  i_rxterm_hiz_ena.data
		.i_rxwidth                         (i_rxwidth),                         //   input,    width = 3,                         i_rxwidth.data
		.i_tstbus_lane                     (i_tstbus_lane),                     //   input,    width = 1,                     i_tstbus_lane.data
		.i_txbeacona                       (i_txbeacona),                       //   input,    width = 1,                       i_txbeacona.data
		.i_txclkdivrate                    (i_txclkdivrate),                    //   input,    width = 3,                    i_txclkdivrate.data
		.i_txdetectrx_reqa                 (i_txdetectrx_reqa),                 //   input,    width = 1,                 i_txdetectrx_reqa.data
		.i_txdrv_levn                      (i_txdrv_levn),                      //   input,    width = 6,                      i_txdrv_levn.data
		.i_txdrv_levnm1                    (i_txdrv_levnm1),                    //   input,    width = 5,                    i_txdrv_levnm1.data
		.i_txdrv_levnm2                    (i_txdrv_levnm2),                    //   input,    width = 3,                    i_txdrv_levnm2.data
		.i_txdrv_levnp1                    (i_txdrv_levnp1),                    //   input,    width = 5,                    i_txdrv_levnp1.data
		.i_txdrv_slew                      (i_txdrv_slew),                      //   input,    width = 4,                      i_txdrv_slew.data
		.i_txelecidle                      (i_txelecidle),                      //   input,    width = 4,                      i_txelecidle.data
		.i_txpstate                        (i_txpstate),                        //   input,    width = 3,                        i_txpstate.data
		.i_txrate                          (i_txrate),                          //   input,    width = 4,                          i_txrate.data
		.i_txwidth                         (i_txwidth),                         //   input,    width = 3,                         i_txwidth.data
		.i_rstxcvrif_xcvrif_tx_rd_rst_n    (i_rstxcvrif_xcvrif_tx_rd_rst_n),    //   input,    width = 1,    i_rstxcvrif_xcvrif_tx_rd_rst_n.data
		.i_rstxcvrif_xcvrif_tx_wr_rst_n    (i_rstxcvrif_xcvrif_tx_wr_rst_n),    //   input,    width = 1,    i_rstxcvrif_xcvrif_tx_wr_rst_n.data
		.o_tx_rst_rd_sync_rst_n            (o_tx_rst_rd_sync_rst_n),            //  output,    width = 1,            o_tx_rst_rd_sync_rst_n.data
		.o_tx_rst_wr_sync_rst_n            (o_tx_rst_wr_sync_rst_n)             //  output,    width = 1,            o_tx_rst_wr_sync_rst_n.data
	);

endmodule
