//__ACDS_USER_COMMENT__ (C) 2001-2024 Intel Corporation. All rights reserved.
//__ACDS_USER_COMMENT__ This simulation model contains highly confidential and
//__ACDS_USER_COMMENT__ proprietary information of Intel and is being provided
//__ACDS_USER_COMMENT__ in accordance with and subject to the protections of the
//__ACDS_USER_COMMENT__ applicable Intel Program License Subscription Agreement
//__ACDS_USER_COMMENT__ which governs its use and disclosure. Your use of Intel
//__ACDS_USER_COMMENT__ Corporation's design tools, logic functions and other
//__ACDS_USER_COMMENT__ software and tools, and its AMPP partner logic functions,
//__ACDS_USER_COMMENT__ and any output files from any of the foregoing (including device
//__ACDS_USER_COMMENT__ programming or simulation files), and any associated
//__ACDS_USER_COMMENT__ documentation or information are expressly subject to the
//__ACDS_USER_COMMENT__ terms and conditions of the Intel Program License Subscription
//__ACDS_USER_COMMENT__ Agreement, Intel FPGA IP License Agreement, or other
//__ACDS_USER_COMMENT__ applicable license agreement, including, without limitation,
//__ACDS_USER_COMMENT__ that your use is for the sole purpose of simulating designs
//__ACDS_USER_COMMENT__ for use exclusively in logic devices manufactured by Intel and sold
//__ACDS_USER_COMMENT__ by Intel or its authorized distributors. Please refer to the
//__ACDS_USER_COMMENT__ applicable agreement for further details. Intel products and
//__ACDS_USER_COMMENT__ services are protected under numerous U.S. and foreign patents,
//__ACDS_USER_COMMENT__ maskwork rights, copyrights and other intellectual property laws.
//__ACDS_USER_COMMENT__ Intel assumes no responsibility or liability arising out of the
//__ACDS_USER_COMMENT__ application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version=1
`pragma protect author="Intel Corporation"
`pragma protect encrypt_agent="Quartus Prime Pro Software"
`pragma protect encrypt_agent_info="23.4"

`pragma protect key_keyowner="Aldec"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ALDEC15_001"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
EgA9JUDd6onDf4tf16+ml7dmaH9Q2WaKZImIq+2AFA1+pPzhK/+5+w/X5KQk
pGCarL0k8Jse6fVqQkjm36sPnBPx63fQs1L17kYv2Yh363Fa8Mbib7q6xkED
H10OXGxkn0cbZ0gPuQ1yVgyWydY6DT5P3eFpvwZ7+euczewiP3RVkkUKjTE2
020HzNr5QwWxCuQ4A2rv4q5eSnxHQcXEextSx2dqrzUr7Li4FvVaRbWb5pU+
8pDEo9RQh2lmLyw8A5rBNw/8K/dH+5dSva6GUL+K2whfXSRnRjAWN7Zs6s/M
6vo5iHckJMHTjThIenwCYEXXTYfjVfRV6qhGO71Mhw==


`pragma protect key_keyowner="Cadence Design Systems."
`pragma protect key_method="rsa"
`pragma protect key_keyname="CDS_RSA_KEY_VER_1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
fY6LTdIDkVM7p+USM54K+scoawFSA/akuhc4TuL9Zd/fmDBxrQAr2WkvkEKN
Ezwcg80+sT3npB+cAErrZzjcKmbziEvzdaW+Mef2BLWgeJv3u7SBm4YizhUp
TF7q0jsPMeH8073FHwEtlpfVQl9C6NfIGfOmxPOH+oX5AEr5t/iQ4fcyXDAu
nZQaqgbTrNCRzPPMvh6aNv12N9V+/PebdTDgN5vqzsIh3iYB5ubz6afb8Gf3
MD0tvV674Ptx79nhJK4p/p5QRd7MhDs3t8c+YmkuS/ZuY47elKVkDB/Plrxr
1B/cbbGxNRu9AhCfC7yZS+ubXwd4nLKPalzKYrNgOQ==


`pragma protect key_keyowner="Metrics Technologies Inc."
`pragma protect key_method="rsa"
`pragma protect key_keyname="DSim"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 256)
`pragma protect key_block
mdvB7bEQrPNl0ZL44NLVw4OVkUKRJ+U44CtsGR5Ebyi9AgDEhLiW3orTtDjV
AywYY4LsK3Ux6d3u14pV9wG2f1ikWGtX8szly/PIm4uACAgpsICG+9OE2SQj
pfxXmnR1Sktxlx0kSytO4PDUY2R8hPYie2B2Atc3Gt04J6CKKYd9qoGp2DMf
qn2vhnY8Bg2tLkh/2sEXsOF6h1FVNxn7YMd7UzPlGI4Qj5LT+QbC/9G/jwc9
AAfhaedo+6Uun3SPq0H6BBcuNCuq33K5MgsS6A82cWVzECALXpxAW+HN9m+H
UnOIIQtOmNLLINJAhCWBq+Q9KIKDyrn+emASeTP2DA==


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VERIF-SIM-RSA-3"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
nhJzvo+7lJmjlp6ncIfZP0aIv7758ooX+oyjUVB9bBP2QBExVmEjP/iQlAEy
QkcxYfyH8g6GVW9oFCpHTDZkWQZ4ngipd+3Ojtt13JmLJH36Wsegcehn5LSj
cOJQeUTQgK99IJCU27cALmmvAUIVXGjm6CiVDc9il6N41HaMp1Y=


`pragma protect key_keyowner="Atrenta"
`pragma protect key_method="rsa"
`pragma protect key_keyname="ATR-SG-RSA-1"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 384)
`pragma protect key_block
U+0afo9uZ6A0ZzQW3jWl7iPFCjQ1Fb7naBcljITGSDEPjIHGsMptZQ6NvoIH
3suRaaX00lCQjNC92ESSCsFYSj9C7S7ufleGHlhp9MsrQfJxBKFvgtRM7KYY
3kz4gHZW9AIkrWJVRAXUHXQTCl+bM3oKPLGJe5cmxfMkFJENzS4z/sGzsWvG
GX/3ObKEHSxB9CvSZMY92ATtY5nH/CY55Butd/H41JwHvdpuTw6MRXXDtKYV
xv1/d4Mb8A4+T4QqBt3hOrLmpK9frlM0BIPatW1WVmuQ6+gaP0VdzOCU66bH
XHtsJftZOTSPpDPqHojI/XuXCXFkjy3UVMQErp0MR2Gi8doz2Dka2cSXon+W
crbcb5G4S0lFd3z5Jb82qTxfRTqWv0UblAUD065goikNyQWCxvOxknDr8o22
tIscXab3ipl3HBiF6bF+teD1e0LqK4E7pwusqfydv+UMFHaSwVrooNGHg+cs
k2ok9iKnqhOZa66gajPNru5reJx7Uprv


`pragma protect key_keyowner="Synopsys"
`pragma protect key_method="rsa"
`pragma protect key_keyname="SNPS-VCS-RSA-2"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
RsGcidey8NJwYeU6pHWfkbfqTI/4BOFC/21ajuaJnzqSNbHdFb/KF3/58EDW
DbEdwpQeQesD6jCWLXKQuE+qeSDIXEK8IYtcJNRSNeTa3DyDvdD8FdKOiHoV
KIUK1rPHzrs1KZl2J3bZV8UrRiYsrlumG1balWXQyTSyo199mT8=


`pragma protect key_keyowner="Mentor Graphics Corporation"
`pragma protect key_method="rsa"
`pragma protect key_keyname="MGC-VELOCE-RSA"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 128)
`pragma protect key_block
oeLOV3jGDnWhZzLaqD6g+v9AdZpapY8zzeUHia8bdn1Jlfn9KeGRmzCZo50x
fAF2+uNVN6gqr0ZahuXwoZ7WNDUf3cgm6icgWJMFfmTNHK98+12v4g4C9S8H
kae2XjIeyjPQxLYiI5WgOCVE+4nhm8LE1JE1z8D2EusLSNeeE8E=


`pragma protect data_method="aes256-cbc"
`pragma protect encoding=(enctype = "base64", line_length = 76, bytes = 6544)
`pragma protect data_block
KDWwyHO/C9vgtux7HBCRRTXfxCAfH5tt3V8+9JH8JJESbXm6vgPkgOM42w4Q
RjnbKuSty3nHEK85BDn/EWGVUaapUMJlLnC9VecMpF3vqilICgokXuwNgGv6
qzwkgmRhR/mCFpP0kMS3lbFTUGoCJN3BjLVzyPZFIWFCBVYzXmu+8xQ17ASc
nkWBs/dv3HG5Ez5/cDKtDnQy/xXUxFSc7KZXFJce6WXmU4IwanxsGrUA1p0p
AySSttY8YbgiBxSkLnihCHNd3wS8lDgYr0882b59dXCFf7OjimuWmsEhaS9K
U7j6CdjYmIl2lxg0kR4YuFj+M9Eym3+KleBBrrwiBvJN3j+RbpDriOOkT7cl
YWn/2y+tTmQPZ7bsawNizxVimaKsEUe/sv4eQkuRtcSyp+6oM+MYWophrBMA
+NkFhwRDNruZE2qBz3nI+AqjQWba0FN6I11joNs3tKiVK98N8TAwNZk/qUVo
V6N+v0JdcqZdw8k2hVl6wl7ddd0JWIVhUcddHYXkpXquHqXEmuBlnZ0ErrS8
YkvS3CF0zuNfd2AFm9fdGuEIoMQtWI+ruZUDggNIhBbOIUfAxNYbRzvo0B+K
P0bJzKY5oPLTPVRSwhHtO1N0Rk4d2I8qr+FfFAMzjlhksQw0AVk+JOcNuoYv
BO0EipZfwxMu5DjNQYKso3X1O3+IBNAeXMA/Xj9GfvBAeL9dHeEI3ycfFkp2
IPN/gERsaQYW4aPEwdZdstWR9I8yOXbp2ZlWVb0hqLRDAPB/LVEbmef+SYxc
o0eGubqbNvrQ5FuE+SpmZ8lQjz5kYqPXxyqIlYURbs98hnfq/n21j2X/rpAb
nyyh+O6TBv8izbqI4llRUt8IZPZOHjgW0h3abNV9xErDWSEuuF/8M6ntmSAA
MK9/4XE0xd9O2LKizQkTQu4dQFVOciZdlmK+6sHDOke0KIVfTZ190sYZQnvA
Og2qAytBKvpyIrX3hp4CY1lJrbv6f392E6czfL8GLBW5Tgn4pH4QYh9DY0JL
7dbMwcbNJC1TW2CFhCP1RgD1J0g464FrizOnD3vjVM2zFwubOAQ/1iIcrSZC
YcJocas4tGYDUovX7cnTyoT9ugrNnVHYl4eZnCjTESzy9MpXlSf78tIK0o6C
uj8zYsGlxfqNjIAqb9xtHiJ/qxtBmlLL1rAVHfJanLdjEAEHIADzrAnAhAh9
c/LYm9q1cBSdx3FKSJzxVLScABmSga93TiBmG38iZAQ/DVrEPghpWi+7wYPO
CgYzFm9Ae8VUyuPFpAoLWtzAeuGNJhgERdp2h6IKOJ3nCcX50eDrTuIaPjKg
khBsHBCBwk+hRO/8SxNHV6NCTAZHeYl4eXZ4f7W6XYVVIrSS1JF/6M2QpIye
sLgpEfDmtN115QrxCmEsRKh7ymrDUGVPa3hEDm0PITDTzdiZX26a8RVsPxVB
ZBy8IhXy6CiOnHKm+lLNyPo9zr+ZtGunsZUFBLwt3FFhYNeHNfcFeXLg95DJ
Qd1hlS16hEp3P5dnTmy4mGdzOf80IR356IoYLyRyktiacuC31JzgaeeBu45Q
7jYSKiOd6z03YPJ64pqvwjyow3h+SF5PaUKfha01XLOIGo2xRLlO07NMDMgs
1+k2t9O87Yi2nY70xzF/IcwqZPWoSSZr8wt6c0KbzTKct4pPJBNmnC6HXlOZ
9GMDgUCFzS+lsHQx+ftEMpDwTZ7ZHxXnrB0gdQL9f2biNil2pi9SYXi66lJ/
K3CgXFi8Abb4S/sK/vxMKF27wRqMrJ0EUfp2S/yNQ0pgxqbRUgR2t2LYMb0c
wFT0atLmcwgVd5HMY72zKnI5N/NPjkIPHAMnAlGTIaiNAEW6R3NVHEua2et4
U0JEZPqJ20B4ZASaan6AKINqMS1XKI0wuGTxD0GHW7h2LwdBRila4v7GhgJf
mUUU8jXjYrOrD+wpczQbis6L980W6JXFuWg07b47qEgUxpdjq7Sm7gKbiVBw
25KvEPqAFMhd2ijSdM+hDxt8FvXxuSu9mtAc1L6iOO+TPP+Oyf3RqdvSDToh
5Tja3ofv/R96XdljIBxFTKRTr54XHPyxvaCj2K7ibDp38mqsQlrSnt4ad6cG
RQHETBbVn3wQi+C3lOR7f0slSYd4hSCRyyMTeW+AJN7FrlEclfMxrdTfoiwQ
o8nxEAgFxhoodb6bC/6T9D0xt+M3msnWv29AjYyKgVSEjfWKakMu1NpsPjfH
pot0kxq4eqWtielygyQqNzKWu/YVajhLmJED1pzEhf4TnoOHyVWkkT2jflR8
Li9jP/U56caKpdwp7yzOBFuRjey4h46bFr+AQcgcF263LgrnMgZZLoemLC3l
G0lH/p+7FovccOa587guk0PPlcQRUSlQxnyzEX/3NVU7AQw6CN1M2i17Bwgd
ZNEd9YPAsfla7dPgO5AnGzfUkySgfKxN7lT+aGc+3M8OHh95MhrwShIQ7F0O
SQGVY1uo04Eq++YA9Tw2zzVul+iAL5thZmfWqK5dIUmTd3e3QspIr9vWsvtf
yxiODUTZ1d0+cCYwMXvd0jgEc8opgM3iTkfpu5/+YjMbKegoN1Z84eGuUc8Q
JV5j2urARfT6v+xrK/JD6HJypNcY6eOFCn41LmjlAQ+XHyAVQ2o440XrrBTD
NRAmTgUdzMkWt8H5rAGTcEUP8BDFFQvfHN29r/Vz8Rd9RUgcdXs2RUUjDeEv
jBCCFPMYfRRWd5OS2QOlJ3S28x4aD/zGSDs/LdTSrfepicbKvyiCCijZ4y/h
spifBfO+oa+TY6rdoC1ar4Q2EpS6cFzbtxnKFryZ68mkiTDnVOz2wWb0BL0Q
JU2Fk8u45lvLWimtmAcqeXiAboA/fIbQSaVLDjQrGKA8E7vtp/v21uCduPC4
uj/TAseWss366K5TP8ztIitn5GicSL5RBkyhvHnsOl2Wq3lL1/+x8YIITJys
RkwqIwDtCoUeHX+3vhKjuEAU79Kj94ARJt1mM9GrTXiqz2h8xE/nsjamS32z
y/i5P+2UQRY/8SOq+Ul4W57XiV1VTmDf0S79vhwq+CQPw1VyjIzXtzINEJF6
s7mrVBtJdl/JaTkCkXfQAA7fpsb4Idq3VCb4qTnT5jRbIChfj7F5/EUx/AjF
zMhYbxl//UU7E0rgp0kDLbXuavTgy/CV9656ZaGaW6Y1QrL9NSd3e7Rxl+06
Mp+G6YhCL6ZGpIi9X40u97xlaiZN1uJ449bw7Y0D/6YlaSWCNSDaoFE0n70O
yeTP5o+Mx3BYtNMCmv2UxTTAXJY4Rlg5KeLYfyzwbADi3YhosfWNnDD9uRRO
epmF84FBviNF6kxejUchC50X5/I49Y7Dtla8iu7ugtA9gxZ3nUlDTbPKPAef
ERgH3T3M5hBU+7tNau5/HZTegcojzYQdGjAS9yGtiXLkJRPqKulmo2q3CZAW
nveM+qy9RxDVY9FSI+ltgBuMOUeScGS6GcT9/qcFRaEcN2jdRTB+Mt+pylPZ
19uwgQNr/AXcnGEZIe67YFbZj4RFUl79W0WlldPuFWDxYOuDX+31LTDU/mNs
tJNCL+vEnMsKrOv+VT0hOZhpex+gduynSIj2lGQnxEeXNU6YEquFGVD9l6bj
JSkt1fDrcWZnOIFXFo7uO+thhVTtBGmBAqw49I9m2LD3ExCyGr2wjkLlmS5B
hs7Ew9qS25MUuYw3hG/NYaCnUDKbECmPj2MHyMxh07Jz96F7VNMpz+iw4LRe
H+2h/qpQ88suEHSdRE56HT1PMq28yMhTSKu++gdaiKXQ2ZBKCg9RFxtzvrPk
L/pWhNk0ncH8D1VbISuZvNKOIrwlnyt5H9i2Ks3bW5drH85hzoYzc3bGgbGs
QBwDLNCECJ+UBrp/eBOTzfBoOKK6zRHqfEm5U9WOQmFSEZRnB723fVOcZm04
bKr+TxGj9cgW1GHqtAaQiMI9e+pgTwOCaxjetF7GhF3IcmF1YUTJfjoOunL5
wQ48XZhW5Uz6N4+wmeNUm00iADeyol0CZ4eulJTlPe6sp829fDIOVQLAUfe0
iNrpT2ScptWd9f3o+4HAU4yP7iVUrGOcxcXyj7+CZHuTZdUt6s/gD/pIJ8x8
uClvc79vgt+upDZOJY/xeQFrtyhC28yZlm8PnX+1oIdp5J5ypFNkKocCOZxI
skX0z477kJtX09t8NZ3UzUBfWj8JqPMvRytBW6UE6+9ZudKhKdtWOeE1Txng
bXY7XnRSF1A1EWXVNZqAR0UhFwPM2ZpH+LcubQDcmFJKynhjIrG/5h7amvIu
tpOsNa4SA6LzGcsh37C12Jv6IC1PF6l1pQ7MktWv1eFFCYa7CKX+6Lx67/fO
0xyGo3hyucjM5eNCYYbV1lMnmXp+z+dXfNR92rLgP6aK0Ne4BPdTTZpGfHKg
dVpWm6rlEqgQbgyxAoVgipJiB+9TnmAc3Ge35w7GokjK4yAbxORoAaR4IRjw
C3VyiXLDws2zkQh0OpSNc8PnmkWn7DNr4BWgPPLUALP9PRxBnXfsXAFyXCAD
Cud6boYYW2jQHNt4SWxVcgBP7ln0GTPe+WnDHnSZqWJyWw+3Q9czIXMj4pbL
8zxabC8VTsn5QvKBMgcZB35hmkh7aIPIpq8EjZjkD/g6QUKLy5OTMcXRY20Q
cVuvRNrVPll0grnBiv7xRLwqQ9FCN4boN8y/1hAjks3kGrvCS8rUMZAIKy9u
loIuuCK6ikjIPrXPU66fO/EqybIcsxBibCTVsMHGdwu9o7KS8Fc2GRi71hyj
BDXzKLDGYiuBk/PR8YFKE/2IaAzDWpTVjrPfedKaDuBEU9LruYwnEokKi2GC
OyItyify1RvhUqxQOonkcG64ojRifSu6sC9rO0NZ9SglcYucdQEwBNsthH8I
RoplFOvQ+QrnDS3ZRxsDakFuPkHTal8NGFhaFxowYXhNouCpPB4zU647mt4B
Hy9ZY8zbtdBIveOjVF28p51QxG9AB5IlGYpSLRNAaqTyeVltAY/4VjutSRN4
lpZKMCUtl2sj+FypeUWqtda4Gl+MaLcQP00HklU7p28GQ/HsoXSiUokIpFGM
Ig9KOV3P8IbaCnrLBAsE3Li+UrBXNow66G57YRHNiFgGrOFBO/kPfeLy4yKL
tZitRHmFb7IxJyC76JiXX/TM9rSkA4YT2FWimSl6cDyQssSZ+hB69b9CIUKm
Sqfi7MqiTT5TNCrMJOsJAud/oRQA2GX8ujHcK5qNAOKjwXZMYOD1HbjRYBL9
uN2zGt4/jFGJXX6sbKTBiE5R/xvgVDG6LvTyoiSwEOv1q+3Ngu7wub8CKHh6
/HZ3YVovCwlndbAEPSPPKnDLx+r/LYE/5CutxPfiJktwAXTeG7n5t3wlSP4+
H0Z/VBpYUA78KcLv4LQP3riV3fWHaochXg0vhxzDMBxhMlkTJiYK6X3gl1LF
oZ2jX0roR47nz51JjLqccMww/UKM1ibkGKj+aRRK5WFxhQ+ojulZUc4njHHY
ukFAcAi40VKi/C/npjKgZe/yeEadLXgc49yrwO0oJgLcykL0ca5yApgC8mPF
ANu95s9RWhunhBEyj5coCbBiRtNFJcgF4A515pjOjZ45YtmL4UV3iLV4wu8S
9TDeiMj8HL+fDIEa7w7jdYoOtwBZnAa+OSLtcgErYOY7Lzu7HpjkGBfDUCt5
5MKRSja5B5a7la1BeQwVeJPDO+/nibZ3w15OpKwjXFxL9YrQMcupAjbedoLK
dQ78sKAMnmDas3EQzwaYogZ4o7qv+P790RQyxLDXnYN4Ao+PLrIc7NTKu+W+
p8IzzkiO/lUAAOecj8YUbgchXAlAGI02JA6nYsJJGAvijy6xSz0u8L6lBu6Z
i/Fn24uxWVZ6hKv8wiB9KSEY44/JclOFrfC26zkRt4CvhDdXcMzy2MJ9QDDk
dk4+68WNYF05P1yFYBPTtA+RGx5Yn68ZtG5Ufn4nM1MzA+oIUS8bP5xlx3Xj
rpFMmaKI77fOu8ZxIrBzuLraGXyj0sv8kksB53OHGTgplGdkwcOTO1jika2D
6C1ZR5IZy11rmqd+zqYnCfOY+49CiHJLTCkZsyYEqTwFBK7/02eT075gI3tR
ZnXZ5HUSIg0DZlspQlakpk3/el0aSxNPV75kyPGXQT/ZUO+bwxRgKDJXU78K
YoUO0nUGkWaSfAh5KqxIAWh001oZfG/iCUAcXjNu5UH85hIWMPK69B01jSe+
ymXJQ2rwPoHpc45B6TO4diwEYXlKqr3NACmYYHiuN4PilRnDt1MnCdnO8GVK
V0EeU0jYopIWCCOIDhhZq9uLVe9qRBCbjzQSYAyXbjbsDwf6gtYfBBmLPM48
MjciFOytU6jxYlF3ixiURRj1LNc99H0AQcy8xWlRY/qQyNQqdHt+aQO0v7lk
nxoA4B1Z1YWlqTPhM4TqoD/T6dHBvER2Nvcn09ZZ1tMOpLr8ZORphEvWDtRw
NB3O9MtdPTDpUpJvbXkhx9k/9U+PfHp491DPzHPaWPHB3wf4OVAvNeJLbTiU
HWEqcb6HyNewOh/+++87B9eHr+6KeopwcII/5VF9mHYOP3HTVTzfyHIjvYoN
o/fU+1EyrK7awUmWKUUQD64qrXv1wmj+iV9h+gJp7V61/5upRKlV75v5Q54x
wLCfwlgaWzIlMWbF2Xx6WblkrPEflQFGHE/EhAonG7NyuJwm6GjqaelPWHxS
U4qRK5XY8PnuoU3HRSqas7+rt6BSzX6tH0uhzZU8Ww5axMP6llSYjA+1C/UL
CUaY2aUc/ajv3Lfz9f3u96kR7BvrA80J1DdzN35ctkLse3M++n91O3dpuTxw
iBUjaIC+DEzEGkolMeHaYOg0qMBvJMvqYW62ghWTX3DglVkp8Yf7nsB3H1rs
7EQLxu9WzHAV91E2cKCKAlnzCeKrnaHtVE/E5XrGDddGYxd6ty5LCqFLMkVp
ykaMMrsngT0JwCCewEyCN1sNee+lbS9LRwp6/fi0f9erz3CV8h+c6WON3zto
yQHx9kCbHSqrNGmxL65JcbUzHLWjeqiV1PYAg97z2sLRhJzqhRkvm5spOmmn
+1vQgfv9tJ17S+ukGOgSHXwONiCo4tJ6r88BmCiuiV9mh2vu7510UyqP+asD
UJeQZPM90+CHtrBw90+/D+7Mzi6M9En15NQYYiQqAeEi72/dRpCqtmAFCgaV
5ZzuE1ioNWbcaIJo5kerKrxZU75iPNybgUgeD4j1uBDZUCRcqLr+mX2Pi7tn
BNUNFedSaV1Jfb8jLD1dFOs1HoTEudP0OjU7WRjNexDZDXVc7bw8IhxQgdiV
rFx+81aNrQk2a5CADZ7vdI/5/T4jLz68gr5CFmeeJZiPynJHfyauO1129Hhn
ymvXLUhsr6NVn96gvizenZ7PZqfFta4J8Ye34zia7jzqyGEOAunoYzaZVrI7
XpGWePdpnro4hRr+IUbXXeqU7UC7TRqc9pQLObCaDV7REEXV38weqgZTnQI6
2SD2nxgOqEptgxiOc4JhIf3DAGlliZv7L7hVKMWmQSN676d6MH1hzbdOS7m1
YyfcQ+0s3otdKDjbt91srRkfxs8O6WQKBTH5xjuQjs3GfOtG4iyInehrY7Fz
vAaOCsJBygpvbgNPSKm6ntBwPMloOZd3XrtBGE9gpDjt59UDGxK4okrDaKDq
rGNGhOezOqn6bXecnf0qEkg2hLeK2trkWtH+6w8VLd70OK3ySFvUutbkLBBy
C9bwId4B4Cg5kQh4Zajl38MbP5wViuWW98QXal5Ofw/eUbRekhoPKtqAuQ55
P70Hsxv9301ANhg3fA36BF0Fm7LJK2Fgv5ola4QFhJixkHVZTGYFVfvyYYmL
cStBaF6mAPRHvAv8xQNpXtWv+JAKMTbLxYN4oHPPVf82tsKOkFw9icnITB5w
P6WzMCcbKn0hwP5trLdGIqNaZCz0mTul8tOS8TXDEYYxmimnJ3FJWclwqeau
vXsbJafqDDcZrTt7cpksYpdfxyp9d3rIPT2rMNAhHbzcuelgI+gm4HXmtWSF
fBffD6jtLWBmMuBQ0FF+AvaJG9UL8TsbUIRuakDF+VE1zYN+/JbUBPwJiZi8
0tFFe23oAdLSAmK7MyQh25r6mjXZn5sfubORpDL73in/vx9D/3dqptp+oN02
pgQMZkXRuEhOPw3t/E6QYqO5kUTUXYJSQPd+EOTeLPjt41oDdmKlTmkQu8I/
L6E1qXmGtUk8/KySh9gJZ0Cg6dCzd8pFj4LVXK4BzvUJESBZ0Mfv/aGU6OXF
gMnAWsXCpNvKJW1h3Nxx61NUjErwsgTr1zGl5PWbtAomvopwAYj0oDO2BN42
z86m6NTXPxdh2oBvm2QstW54AYlZUyHS8gMiNlblso7bmyy//WwPjVo4G35m
MFW2ZqRoQVGrat3VcGKOofQCfL/I+jikK8HORT4sQdSnW4AV0yUWiHu6ifF0
hAXubD7B8/CWVB6DDQkERO/x5ZyCqAmV3KajRCiohruQHe7+iqnURBHNf9TP
Z+270M7irOz5BoH0TzbqpDN8+pDz6gfEXbCEGJcDVIVCfUMbWsqMaSEweDco
TbRSMWHwltsZelFJQ2hm08TdePAIvQFpnYrIxuqGOHwNMKNTS+issaaaHRUC
zhjgIvWThizVaz9ROy66otK4P9negABNBSbB0I7lHorot+PXC4HvOFEwfFzC
XGL8CnG9O2T6tEKxPbEDgnAOyQiO8Fa4RcT8OcuGKZoDeLj+BoVm3W/R5EHb
gJ4NP5+cKHNE03UB/ZP77ZM2fA==

`pragma protect end_protected
`ifdef QUESTA_INTEL_OEM
`pragma questa_oem_00 "CbILi0GnYjtEWmRNKNj5RgNJK0IIz5zHSE9Rn/kaB55CqsFyqlUKVKseihpN4QkCK4D726Y9yxpvlkEEsZuFI92T0NPCHL9iV6nI+RWTU0V3MdmpYPJwm+nH5bs2hSnHBSgZxX18LPDGkO2/sGZW4UdapTeyyaVpJ6ym1liwBhwGIdZtW4LQKQJrPf/6wnW3RDZ6dM4mMlryGqZ7J4MUifJGwse2OmTGHm1yGaKAJ+nJbOBbeStJFbgxI1uAamJIr2978BFFP6KjGY4E3LOqPVpBrJWvJ1mx9keP9MSmUCT8tIrLZPyn1lT7AqKvL9m75uPELDtBLUEWYTxxhQCJP8p7QtvDTEZQbOJDE1AIOTQMBOpy4lvHO562+1Ru/kk9b2CYtfPdYBDv2TjPkgzOi80kRb//JwXkIQUISLUIIA26x8JzouRVhuHno92VLPbNqnCuDvJfKfukyVdMK4bR87vv2ccFMFJB+iECFZjzN4KO1iVEMfKWJ5iJZ0ffS/W6PZiIN7scmWOL8F0/cFPuSGOE1R8arhu8Q+X5jEIFlTqWF0rcF23PUSzb6x92vXdiOKtGadnTORVOUvtWoPIdPO5e55J6YOlb5UpAnoM/kwy8KeuoWBJWlHX3sEt2N4kBsQ4Ka7hVfuqIjMfR7lIMQxUqvtaK6S2sSkR0O8A0Lh0/3pYN0k+DheRT3cDYtnd0yUNNEhQ4pERNFpeZw7luUHjwyM5X2NSgQS8WMC3378KFow1AA6hGTjDxcxqVQ4kgkam3GZNpq63PlspzbqQ7jhZJPZrTyyK597e0B0LE4NKTP1mMJCYagid2fxBTEvgRJK3aC65ZeOUcg/Sg1Y6JO3btPi52rKal6xWDfeB6ETiybMplDxl0gMXSUXCpFvfHDWvVConEo7XNYVCzLrbXhOS6/o3gJBmtCfWwDGlS8esE5Zm6YZgCyQ1u0eSmHf2sJ0bCUA2cOL24/vgd3+g/Y2QbT7qXp3hPkOJx73sjPyEr1OjvHu79jqCvpMz57pmM"
`endif